Då skall Moab komma på skam med Kemos, likasom Israels hus kom på skam med Betel, som det förlitade sig på.
Huru kunnen I säga: »Vi äro hjältar och tappra män i striden»?
Moab skall ändå bliva förstört, dess städer skola gå upp i rök, och dess utvalda unga manskap måste ned till att slaktas; så säger konungen, han vilkens namn är HERREN Sebaot.
Snart kommer Moabs ofärd, och hans olycka hastar fram med fart.
Ömken honom, I alla som bon omkring honom, I alla som kännen hans namn.
Sägen: »Huru sönderbruten är icke den starka spiran, den präktiga staven!»
Stig ned från din härlighet och sätt dig på torra marken, du dottern Dibons folk; ty Moabs förhärjare drager upp mot dig och förstör dina fästen.
Ställ dig vid vägen och spela omkring dig, du Aroers folk; fråga männen som fly och kvinnorna som söka rädda sig, säg: »Vad har hänt?»
Moab har kommit på skam, ja, det är krossat; jämren eder och ropen Förkunnen vid Arnon att Moab är förstört.
Domen har kommit över slättlandet, över Holon, Jahas och Mofaat,
över Dibon, Nebo och Bet-Diblataim,
över Kirjataim, Bet-Gamul och Bet-Meon,
över Keriot och Bosra och över alla andra städer i Moabs land, vare sig de ligga fjärran eller nära.
Avhugget är Moabs horn, och hans arm är sönderbruten, säger HERREN.
Gören honom drucken, ty han har förhävt sig mot HERREN; ja, må Moab ragla omkull i sina egna spyor och bliva till åtlöje, också han.
Eller var icke Israel till ett åtlöje för dig?
Blev han då ertappad bland tjuvar, eftersom du skakar huvudet, så ofta du talar om honom?
Övergiven edra städer och byggen bo i klipporna, I Moabs inbyggare, och bliven lika duvor som bygga sina nästen bortom klyftans gap.
Vi hava hört om Moabs högmod, det övermåttan höga, om hans stolthet, högmod och högfärd och hans hjärtas förhävelse.
Jag känner, säger HERREN, hans övermod och opålitlighet, hans lösa tal och opålitliga handlingssätt.
Därför måste jag jämra mig för Moabs skull; över hela Moab måste jag klaga.
Över Kir-Heres' män må man sucka.
Mer än Jaeser gråter, måste jag gråta över dig, du Sibmas vinträd, du vars rankor gingo över havet och nådde till Jaesers hav; mitt i din sommar och din vinbärgning har ju en förhärjare slagit ned.
Glädje och fröjd är nu avbärgad från de bördiga fälten och från Moabs land.
På vinet i pressarna har jag gjort slut; man trampar ej mer vin under skördeskri, skördeskriet är intet skördeskri mer.
Från Hesbon, jämmerstaden, ända till Eleale, ända till Jahas upphäver man rop, och från Soar ända till Horonaim, till Eglat-Selisia; ty också Nimrims vatten bliva torr ökenmark.
Och jag skall i Moab så göra, säger HERREN, att ingen mer frambär offer på offerhöjden och ingen mer tänder offereld åt sin gud.
Därför klagar mitt hjärta såsom en flöjt över Moab, ja, mitt hjärta klagar såsom en flöjt över Kir-Heres' män: vad de hava kvar av sitt förvärv går ju förlorat.
Ty alla huvuden äro skalliga och alla skägg avskurna; på alla händer äro sårmärken och omkring länderna säcktyg.
På alla Moabs tak och på dess torg höres allenast dödsklagan, ty jag har krossat Moab såsom ett värdelöst kärl, säger HERREN.
Huru förfärad är han icke!
I mån jämra eder.
Huru vänder icke Moab ryggen till med blygd!
Ja, Moab bliver ett åtlöje och en skräck för alla dem som bo däromkring.
Ty så säger HERREN: Se, en som liknar en örn svävar fram och breder ut sina vingar över Moab.
Keriot bliver intaget, bergfästena bliva erövrade.
Och Moabs hjältars hjärtan bliva på den dagen såsom en kvinnas hjärta, när hon är barnsnöd.
Ja, Moab skall förgöras så att det icke mer är ett folk, ty det har förhävt sig mot HERREN.
Faror, fallgropar och fällor vänta eder, I Moabs inbyggare, säger HERREN.
Om någon flyr undan faran, så störtar han i fallgropen, och om han kommer upp ur fallgropen, så fångas han i fällan.
Ty jag skall låta ett hemsökelsens år komma över dem, över Moab, säger HERREN.
I Hesbons skugga stanna de, det är ute med flyktingarnas kraft.
Ty eld gick ut från Hesbon, en låga från Sihons land; och den förtärde Moabs tinning, hjässan på stridslarmets söner.
Ve dig, Moab!
Förlorat är Kemos' folk.
Ty dina söner äro tagna till fånga, och dina döttrar förda bort i fångenskap.
Men i kommande dagar skall jag åter upprätta Moab, säger HERREN.
Så långt om domen över Moab.
Om Ammons barn.
Så säger HERREN: Har Israel nu inga barn, eller har han ingen arvinge mer?
Eller varför har Malkam tagit arv, efter Gad, och varför bor hans folk i dess städer?
Se, därför skola dagar komma, säger HERREN då jag skall låta höra ett härskri mot Rabba i Ammons barns land; och då skall det bliva en öde grushög, och dess lydstäder skola brännas upp i eld; och Israel skall då taga arv efter dem som hava tagit hans arv, säger HERREN.
Jämra dig, du Hesbon, ty Ai är förstört; ropen, I Rabbas döttrar.
Höljen eder i sorgdräkt, klagen, och gån omkring i gårdarna; ty Malkam måste vandra bort i fångenskap, och hans präster och furstar med honom.
Varför berömmer du dig av dina dalar, av att din dal flödar över, du avfälliga dotter?
Du som förlitar dig på dina skatter och säger: »Vem skall väl komma åt mig?»,
se, jag skall låta förskräckelse komma över dig från alla dem som bo omkring dig, säger Herren, HERREN Sebaot.
Och I skolen varda bortdrivna, var och en åt sitt håll och ingen skall församla de flyktande.
Men därefter skall jag åter upprätta Ammons barn, säger HERREN.
Om Edom.
Så säger HERREN Sebaot: Finnes då ingen vishet mer i Teman?
Har all rådighet försvunnit ifrån de förståndiga?
Är deras vishet uttömd?
Flyn, vänden om, gömmen eder djupt nere, I Dedans inbyggare.
Ty över Esau skall jag låta ofärd komma på hans hemsökelses tid.
När vinbärgare komma över dig, skola de icke lämna kvar någon efterskörd.
När tjuvar komma om natten, skola de fördärva så mycket dem lyster.
Ty jag skall blotta Esau, jag skall uppenbara hans gömslen, och han skall icke lyckas hålla sig dold; fördärv skall drabba hans barn, hans bröder och grannar, och han skall icke mer vara till.
Bekymra dig ej om dina faderlösa, jag vill behålla dem vid liv; och må dina änkor förtrösta på mig.
Ty så säger HERREN: Se, de som icke hade förskyllt att dricka kalken, de nödgas att dricka den; skulle då du bliva ostraffad?
Nej, du skall icke bliva ostraffad, utan skall nödgas att dricka den.
Ty vid mig själv har jag svurit, säger HERREN, att Bosra skall bliva ett föremål för häpnad och smälek; det skall förödas och bliva ett exempel som man nämner, när man förbannar; och alla dess lydstäder skola bliva ödemarker för evärdlig tid.
Ett budskap har jag hört från HERREN, och en budbärare är utsänd bland folken: »Församlen eder och kommen emot det, och stån upp till strid.
Ty se, jag skall göra dig ringa bland folken, föraktad bland människorna.
Den förfäran du väckte har bedragit dig, ja, ditt hjärtas övermod, där du sitter ibland bergsklyftorna och håller dig fast högst uppe på höjden.
Om du än byggde ditt näste så högt uppe som örnen, så skulle jag dock störta dig ned därifrån, säger HERREN.
Och Edom skall bliva ett föremål för häpnad; alla som gå där fram skola häpna och vissla vid tanken på alla dess plågor.
Likasom när Sodom och Gomorra med sina grannstäder omstörtades, säger HERREN, så skall ingen mer bo där och intet människobarn där vistas.
Se, lik ett lejon som drager upp från Jordanbygdens snår och bryter in på frodiga betesmarker skall jag i ett ögonblick jaga dem bort därifrån; och den som jag utväljer skall jag sätta till herde över dem.
Ty vem är min like, och vem kan ställa mig till ansvar?
Och vilken är den herde som kan bestå inför mig?
Hören därför det råd som HERREN har lagt mot Edom, och de tankar som han har mot Temans inbyggare: Ja, herdegossarna skola sannerligen släpas bort; sannerligen, deras betesmark skall häpna över dem.
Vid dånet av deras fall bävar jorden; man skriar så, att ljudet höres ända borta vid Röda havet.
Se, en som liknar en örn lyfter sig och svävar fram och breder ut sina vingar över Bosra.
Och Edoms hjältars hjärtan bliva på den dagen såsom en kvinnas hjärta, när hon är i barnsnöd.
Om Damaskus.
Hamat och Arpad komma på skam; ty ett ont budskap få de höra, och de betagas av ångest.
I havet råder oro; det kan ej vara stilla.
Damaskus förlorar modet, det vänder sig om till flykt, ty skräck har fattat det; ångest och vånda har gripit det, lik en barnaföderskas.
Varför lät man den icke vara, den berömda staden, min glädjes stad?
Så måste nu dess unga män falla på dess gator, och alla dess stridsmän förgöras på den dagen, säger HERREN Sebaot.
Och jag skall tända eld på Damaskus' murar, och elden skall förtära Ben-Hadads palatser.
Om Kedar och Hasors riken, som blevo slagna av Nebukadressar, konungen i Babel.
Så säger HERREN: Upp, ja, dragen åstad upp mot Kedar, och fördärven Österlandets söner.
Deras hyddor och deras hjordar må man taga, deras tält och allt deras bohag och deras kameler må föras bort ifrån dem och man må ropa över dem; »Skräck från alla sidor!»
Flyn, ja, flykten med hast, gömmen eder djupt nere, I Hasors inbyggare, säger HERREN, ty Nebukadressar, konungen i Babel, har lagt råd mot eder och tänkt ut mot eder ett anslag.
Upp, säger HERREN, ja, dragen ditupp mot ett fredligt folk, som bor där i trygghet, utan både portar och bommar, i sin avskilda boning.
Deras kameler skola bliva edert byte, och deras myckna boskap skall bliva edert rov; och jag skall förströ dem åt alla väderstreck, männen med det kantklippta håret och från alla sidor skall jag låta ofärd komma över dem, säger HERREN.
Och Hasor skall bliva en boning för schakaler en ödemark till evärdlig tid; ingen skall mer bo där och intet människobarn där vistas.
Detta är vad som kom till profeten Jeremia såsom HERRENS ord om Elam, i begynnelsen av Sidkias, Juda konungs, regering; han sade:
Så säger HERREN Sebaot: Se, jag skall bryta sönder Elams båge, deras yppersta makt.
Och från himmelens fyra ändar skall jag låta fyra vindar komma mot Elam, och skall förströ dess folk åt alla dessa väderstreck; och intet folk skall finnas, dit icke de fördrivna ifrån Elam skola komma.
Och jag skall göra elamiterna förfärade för sina fiender och för dem som stå efter deras liv, och jag skall låta olycka komma över dem, min vredes glöd, säger HERREN.
Jag skall sända svärdet efter dem, till dess att jag har gjort ände på dem.
Och jag skall sätta upp min tron i Elam och förgöra där både konung och furstar, säger HERREN.
Men i kommande dagar skall jag åter upprätta Elam, säger HERREN.
Detta är det ord som HERREN talade om Babel, om kaldéernas land, genom profeten Jeremia.
Förkunnen detta bland folken och kungören det, och resen upp ett baner; kungören det, döljen det icke.
Sägen: Babel är intaget, Bel har kommit på skam, Merodak är krossad, ja, dess avgudar hava kommit på skam, dess eländiga avgudar äro krossade.
Ty ett folk drager upp mot det norrifrån, som skall göra dess land till en ödemark, så att ingen kan bo däri; både människor och djur skola fly bort.
I de dagarna och på den tiden, säger HERREN, skola Israels barn komma vandrande tillsammans med Juda barn; under gråt skola de gå åstad och söka HERREN, sin Gud.
De skola fråga efter Sion; hitåt skola deras ansikten vara vända: »Kommen!
Må man nu hålla fast vid HERREN i ett evigt förbund, som aldrig varder förgätet.»
En vilsekommen hjord var mitt folk.
Deras herdar hade fört dem vilse och läto dem irra omkring på bergen.
Så strövade de från berg till höjd och glömde sin rätta lägerplats.
Alla som träffade på dem åto upp dem, och deras ovänner sade: »Vi ådraga oss ingen skuld därmed.»
Så skedde, därför att de hade syndat mot HERREN, rättfärdighetens boning, mot HERREN, deras fäders hopp.
Flyn ut ur Babel, dragen bort ifrån kaldéernas land, och bliven lika bockar som hasta framför hjorden.
Ty se, jag skall uppväcka från nordlandet en hop av stora folk och föra dem upp mot Babel, och de skola rusta sig till strid mot det; från det hållet skall det bliva intaget.
Deras pilar skola vara såsom en lyckosam hjältes, som icke vänder tillbaka utan seger.
Och Kaldeen skall lämnas till plundring; dess plundrare skola alla få nog, säger HERREN.
Ja, om I än glädjens och fröjden eder, I som skövlen min arvedel, om I än hoppen såsom kvigor på tröskplatsen och frusten såsom hingstar,
eder moder skall dock komma storligen på skam; hon som har fött eder skall få blygas.
Se, bland folken skall hon bliva den yttersta -- en öken, ett torrt land och en hedmark!
För HERRENS förtörnelses skull måste det ligga obebott och alltigenom vara en ödemark.
Alla som gå fram vid Babel skola häpna och vissla vid tanken på alla dess plågor.
Rusten eder till strid mot Babel från alla sidor, I som spännen båge; skjuten på henne, sparen icke på pilarna; ty mot HERREN har hon syndat.
Höjen segerrop över henne på alla sidor: »Hon har måst giva sig; fallna äro hennes stödjepelare, nedrivna hennes murar!»
Detta är ju HERRENS hämnd, så hämnens då på henne.
Såsom hon har gjort, så mån I göra mot henne.
Utroten ur Babel både dem som så och dem som i skördens tid föra lien.
Undan det härjande svärdet må envar nu vända om till sitt folk och envar fly hem till sitt land.
Israel var ett vilsekommet får som jagades av lejon.
Först åts det upp av konungen i Assyrien, och sist har Nebukadressar, konungen i Babel, gnagt dess ben.
Därför säger HERREN Sebaot, Israels Gud, så: Se, jag skall hemsöka konungen i Babel och hans land, likasom jag har hemsökt konungen i Assyrien.
Och jag skall föra Israel tillbaka till hans betesmarker, och han skall få gå bet på Karmel och i Basan; och på Efraims berg och i Gilead skall han få äta sig mätt.
I de dagarna och på den tider säger HERREN, skall man söka efter Israels missgärning, och den skall icke mer vara till, och efter Juda synder, och de skola icke mer bliva funna; ty jag skall förlåta dem som jag låter leva kvar.
Drag ut mot Merataims land och mot inbyggarna i Pekod.
Förfölj dem och döda dem och giv dem till spillo, säger HERREN, och gör i alla stycken såsom jag har befallt dig.
Krigsrop höras i landet, och stort brak.
Huru sönderbruten och krossad är den icke, den hammare som slog hela jorden!
Huru har icke Babel blivit till häpnad bland folken!
Jag lade ut en snara för dig, och så blev du fångad, Babel, förrän du visste därav; du blev ertappad och gripen, ty det var med HERREN som du hade givit dig i strid.
HERREN öppnade sin rustkammare och tog fram sin vredes vapen.
Ty ett verk hade Herren, HERREN Sebaot, att utföra i kaldéernas land.
Ja, kommen över det från alla sidor, öppnen dess förrådskammare, kasten i en hög vad där finnes, såsom man gör med säd, och given det till spillo; låten intet därav bliva kvar.
Nedgören alla dess tjurar, fören dem ned till att slaktas.
Ve dem, ty deras dag har kommit, deras hemsökelses tid!
Hör huru de fly och söka rädda sig ur Babels land, för att i Sion förkunna HERRENS, vår Guds, hämnd, hämnden för hans tempel.
Båden upp mot Babel folk i mängd, allt vad bågskyttar heter; lägren eder runt omkring det, låten ingen undkomma.
Vedergällen det efter dess gärningar; gören mot det alldeles såsom det självt har gjort.
Ty mot HERREN har det handlat övermodigt, mot Israels Helige.
Därför skola dess unga man falla på dess gator, och alla dess stridsmän skola förgöras på den dagen, säger HERREN.
Se, jag skall vända mig mot dig, du övermodige, säger Herren, HERREN Sebaot, ty din dag har kommit, den tid då jag vill hemsöka dig.
Då skall den övermodige stappla och falla, och ingen skall kunna upprätta honom.
Och jag skall tända eld på hans städer, och elden skall förtära allt omkring honom.
Så säger HERREN Sebaot: Förtryckta äro Israels barn, och Juda barn jämte dem.
Alla de som hava fart dem i fångenskap hålla dem fast och vilja icke släppa dem.
Men deras förlossare är stark; HERREN Sebaot är hans namn.
Han skall förvisso utföras deras sak, så att han skaffar ro åt jorden -- men oro åt Babels invånare.
Svärd komme över kaldéerna, säger HERREN, över Babels invånare, över dess furstar och dess visa män!
Svärd komme över lögnprofeterna, så att de stå där såsom dårar!
Svärd komme över dess hjältar, så att de bliva förfärade!
Svärd komme över dess hästar och vagnar och över allt främmande folk därinne, så att de bliva såsom kvinnor!
Svärd komme över dess skatter, så att de bliva tagna såsom byte!
Torka komme över dess vatten, så att de bliva uttorkade!
Ty det är ett belätenas land, och skräckgudar dyrka de såsom vanvettiga människor.
Därför skola nu schakaler bo där tillsammans med andra ökendjur, och strutsar skola där få sin boning.
Aldrig mer skall det bliva bebyggt, från släkte till släkte skall det vara obebott.
Likasom när Sodom och Gomorra med sina grannstäder omstörtades av Gud, säger HERREN, så skall ingen mer bo där och intet människobarn där vistas.
Se, ett folk kommer norrifrån; ett stort folk och många konungar resa sig och komma från jordens yttersta ända.
De föra båge och lans, de äro grymma och utan förbarmande.
Dånet av dem är såsom havets brus, och på sina hästar rida de fram, rustade såsom kämpar till strid, mot dig, du dotter Babel.
När konungen i Babel hör ryktet om dem, sjunka hans händer ned; ängslan griper honom, ångest lik en barnaföderskas.
Se, lik ett lejon som drager upp från Jordanbygdens snår och bryter in på frodiga betesmarker skall jag i ett ögonblick jaga dem bort därifrån; och den som jag utväljer skall jag sätta till herde över dem.
Ty vem är min like, och vem kan ställa mig till ansvar?
Och vilken är den herde som kan bestå inför mig?
Hören därför det råd som HERREN har lagt mot Babel, och de tankar som han har mot kaldéernas land: Ja, herdegossarna skola sannerligen släpas bort; sannerligen, deras betesmark skall häpna över dem.
När man ropar: »Babel är intaget», då bävar jorden, och ett skriande höres bland folken.
Så säger HERREN: Se, jag skall uppväcka mot Babel och mot Leb-Kamais inbyggare en fördärvares ande.
Och jag skall sända främlingar mot Babel, och de skola kasta det med kastskovlar och ödelägga dess land.
Ja, från alla sidor skola de komma emot det på olyckans dag.
Skyttar skola spänna sina bågar mot dem som där spänna båge, och mot dem som där yvas i pansar.
Skonen icke dess unga män, given hela dess här till spillo.
Dödsslagna män skola då falla i kaldéernas land och genomborrade man på dess gator.
Ty Israel och Juda äro icke änkor som hava blivit övergivna av sin Gud, av HERREN Sebaot, därför att deras land var fullt av skuld mot Israels Helige.
Flyn ut ur Babel; må var och en söka rädda sitt liv, så att I icke förgås genom dess missgärning.
Ty detta är för HERREN en hämndens tid, då han vill vedergälla det vad det har gjort.
Babel var i HERRENS hand en gyllene kalk som gjorde hela jorden drucken.
Av dess vin drucko folken, och så blevo folken såsom vanvettiga.
Men plötsligt är nu Babel fallet och krossat.
Jämren eder över henne, hämten balsam för hennes plåga, om hon till äventyrs kan helas.
»Ja, vi hava sökt hela Babel, men hon har icke kunnat helas; låt oss lämna henne och gå var och en till sitt land.
Ty hennes straffdom räcker upp till himmelen och når allt upp till skyarna.
HERREN har låtit vår rätt gå fram; kom, låt oss förtälja i Sion HERRENS, vår Guds, verk.»
Vässen pilarna, fatten sköldarna.
HERREN har uppväckt de mediska konungarnas ande; ty hans tankar äro vända mot Babel till att fördärva det.
Ja, HERRENS hämnd är här, hämnden för hans tempel.
Resen upp ett baner mot Babels murar, hållen sträng vakt, ställen ut väktare, läggen bakhåll; ty HERREN har fattat sitt beslut, och han gör vad han har talat mot Babels invånare.
Du som bor vid stora vatten och är så rik på skatter, din ände har nu kommit, din vinningslystnads mått är fyllt.
HERREN Sebaot har svurit vid sig själv: sannerligen, om jag än har uppfyllt dig med människor så talrika som gräshoppor, så skall man dock få upphäva skördeskri över dig.
Han har gjort jorden genom sin kraft, han har berett jordens krets genom sin vishet, och genom sitt förstånd har han utspänt himmelen.
När han vill låta höra sin röst, då brusa himmelens vatten, då låter han regnskyar stiga upp från jordens ända; han låter ljungeldar komma med regn och för vinden ut ur dess förvaringsrum.
Såsom dårar stå då alla människor där och begripa intet; guldsmederna komma då alla på skam med sina beläten, ty deras gjutna beläten äro lögn, och ingen ande är i dem.
De äro fåfänglighet, en tillverkning att le åt; när hemsökelsen kommer över dem, måste de förgås.
Men sådan är icke han som är Jakobs del; nej, det är han som har skapat allt, och särskilt sin arvedels stam.
HERREN Sebaot är hans namn.
Du var min hammare, mitt stridsvapen; med dig krossade jag folk, med dig fördärvade jag riken.
Med dig krossade jag häst och ryttare; med dig krossade jag vagn och körsven.
Med dig krossade jag man och kvinna; med dig krossade jag gammal och ung; med dig krossade jag yngling och jungfru.
Med dig krossade jag herden och hans hjord; med dig krossade jag åkermannen och hans oxpar; med dig krossade jag ståthållare och landshövding.
Men nu skall jag vedergälla Babel och alla Kaldeens inbyggare allt det onda som de hava förövat mot Sion, inför edra ögon, säger HERREN.
Se, jag skall vända mig mot dig, du fördärvets berg, säger HERREN, du som fördärvade hela jorden; och jag skall uträcka min hand mot dig och vältra dig ned från klipporna och göra dig till ett förbränt berg,
så att man icke av dig skall kunna taga vare sig hörnsten eller grundsten, utan du skall bliva en ödemark för evärdlig tid, säger HERREN.
Resen upp ett baner på jorden, stöten i basun ibland folken, invigen folk till strid mot det, båden upp mot det riken, både Ararats, Minnis och Askenas', tillsätten hövdingar mot det, dragen ditupp med hästar som likna borstiga gräshoppor.
Invigen folk till strid mot det: Mediens konungar, dess ståthållare och alla dess landshövdingar, och hela det land som lyder under deras välde.
Då darrar jorden och bävar, ty nu fullbordas vad HERREN tänkte mot Babel: att han ville göra Babels land till en ödemark, där ingen skulle bo.
Babels hjältar upphöra att strida, de sitta stilla i sina fästen; deras styrka har försvunnit, de hava blivit såsom kvinnor.
Man har tänt eld på dess boningar; dess bommar äro sönderbrutna.
Löparna löpa mot varandra, den ene budbäraren korsar den andres väg, med bud till konungen i Babel om att hela hans stad år intagen,
att vadställena äro besatta och dammarna förbrända i eld och krigsmännen gripna av skräck.
Ty så säger HERREN Sebaot, Israels Gud: Dottern Babel är såsom en tröskplats, när man just har trampat till den; ännu en liten tid, och skördetiden kommer för henne.
Uppätit mig och förgjort mig har han, Nebukadressar, konungen i Babel.
Han har gjort mig till ett tomt kärl; lik en drake har han uppslukat mig, han har fyllt sin buk med mina läckerheter och drivit mig bort.
»Den orätt mig har skett och det som har vederfarits mitt kött, det komme över Babel», så må Sions invånare säga; och »Mitt blod komme över Kaldeens inbyggare», så må Jerusalem säga.
Därför säger HERREN så: Se, jag skall utföra din sak och utkräva din hämnd.
Jag skall låta dess hav sina bort och dess brunn uttorka,
och Babel skall bliva en stenhop, en boning för schakaler, ett föremål för häpnad och begabberi, så att ingen kan bo där.
Alla ryta de nu såsom lejon; de skria såsom lejonungar.
Men när de äro som mest upptända, skall jag tillreda åt dem ett gästabud; jag skall göra dem druckna, så att de jubla.
Så skola de somna in i en evig sömn, ur vilken de aldrig skola uppvakna, säger HERREN.
Jag skall föra dem ned till att slaktas såsom lamm, likasom vädurar och bockar.
Huru har icke Sesak blivit intaget och hon som var hela jordens berömmelse erövrad!
Huru har icke Babel blivit ett föremål för häpnad bland folken!
Havet steg upp över Babel; av dess brusande böljor blev det övertäckt.
Så blev av dess städer en ödemark, ett torrt land och en hedmark, ett land där ingen bor, och där intet människobarn går fram.
Ja, jag skall hemsöka Bel i Babel och taga ut ur hans gap vad han har slukat; och folken skola icke mer strömma till honom.
Babels murar skola ock falla.
Dragen ut därifrån, mitt folk; må var och en söka rädda sitt liv undan HERRENS vredes glöd.
Varen icke försagda i edra hjärtan, och frukten icke för de olycksbud som höras i landet, om än ett olycksbud kommer det ena året och sedan nästa år ett nytt olycksbud, och om än våld råder på jorden och härskare står mot härskare.
Se, därför skola dagar komma, då jag skall hemsöka Babels beläten, och då hela dess land skall stå med skam och alla skola falla slagna därinne.
Då skola himmel och jord jubla över Babel, de och allt vad i dem är, då nu förhärjarna komma över det norrifrån, säger HERREN.
Ja, I slagna av Israel, också Babel måste falla, likasom för Babel människor föllo slagna över hela jorden.
I som haven lyckats rädda eder undan svärdet, gån åstad, stannen icke.
Kommen ihåg HERREN, i fjärran land, och tänken på Jerusalem.
Vi stå här med skam, ja vi måste höra smädelse; blygsel höljer vårt ansikte, ty främlingar hava kastat sig över vad heligt som fanns i HERRENS hus.
Se, därför skola dagar komma, säger HERREN, då jag skall hemsöka dess beläten, och då slagna män skola jämra sig i hela dess land.
Om Babel än stege upp till himmelen, och om det gjorde sin befästning än så hög och stark så skulle dock förhärjare ifrån mig komma över det, säger HERREN.
Klagorop höras från Babel, och stort brak från kaldéernas land.
Ty HERREN förhärjar Babel och gör slut på det stora larmet därinne.
Och deras böljor brusa såsom stora vatten; dånet av dem ljuder högt.
Ty över det, över Babel, kommer en förhärjare, och dess hjältar tagas till fånga, deras bågar brytas sönder.
Se, HERREN är en vedergällningens Gud; han lönar till fullo.
Ja, jag skall göra dess furstar druckna, så ock dess visa män, dess ståthållare, dess landshövdingar och dess hjältar, och de skola somna in i en evig sömn, ur vilken de aldrig skola uppvakna, säger konungen, han vilkens namn är HERREN Sebaot.
Så säger HERREN Sebaot: Det vida Babels murar skola i grund omstörtas, och dess höga portar skola brännas upp i eld.
Så möda sig folken för det som skall bliva till intet, och folkslagen arbeta sig trötta för det som skall förbrännas av elden.
Detta är vad profeten Jeremia bjöd Seraja, son till Neria, son till Mahaseja, när denne begav sig till Babel med Sidkia, Juda konung, i hans fjärde regeringsår.
Seraja var nämligen den som hade bestyret med lägerplatserna.
Och Jeremia tecknade i en och samma bok upp alla de olyckor som skulle komma över Babel, allt detta som nu är skrivet om Babel.
Jeremia sade till Seraja: »När du kommer till Babel, så se till, att du läser upp allt detta.
Och du skall säga: 'HERRE, du har själv talat om denna ort att du vill fördärva den, så att ingen mer skall bo där, varken någon människa eller något djur; ty den skall vara en ödemark för evärdlig tid.'
Och när du har läst upp boken till slut, så bind en sten vid den och kasta den ut i Frat,
och säg: 'På detta sätt skall Babel sjunka ned och icke mer komma upp, för den olyckas skull som jag skall låta komma över det, mitt under deras ävlan.'»
Så långt Jeremias ord.
Sidkia var tjuguett år gammal, när han blev konung, och han regerade elva år i Jerusalem.
Hans moder hette Hamital, Jeremias dotter, från Libna.
Han gjorde vad ont var i HERRENS ögon, alldeles såsom Jojakim hade gjort.
Ty på grund av HERRENS vrede skedde vad som skedde med Jerusalem och Juda, till dess att han kastade dem bort ifrån sitt ansikte.
Och Sidkia avföll från konungen i Babel.
Då, i hans nionde regeringsår, i tionde månaden, på tionde dagen i månaden, kom Nebukadressar, konungen i Babel, med hela sin här till Jerusalem, och de belägrade det; och de byggde en belägringsmur runt omkring det.
Så blev staden belägrad och förblev så ända till konung Sidkias elfte regeringsår.
Men i fjärde månaden, på nionde dagen i månaden, var hungersnöden så stor i staden, att mängden av folket icke hade något att äta.
Och staden stormades, och allt krigsfolket flydde och drog ut ur staden om natten genom porten mellan de båda murarna (den port som ledde till den kungliga trädgården), medan kaldéerna lågo runt omkring staden; och de togo vägen åt Hedmarken till.
Men kaldéernas här förföljde konungen, och de hunno upp Sidkia på Jerikos hedmarker, sedan hela hans här hade övergivit honom och skingrat sig.
Och de grepo konungen och förde honom till den babyloniske konungen i Ribla i Hamats land; där höll denne rannsakning och dom med honom.
Och konungen i Babel lät slakta Sidkias barn inför hans ögon; därjämte lät han ock slakta alla Juda furstar i Ribla.
Och på Sidkia själv lät han sticka ut ögonen och lät fängsla honom med kopparfjättrar.
Och konungen i Babel förde honom därefter till Babel och lät honom sitta i fängelsehuset ända till hans dödsdag.
I femte månaden, på tionde dagen i månaden, detta i den babyloniske konungen Nebukadressars nittonde regeringsår, kom Nebusaradan, översten för drabanterna; denne var den babyloniske konungens förtroendeman vid Jerusalem.
Han brände upp HERRENS hus och konungshuset; ja, alla hus i Jerusalem, i synnerhet alla de förnämas hus, brände han upp i eld.
Och alla murar runt omkring Jerusalem brötos ned av hela den här av kaldéer, som översten för drabanterna hade med sig.
Och en del av de ringaste bland folket och den övriga återstoden av folket, dem som voro kvar i staden, och de överlöpare som hade gått över till konungen i Babel, så ock det hantverksfolk som fanns kvar, dem förde Nebusaradan, översten för drabanterna, bort i fångenskap.
Men av de ringaste i landet lämnade Nebusaradan, översten för drabanterna, några kvar till vingårdsmän och åkermän.
Kopparpelarna i HERRENS hus, bäckenställen och kopparhavet i HERRENS hus slogo kaldéerna sönder och förde all kopparen till Babel.
Och askkärlen, skovlarna, knivarna, de båda slagen av skålar och alla kopparkärl som hade begagnats vid gudstjänsten togo de bort.
Likaledes tog översten för drabanterna bort faten, fyrfaten, offerskålarna, askkärlen, ljusstakarna, de andra skålarna och bägarna, allt vad som var av rent guld eller av rent silver.
Vad angår de två pelarna, havet som var allenast ett, och de tolv kopparoxarna under bäckenställen, som konung Salomo hade låtit göra till HERRENS hus, så kunde kopparen i alla dessa föremål icke vägas.
Och vad pelarna angår, så var den ena pelaren aderton alnar hög, och en tolv alnar lång tråd mätte dess omfång, och den var fyra finger tjock och ihålig.
Och ovanpå den var ett pelarhuvud av koppar; och detta ena pelarhuvud var fem alnar högt, och ett nätverk och granatäpplen funnos på pelarhuvudet runt omkring, alltsammans av koppar.
Och likadant var det på den andra pelaren med fina granatäpplen.
Och granatäpplena voro nittiosex utåt; men tillsammans voro granatäpplena på nätverket runt omkring ett hundra.
Och översten för drabanterna tog översteprästen Seraja jämte Sefanja prästen näst under honom, så ock de tre som höllo vakt vid tröskeln,
och från staden tog han en hovman, den som var anförare för krigsfolket, och sju av konungens närmaste män, som påträffades i staden, så ock härhövitsmannens sekreterare, som plägade utskriva folket i landet till krigstjänst, och sextio andra män av landets folk, som påträffades i staden --
dessa tog Nebusaradan, översten för drabanterna, och förde dem till den babyloniske konungen i Ribla.
Och konungen i Babel lät avliva dem där, i Ribla i Hamats land.
Så blev Juda bortfört från sitt land.
Detta är antalet av dem som Nebukadressar förde bort: i det sjunde året tre tusen tjugutre judar,
och i Nebukadressars adertonde: regeringsår åtta hundra trettiotvå personer från Jerusalem.
Men i Nebukadressars tjugutredje regeringsår bortförde Nebusaradan, översten för drabanterna, av judarna sju hundra fyrtiofem personer.
Hela antalet utgjorde fyra tusen sex hundra personer.
Men i det trettiosjunde året sedan Jojakin, Juda konung, hade blivit bortförd i fångenskap, i tolfte månaden, på tjugufemte dagen i månaden, tog Evil-Merodak, konungen i Babel -- samma år han blev konung -- Jojakin, Juda konung, till nåder och förde honom ut ur fängelset.
Och han talade vänligt med honom och gav honom översta platsen bland de konungar som voro hos honom i Babel.
Han fick lägga av sin fångdräkt och beständigt äta vid hans bord, så länge han levde.
Och ett ständigt underhåll gavs honom från konungen i Babel, visst för var dag, ända till hans dödsdag, så länge han levde.
Huru övergiven sitter hon icke, den folkrika staden!
Hon har blivit lik en änka.
Hon som var så mäktig bland folken, en furstinna bland länderna, hon måste nu göra trältjänst.
Bittert gråter hon i natten, och tårar rinna utför hennes kind.
Ingen finnes, som tröstar henne, bland alla hennes vänner.
Alla hennes närmaste hava varit trolösa mot henne; de hava blivit hennes fiender.
Juda har måst gå i landsflykt efter att hava utstått elände och svåra vedermödor; hon bor nu bland hedningarna och finner ingen ro.
Alla hennes förföljare hava fallit över henne, mitt i hennes trångmål.
Vägarna till Sion ligga sörjande, då nu ingen kommer till högtiderna.
Alla hennes portar äro öde, hennes präster sucka.
Hennes jungfrur äro bedrövade, och själv sörjer hon bittert.
Hennes ovänner hava fått övermakten, för hennes fiender går allt väl.
Ty HERREN har sänt henne bedrövelser för hennes många överträdelsers skull.
Hennes barn hava måst gå i fångenskap, bortdrivna av ovännen.
Så har all dottern Sions härlighet försvunnit ifrån henne.
Hennes furstar likna hjortar som icke finna något bete; vanmäktiga söka de fly bort, undan sina förföljare.
I denna sitt eländes och sin husvillhets tid kommer Jerusalem ihåg allt vad dyrbart hon ägde i forna dagar.
Nu då hennes folk har fallit för ovännens hand och hon icke har någon hjälpare nu se hennes ovänner med hån på hennes undergång.
Svårt hade Jerusalem försynda sig; därför har hon blivit en styggelse.
Alla som ärade henne förakta henne nu, då de se hennes blygd.
Därför suckar hon ock själv och drager sig undan.
Orenhet fläckar hennes klädesfållar; hon tänkte icke på anden.
Därför vart hennes fall så gruvligt; ingen finnes, som tröstar henne.
Se, HERRE, till mitt elände, ty fienden förhäver sig.
Ovännen räckte ut sin hand efter allt vad dyrbart hon ägde; ja, hon fick se huru hedningar kommo in i hennes helgedom, just sådana som du hade förbjudit att komma in i din församling.
Allt hennes folk måste med suckan tigga sitt bröd; för vad dyrbart de ägde måste de köpa sig mat till att stilla sin hunger.
Se, HERRE, och akta på huru föraktad jag har blivit.
Går detta eder ej till sinnes, I alla som dragen vägen fram?
Akten härpå och sen till: kan någon plåga vara lik den varmed jag har blivit hemsökt, den varmed HERREN har bedrövat mig på sin glödande vredes dag?
Från höjden sände han en eld i mina ben och fördärvade dem.
Han bredde ut ett nät för mina fötter, han stötte mig tillbaka.
Förödelse lät han gå över mig, han gjorde mig maktlös för alltid.
Mina överträdelser knötos samman av hans hand till ett ok, hopbundna lades de på min hals; så bröt han ned min kraft.
Herren gav mig i händerna på människor som jag ej kan stå emot.
Alla de tappra kämpar jag hyste aktade Herren för intet.
Han lyste ut högtid, mig till fördärv, för att krossa mina unga män.
Ja, vinpressen trampade Herren till ofärd för jungfrun dottern Juda.
Fördenskull gråter jag; mitt öga, det flyter i tårar; ty fjärran ifrån mig äro de som skulle trösta mig och vederkvicka min själ.
Förödelse har gått över mina barn, ty fienden har blivit mig övermäktig.
Sion räcker ut sina händer, men ingen finnes, som tröstar henne; mot Jakob bådade HERREN upp ovänner från alla sidor; Jerusalem har blivit en styggelse ibland dem.
Ja, HERREN är rättfärdig, ty jag var gensträvig mot hans bud.
Hören då, alla I folk, och sen min plåga: mina jungfrur och mina unga män fingo gå i fångenskap.
Jag kallade på mina vänner, men de bedrogo mig.
Mina präster och mina äldste förgingos i staden, medan de tiggde sig mat för att stilla sin hunger.
Se HERRE, huru jag är i nöd, mitt innersta är upprört.
Mitt hjärta vänder sig i mitt bröst, därför att jag var så gensträvig.
Ute har svärdet förgjort mina barn, och inomhus pesten.
Väl hör man huru jag suckar, men ingen finnes, som tröstar mig; alla mina fiender höra om min olycka och fröjda sig över att du har gjort detta.
Den dag du förkunnade har du låtit komma.
Dock, dem skall det gå såsom mig.
Låt all deras ondska komma inför ditt ansikte, och hemsök dem, likasom du har hemsökt mig för alla mina överträdelsers skull ty många äro mina suckar, och mitt hjärta är sjukt.
Huru höljer icke Herren genom sin vrede dottern Sion i mörker!
Från himmelen ned till jorden kastade han Israels härlighet.
Han vårdade sig icke om sin fotapall på sin vredes dag.
Utan skonsamhet fördärvade Herren alla Jakobs boningar; i sin förgrymmelse bröt han ned dottern Judas fästen, ja, han slog dem till jorden, han oskärade riket och dess furstar.
I sin vredes glöd högg han av vart Israels horn; han höll sin högra hand tillbaka, när fienden kom.
Jakob förbrände han lik en lågande eld, som förtär allt runt omkring.
Han spände sin båge såsom en fiende, med sin högra hand stod han fram såsom en ovän och dräpte alla som voro våra ögons lust.
Över dottern Sions hydda utgöt han sin vrede såsom en eld.
Herren kom såsom en fiende och fördärvade Israel, han fördärvade alla dess palats, han förstörde dess fästen; så hopade han över dottern Juda jämmer på jämmer.
Och han bröt ned sin hydda såsom en trädgård, han förstörde sin högtidsplats.
Både högtid och sabbat lät HERREN bliva förgätna i Sion, och i sin vredes förgrymmelse försköt han både konung och präst.
Herren förkastade sitt altare, han gav sin helgedom till spillo.
Murarna omkring hennes palatser gav han i fiendernas hand.
De hovo upp rop i HERRENS hus såsom på en högtidsdag.
HERREN hade beslutit att förstöra dottern Sions murar; han spände mätsnöret till att fördärva och drog sin hand ej tillbaka.
Han lät sorg komma över vallar och murar; förfallna ligga de nu alla.
Hennes portar sjönko ned i jorden, han bräckte och krossade hennes bommar.
Hennes konung och furstar leva bland hedningar, ingen lag finnes mer; hennes profeter undfå ej heller någon syn från HERREN.
Dottern Sions äldste sitta där stumma på jorden, de hava strött stoft på sina huvuden och höljt sig i sorgdräkt; Jerusalems jungfrur sänka sina huvuden mot jorden.
Mina ögon äro förtärda av gråt, mitt innersta är upprört, min lever är såsom utgjuten på jorden för dottern mitt folks skada; ty barn och spenabarn försmäkta på gatorna i staden.
De ropa till sina mödrar: »Var få vi bröd och vin?»
Ty försmäktande ligga de såsom slagna på gatorna i staden; ja, de uppgiva sin anda i sina mödrars famn.
Vad jämförligt skall jag framlägga för dig, du dotter Jerusalem?
Vilket liknande öde kan jag draga fram till din tröst, du jungfru dotter Sion?
Din skada är ju stor såsom ett hav; vem kan hela dig?
Dina profeters syner voro falskhet och flärd, de blottade icke för dig din missgärning, så att du kunde bliva upprättad; de utsagor de förkunnade för dig voro falskhet och förförelse.
Alla vägfarande slå ihop händerna, dig till hån; de vissla och skaka huvudet åt dottern Jerusalem: »Är detta den stad som man kallade 'skönhetens fullhet', 'hela jordens fröjd'?»
Alla dina fiender spärra upp munnen emot dig, de vissla och bita samman tänderna, de säga: »Vi hava fördärvat henne.
Ja, detta är den dag som vi bidade efter; nu hava vi upplevat och sett den.»
HERREN har gjort vad han hade beslutit, han har fullbordat sitt ord, vad han för länge sedan hade förordnat; han har brutit ned utan förskoning.
Och han har låtit fienden glädjas över dig, han har upphöjt dina ovänners horn.
Deras hjärtan ropa till Herren.
Du dottern Sions mur, låt dina tårar rinna som en bäck, både dag och natt; låt dig icke förtröttas, unna ditt öga ingen ro.
Stå upp, ropa högt i natten, när dess väkter begynna, utgjut ditt hjärta såsom vatten inför Herrens ansikte; lyft upp till honom dina händer för dina barns liv, ty de försmäkta av hunger i alla gators hörn.
Se, HERRE, och akta på vem du så har hemsökt.
Skola då kvinnor nödgas äta sin livsfrukt, barnen som de hava burit i sin famn?
Skall man i Herrens helgedom dräpa präster och profeter?
På jorden, ute på gatorna, ligga de, både unga och gamla; mina jungfrur och mina unga män hava fallit för svärd.
Du dräpte på din vredes dag, du slaktade utan förskoning.
Såsom till en högtidsdag kallade du samman mot mig förskräckelser ifrån alla sidor; och på HERRENS vredes dag fanns ingen som blev räddad och slapp undan.
Dem som jag hade burit i min famn och fostrat, dem förgjorde min fiende.
Jag är en man som har prövat elände under hans vredes ris.
Mig har han fört och låtit vandra genom mörker och genom ljus.
Ja, mot mig vänder han sin hand beständigt, åter och åter.
Han har uppfrätt mitt kött och min hud, han har krossat benen i mig.
Han har kringskansat och omvärvt mig med gift och vedermöda.
I mörker har han lagt mig såsom de längesedan döda.
Han har kringmurat mig, så att jag ej kommer ut, han har lagt på mig tunga fjättrar.
Huru jag än klagar och ropar, tillstoppar han öronen för min bön.
Med huggen sten har han murat för mina vägar, mina stigar har han gjort svåra.
En lurande björn är han mot mig, ett lejon som ligger i försåt.
Han förde mig på villoväg och rev mig i stycken, förödelse lät han gå över mig.
Han spände sin båge och satte mig upp till ett mål för sin pil.
Ja, pilar från sitt koger sände han in i mina njurar.
Jag blev ett åtlöje för hela mitt folk en visa för dem hela dagen.
Han mättade mig med bittra örter, han gav mig malört att dricka.
Han lät mina tänder bita sönder sig på stenar, han höljde mig med aska.
Ja, du förkastade min själ och tog bort min frid; jag visste ej mer vad lycka var.
Jag sade: »Det är ute med min livskraft och med mitt hopp till HERREN.»
Tänk på mitt elände och min husvillhet, på malörten och giftet!
Stadigt tänker min själ därpå och är bedrövad i mig.
Men detta vill jag besinna, och därför skall jag hoppas:
HERRENS nåd är det att det icke är ute med oss, ty det är icke slut med hans barmhärtighet.
Den är var morgon ny, ja, stor är din trofasthet.
HERREN är min del, det säger min själ mig; därför vill jag hoppas på honom.
HERREN är god mot dem som förbida honom, mot den själ som söker honom.
Det är gott att hoppas i stillhet på hjälp från HERREN.
Det är gott för en man att han får bära ett ok i sin ungdom.
Må han sitta ensam och tyst, när ett sådant pålägges honom.
Må han sänka sin mun i stoftet; kanhända finnes ännu hopp.
Må han vända kinden till åt den som slår honom och låta mätta sig med smälek.
Ty Herren förkastar icke för evig tid;
utan om han har bedrövat, så förbarmar han sig igen, efter sin stora nåd.
Ty icke av villigt hjärta plågar han människors barn och vållar dem bedrövelse.
Att man krossar under sina fötter alla fångar i landet,
att man vränger en mans rätt inför den Högstes ansikte,
att man gör orätt mot en människa i någon hennes sak, skulle Herren icke se det?
Vem sade, och det vart, om det ej var Herren som bjöd?
Kommer icke från den Högstes mun både ont och gott?
Varför knorrar då en människa här i livet, varför en man, om han drabbas av sin synd?
Låtom oss rannsaka våra vägar och pröva dem och omvända oss till HERREN.
Låtom oss upplyfta våra hjärtan, såväl som våra händer, till Gud i himmelen.
Vi hava varit avfälliga och gensträviga, och du har icke förlåtit det.
Du har höljt dig i vrede och förföljt oss, du har dräpt utan förskoning.
Du har höljt dig i moln, så att ingen bön har nått fram.
Ja, orena och föraktade låter du oss stå mitt ibland folken.
Alla våra fiender spärra upp munnen emot oss.
Faror och fallgropar möta oss fördärv och skada.
Vattenbäckar rinna ned från mitt öga för dottern mitt folks skada.
Mitt öga flödar utan uppehåll och förtröttas icke,
till dess att HERREN blickar ned från himmelen och ser härtill.
Mitt öga vållar mig plåga för alla min stads döttrars skull.
Jag bliver ivrigt jagad såsom en fågel av dem som utan sak äro mina fiender.
De vilja förgöra mitt liv här i djupet, de kasta stenar på mig.
Vatten strömma över mitt huvud, jag säger: »Det är ute med mig.»
Jag åkallar ditt namn, o HERRE, har underst i djupet.
Du hör min röst; tillslut icke ditt öra, bered mig lindring, då jag nu ropar.
Ja, du nalkas mig, när jag åkallar dig; du säger: »Frukta icke.»
Du utför, Herre, min själs sak, du förlossar mitt liv.
Du ser, HERRE, den orätt mig vederfares; skaffa mig rätt.
Du ser all deras hämndgirighet, alla deras anslag mot mig.
Du hör deras smädelser, HERRE, alla deras anslag mot mig.
Vad mina motståndare tala och tänka ut är beständigt riktat mot mig.
Akta på huru de hava mig till sin visa, evad de sitta eller stå upp.
Du skall giva dem vedergällning, HERRE, efter deras händers verk.
Du skall lägga ett täckelse över deras hjärtan; din förbannelse skall komma över dem.
Du skall förfölja dem i vrede och förgöra dem, så att de ej bestå under HERRENS himmel.
Huru har icke guldet berövats sin glans, den ädla metallen förvandlats!
Heliga stenar ligga kringkastade i alla gators hörn.
Sions ädlaste söner som aktades lika med fint guld, huru räknas de icke nu såsom lerkärl, krukmakarhänders verk!
Själva schakalerna räcka spenarna åt sina ungar för att giva dem di; men dottern mitt folk har blivit grym, lik strutsen i öknen.
Spenabarnets tunga låder av törst vid dess gom; le späda barnen bedja om bröd, men ingen bryter sådant åt dem.
De som förr åto läckerheter försmäkta nu på gatorna; de som uppföddes i scharlakan måste nu ligga i dyn.
Så var dottern mitt folks missgärning större än Sodoms synd, Sodoms, som omstörtades i ett ögonblick, utan att människohänder kommo därvid.
Hennes furstar voro mer glänsande än snö, de voro vitare än mjölk, deras hy var rödare än korall, deras utseende var likt safirens.
Nu hava deras ansikten blivit mörkare än svart färg, man känner icke igen dem på gatorna; deras hud sitter fastklibbad vid benen, den har förtorkats och blivit såsom trä.
Lyckligare voro de som dräptes med svärd, än de äro, som dräpas av hunger, de som täras bort under kval, utan näring från marken.
Med egna händer måste ömsinta kvinnor koka sina barn för att hava dem till föda vid dottern mitt folks skada.
HERREN har uttömt sin förtörnelse, utgjutit sin vredes glöd; i Sion har han tänt upp en eld, som har förtärt dess grundvalar.
Ingen konung på jorden hade trott det, ingen som bor på jordens krets, att någon ovän eller fiende skulle komma in genom Jerusalems portar.
För dess profeters synders skull har så skett, för dess prästers missgärningar, därför att de därinne utgöto de rättfärdigas blod.
Såsom blinda irra de omkring på gatorna, fläckade av blod. så att ingen finnes, som vågar komma vid deras kläder.
»Viken undan!» »Oren!», så ropar man framför dem; »Viken undan, viken undan, kommen icke vid den!» ja, flyktiga och ostadiga måste de vara; bland hedningarna säger man om dem: »De skola ej mer finna någon boning.»
HERRENS åsyn förskingrar dem, han vill icke mer akta på dem; mot prästerna visas intet undseende, mot de äldste ingen misskund.
Ännu försmäkta våra ögon i fåfäng väntan efter hjälp; från vårt vårdtorn speja vi efter ett folk som ändå ej kan frälsa oss.
Han lurar på vara steg, så att vi ej våga gå på våra gator.
Vår ände är nära, vara dagar äro ute; ja, vår ande har kommit.
Våra förföljare voro snabbare än himmelens örnar; på bergen jagade de oss, i öknen lade de försåt för oss.
HERRENS smorde, han som var vår livsfläkt, blev fångad i deras gropar, han under vilkens skugga vi hoppades att få leva bland folken.
Ja, fröjda dig och var glad, du dotter Edom, du som bor i Us' land!
Också till dig skall kalken komma; du skall varda drucken och få ligga blottad.
Din missgärning är ej mer, du dotter Sion; han skall ej åter föra dig bort i fångenskap.
Men din missgärning, du dotter Edom, skall han hemsöka; han skall uppenbara dina synder.
Tänk, HERRE, på vad som har vederfarits oss skåda ned och se till vår smälek.
Vår arvedel har kommit i främlingars ägo, våra hus i utlänningars.
Vi hava blivit värnlösa, vi hava ingen fader; våra mödrar äro såsom änkor.
Vattnet som tillhör oss få vi dricka allenast för penningar; vår egen ved måste vi betala.
Våra förföljare äro oss på halsen; huru trötta vi än äro, unnas oss dock ingen vila.
Vi hava måst giva oss under Egypten, under Assyrien, för att få bröd till att mätta oss med.
Våra fäder hava syndat, de äro icke mer, vi måste bära deras missgärningar.
Trälar få råda över oss; ingen finnes, som rycker oss ur deras våld.
Med fara för vårt liv hämta vi vårt bröd, bärga det undan öknens svärd.
Vår hud är glödande såsom en ugn, för brännande hungers skull.
Kvinnorna kränkte man i Sion, jungfrurna i Juda städer.
Furstarna blevo upphängda av deras händer, för de äldste visade de ingen försyn.
Ynglingarna måste bära på kvarnstenar, och gossarna dignade under vedbördor.
De gamla sitta icke mer i porten, de unga hava upphört med sitt strängaspel.
Våra hjärtan hava icke mer någon fröjd i sorgelåt är vår dans förvandlad.
Kronan har fallit ifrån vårt huvud; ve oss, att vi syndade så!
Därför hava ock våra hjärtan blivit sjuka, därför äro våra ögon förmörkade,
för Sions bergs skull, som nu ligger öde, så att rävarna ströva omkring därpå.
Du, HERRE, tronar evinnerligen; din tron består från släkte till släkte.
Varför vill du för alltid förgäta oss, förkasta oss för beständigt?
Tag oss åter till dig, HERRE, så att vi få vända åter; förnya våra dagar, så att de bliva såsom fordom.
Eller har du alldeles förkastat oss?
Förtörnas du på oss så övermåttan?
I det trettionde året, på femte dagen i fjärde månaden, när jag var bland de fångna vid strömmen Kebar, öppnades himmelen, och jag såg en syn från Gud.
På femte dagen i månaden, när femte året gick, efter att konung Jojakin hade blivit bortförd i fångenskap,
kom HERRENS ord till prästen Hesekiel, Busis son, i kaldéernas land vid strömmen Kebar, och HERRENS hand kom där över honom.
Och jag fick se en stormvind komma norrifrån, ett stort moln med flammande eld, och ett sken omgav det; och mitt däri, mitt i elden, syntes något som var såsom glänsande malm.
Och mitt däri syntes något som liknade fyra väsenden, och dessa sågo ut på följande sätt: de liknade människor,
men vart väsende hade fyra ansikten, och vart och ett av dem hade fyra vingar,
och deras ben voro raka och deras fötter såsom fötterna på en kalv och de glimmade såsom glänsande koppar.
Och de hade människohänder under sina vingar på alla fyra sidorna.
Och med de fyras ansikten och vingar förhöll det sig så:
deras vingar slöto sig intill varandra; och när de gingo, behövde de icke vända sig, utan gingo alltid rakt fram.
Och deras ansikten liknade människoansikten, och alla fyra hade lejonansikten på högra sidan, och alla fyra hade tjuransikten på vänstra sidan, och alla fyra hade ock örnansikten.
Så var det med deras ansikten.
Och deras vingar voro utbredda upptill; vart väsende hade två vingar med vilka de slöto sig intill varandra, och två som betäckte deras kroppar.
Och de gingo alltid rakt fram; vart anden ville gå, dit gingo de, och när de gingo, behövde de icke vända sig.
Och väsendena voro till sitt utseende lika eldsglöd, som brunno likasom bloss, under det att elden for omkring mellan väsendena; och den gav ett sken ifrån sig, och ljungeldar foro ut ur elden.
Och väsendena hastade fram och tillbaka likasom blixtar.
När jag nu såg på väsendena, fick jag se ett hjul stå på jorden, invid väsendena, vid var och en av deras fyra framsidor.
Och det såg ut som om hjulen voro gjorda av något som liknade krysolit, och alla fyra voro likadana; och det såg vidare ut som om de voro så gjorda, att ett hjul var insatt i ett annat.
När de skulle gå, kunde de gå åt alla fyra sidorna, de behövde icke vända sig, när de gingo.
Och deras lötar voro höga och förskräckliga, och på alla fyra voro lötarna fullsatta med ögon runt omkring.
Och när väsendena gingo, gingo ock hjulen invid dem, och när väsendena lyfte sig upp över jorden lyfte sig ock hjulen.
Vart anden ville gå, dit gingo de, ja, varthelst anden ville gå; och hjulen lyfte sig jämte dem, ty väsendenas ande var i hjulen.
När väsendena gingo, gingo ock dessa; när de stodo stilla, stodo ock dessa stilla; när de lyfte sig upp över jorden, lyfte sig ock hjulen jämte dem, ty väsendenas ande var i hjulen.
Och över väsendenas huvuden syntes något som liknade ett himlafäste, till utseendet såsom underbar kristall, utspänt ovanpå deras huvuden.
Och under fästet voro deras vingar utbredda rätt emot varandra Vart särskilt väsende hade två vingar med vilka det kunde betäcka sin kropp.
Och när de gingo, lät dånet av deras vingar i mina öron såsom dånet av stora vatten, såsom den Allsmäktiges röst; ja, det var ett väldigt dån, likt dånet från en härskara.
Men när de stodo stilla, höllo de sina vingar nedsänkta.
Och ovan fästet, som vilade på deras huvuden, dånade det; när de då stodo stilla, höllo de sina vingar nedsänkta.
Och ovanpå fästet, som vilade på deras huvuden, syntes något som såg ut att vara av safirsten, och som liknade en tron; och ovanpå det som liknade en tron satt en som till utseendet liknade en människa,
Och jag såg något som var såsom glänsande malm och omgivet runt omkring av något som såg ut såsom eld, ända ifrån det som såg ut att vara hans länder och sedan allt uppåt.
Men nedåt från det som såg ut att vara hans länder såg jag något som såg ut såsom eld; och ett sken omgav honom.
Såsom bågen som synes i skyn, när det regnar, så såg skenet ut där runt omkring.
Så såg det ut, som tycktes mig vara HERRENS härlighet; och när jag såg det, föll jag ned på mitt ansikte, och jag hörde rösten av en som talade
Och han sade till mig: »Du människobarn, stå upp på dina fötter, så vill jag tala med dig.»
När han så talade till mig, kom en andekraft i mig och reste upp mig på mina fötter; och jag hörde på honom som talade till mig.
Och han sade till mig: »Du människobarn, jag sänder dig till Israels barn, de avfälliga hedningarna som hava avfallit från mig; de och deras fäder hava begått överträdelser mot mig allt intill den dag som i dag är.
Till barnen med hårda pannor och förstockade hjärtan sänder jag dig, och du skall säga till dem: 'Så säger Herren, HERREN'
Och evad de höra därpå eller icke -- ty de äro ett gensträvigt släkte -- så skola de dock förnimma att en profet har varit ibland dem.
Och du, människobarn, frukta icke för dem, och frukta icke för deras ord, fastän du omgives av tistlar och törnen och bor ibland skorpioner.
Nej, frukta icke för deras ord, och var icke förfärad för dem själva, då de nu äro ett gensträvigt släkte.
Utan tala mina ord till dem, evad de höra på dem eller icke, då de nu äro så gensträviga.
Men du, människobarn, hör nu vad jag talar till dig; var icke gensträvig såsom detta gensträviga släkte.
Öppna din mun och ät vad jag giver dig.»
Och jag fick se en hand uträckas mot mig, och i den såg jag en bokrulle.
Och denna breddes ut framför mig, och den var fullskriven innan och utan; och där voro uppskrivna klagosånger, suckan och verop.
Och han sade till mig: »Du människobarn, ät vad du här finner, ät upp denna rulle, och gå sedan åstad och tala till Israels hus.»
Då öppnade jag min mun, och han gav mig rullen att äta.
Och han sade till mig: »Du människobarn, du måste mätta din buk och fylla dina inälvor med den rulle som jag nu giver dig.»
Och jag åt, och den var i min mun söt såsom honung.
Och han sade till mig: »Du människobarn, gå bort till Israels hus och tala till dem med mina ord.
Ty du bliver ju icke sänd till ett folk med obegripligt språk och trög tunga, utan till Israels hus,
icke till mångahanda folk med obegripligt språk och trög tunga, vilkas tal du icke förstår; sannerligen, sände jag dig till sådana, så skulle de höra på dig
Men Israels hus vill icke höra på dig, ty de vilja icke höra på mig; hela Israels hus har hårda pannor och förhärdade hjärtan.
Men se, jag gör ditt ansikte hårt såsom deras ansikten, och din panna hård såsom deras pannor.
Ja, jag gör din panna hård såsom diamant, hårdare än flinta.
Du skall icke frukta för dem och icke förfäras för dem, då de nu äro ett gensträvigt släkte.»
Och han sade till mig: »Du människobarn, allt vad jag talar till dig skall du upptaga i ditt hjärta och höra med dina öron.
Och gå bort till dina fångna landsmän, och tala till dem och säg till dem: 'Så säger Herren, HERREN' -- evad de nu höra därpå eller icke.»
Och en andekraft lyfte upp mig, och jag hörde bakom mig ljudet av ett väldigt dån: »Lovad vare HERRENS härlighet, där varest den är!»,
så ock ljudet av väsendenas vingar, som rörde vid varandra, och ljudet av hjulen jämte dem och ljudet av ett väldigt dån.
Och en andekraft lyfte upp mig och förde mig bort, och jag färdades åstad, bedrövad och upprörd i min ande, och HERRENS hand var stark över mig.
Och jag kom till de fångna i Tel-Abib, till dem som bodde vid strömmen Kebar, till den plats där de bodde; och jag satt där ibland dem i sju dagar, försänkt i djup sorg.
Men efter sju dagar kom HERRENS ord till mig; han sade:
»Du människobarn, jag har satt dig till en väktare för Israels hus, för att du å mina vagnar skall varna dem, när du hör ett ord från min mun.
Om jag säger till den ogudaktige: 'Du måste dö' och du då icke varnar honom, ja, om du icke säger något till att varna den ogudaktige för hans ogudaktiga väg och rädda hans liv, då skall väl den ogudaktige dö genom sin missgärning, men hans blod skall jag utkräva av din hand.
Men om du varnar den ogudaktige och han likväl icke vänder om från sin ogudaktighet och sin ogudaktiga väg, då skall visserligen han dö genom sin missgärning, men du själv har räddat din själ.
Och om en rättfärdig man vänder om från sin rättfärdighet och gör vad orätt är, så skall jag lägga en stötesten i hans väg, och han skall dö.
Om du då icke har varnat honom, så skall han väl dö genom sin synd, och den rättfärdighet som han förr har övat skall icke varda ihågkommen, men hans blod skall jag utkräva av din hand.
Men om du har varnat den rättfärdige, för att han, den rättfärdige, icke skall synda, och han så avhåller sig från synd, då skall han förvisso få leva, därför att han lät varna sig, och du själv har då räddat din själ.»
Och HERRENS hand kom där över mig, och han sade till mig: »Stå upp och gå ut på slätten; där skall jag tala med dig.»
Då stod jag upp och gick ut på slätten; och se, där stod HERRENS härlighet, alldeles sådan som jag hade sett den vid strömmen Kebar; och jag föll ned på mitt ansikte.
Men en andekraft kom i mig och reste upp mig på mina fötter.
Och han talade med mig och sade till mig: »Gå och stäng dig inne i ditt hus.
Och se, du människobarn, bojor skola läggas på dig, och du skall bliva bunden med sådana, så att du icke kan gå ut bland de andra.
Och jag skall låta din tunga låda vid din gom, så att du bliver stum och icke kan bestraffa dem, då de nu äro ett gensträvigt släkte.
Men när jag talar med dig, skall jag upplåta din mun, så att du kan säga till dem: 'Så säger Herren, HERREN.'
Den som då vill höra, han höre, och den som icke vill, han höre icke, då de nu äro ett gensträvigt släkte.»
Och du, människobarn, tag dig en tegeltavla och lägg den framför dig och rista på den in en stad, nämligen Jerusalem.
Och res upp bålverk mot den och bygg en belägringsmur mot den och kasta upp en vall mot den och slå upp läger mot den och sätt upp murbräckor mot den runt omkring.
Och tag dig en järnplåt och sätt upp den såsom en järnvägg mellan dig och staden; och vänd så ditt ansikte emot den och håll den belägrad och ansätt den.
Detta skall vara ett tecken för Israels hus.
Och lägg du dig på din vänstra sida och lägg Israels hus' missgärning ovanpå; lika många dagar som du ligger så, skall du bära på deras missgärning.
Jag skall låta deras missgärningsår för dig motsvaras av ett lika antal dagar, nämligen av tre hundra nittio dagar; så länge skall du bara på Israels hus' missgärning.
Och sedan, när du har fullgjort detta, skall du lägga dig på din högra sida och bära på Juda hus' missgärning; i fyrtio dagar, var dag svarande mot ett år, skall denna min föreskrift gälla för dig.
Och du skall vända ditt ansikte och din blottade arm mot det belägrade Jerusalem och profetera mot det.
Och se, jag skall lägga bojor på dig, så att du icke kan vända dig från den ena sidan på den andra, förrän dina belägringsdagar äro slut.
Och tag dig vete, korn, bönor, linsärter, hirs och spält och lägg detta i ett och samma kärl och baka dig bröd därav; lika många dagar som du ligger på ena sidan, alltså tre hundra nittio dagar, skall detta vara vad du har att äta.
Den mat som du får att äta skall du äta efter vikt, tjugu siklar om dagen; detta skall du hava att äta från en viss timme ena dagen till samma timme nästa dag
Du skall ock dricka vatten efter mått, nämligen en sjättedels hin; så mycket skall du hava att dricka från en viss timme ena dagen till samma timme nästa dag.
Tillredd såsom kornkakor skall maten ätas av dig, och du skall tillreda den inför deras ögon på bränsle av människoträck.
Och HERREN tillade: »Likaså skola Israels barn äta sitt bröd orent bland hedningarna, till vilka jag skall fördriva dem.»
Men jag svarade: »Ack, Herre, HERRE!
Se, jag har ännu aldrig blivit orenad.
Jag har aldrig, från min ungdom och intill nu, ätit något självdött eller ihjälrivet djur; och sådant kött som räknas för vederstyggligt har aldrig kommit i min mun.»
Då sade han till mig: »Välan, jag vill låta dig taga kospillning i stället för människoträck; vid sådan må du baka ditt bröd.»
Och han sade åter till mig: »Du människobarn, se, jag vill fördärva livsuppehället för Jerusalem, så att de skola äta bröd efter vikt, och det med oro, och dricka vatten efter mått, och det med förfäran;
ja, så att de lida brist på bröd och vatten och gripas av förfäran, den ene med den andre, och försmäkta genom sin missgärning.
Och du, människobarn, tag dig ett skarpt svärd och bruka det såsom rakkniv, och för det över ditt huvud och din haka; tag dig så en vågskål och dela det avrakade håret.
En tredjedel skall du bränna upp i eld mitt i staden, när belägringsdagarna hava gått till ända; en tredjedel skall du taga ut och slå den med svärdet där runt omkring; och en tredjedel skall du strö ut för vinden, och mitt svärd skall jag draga ut efter dem.
Men några få strån skall du taga undan därifrån, och dem skall du knyta in i flikarna av din mantel.
Och av dessa strån skall du återigen taga några och kasta dem i elden och bränna upp dem i eld.
Härifrån skall en eld gå ut över hela Israels hus.
Så säger Herren, HERREN: Detta år Jerusalem, som jag har satt mitt ibland hednafolken, med länder runt däromkring.
Men det var gensträvigt mot mina rätter på ett ännu ogudaktigare sätt än hednafolken, och var ännu mer gensträvigt mot mina stadgar än länderna runt däromkring; ty de förkastade mina rätter och vandrade icke efter mina stadgar.
Därför säger Herren, HERREN så: Eftersom I haven rasat värre än hednafolken runt omkring eder, och icke haven vandrat efter mina stadgar och icke gjort efter mina rätter, ja, icke ens gjort efter de hednafolks rätter, som bo runt omkring eder,
därför säger Herren, HERREN så: Se, fördenskull skall jag också komma över dig och skipa rätt mitt ibland dig inför hednafolkens ögon;
jag skall göra med dig vad jag aldrig förr har gjort, och sådant som jag aldrig mer vill göra, för alla dina styggelsers skull.
Därför skola i dig föräldrar äta sina barn, och barn sina föräldrar; och jag skall skipa rätt i dig och strö ut för alla vindar allt som bliver kvar av dig.
Ja, så sant jag lever, säger Herren, HERREN: sannerligen, därför att du har orenat min helgedom med alla dina skändligheter och alla dina styggelser, skall jag också utan skonsamhet vända bort mitt öga och icke hava någon misskund.
En tredjedel av dig skall dö av pest och förgås av hunger i dig, en tredjedel skall falla för svärd runt omkring dig; och en tredjedel skall jag strö ut för alla vindar, och mitt svärd skall jag draga ut efter dem.
Ja, min vrede skall få uttömma sig, och jag skall släcka min förtörnelse på dem och hämnas på dem; och när jag så uttömmer min förtörnelse på dem, skola de förnimma att jag, HERREN, har talat i min nitälskan.
Och jag skall låta dig bliva en ödemark och en smälek bland folken runt omkring dig, inför var mans ögon, som går där fram.
Ja, det skall bliva till smälek och hån, till varnagel och skräck för folken runt omkring dig, när jag så skipar rätt i dig med vrede och förtörnelse och förtörnelses tuktan.
Jag, HERREN, har talat.
När jag sänder bland dem hungerns onda pilar, som bliva till fördärv, ja, när jag sänder dessa till att fördärva eder och så låter eder hunger bliva allt värre, då skall jag förstöra för eder edert livsuppehälle.
Jag skall sända över eder hungersnöd och vilddjur, som skola döda edra barn; och pest och blodsutgjutelse skall gå över dig, och svärd skall jag låta komma över dig.
Jag, HERREN, har talat.
Och HERRENS ord kom till mig; han sade:
Du människobarn, vänd ditt ansikte mot Israels berg och profetera mot dem
och säg: I Israels berg, hören Herrens, HERRENS ord: Så säger Herren, HERREN till bergen och höjderna, till bäckarna och dalarna: Se, jag skall låta svärd komma över eder och förstöra edra offerhöjder.
Och edra altaren skola varda förödda och edra solstoder sönderkrossade, och dem av eder, som bliva slagna, skall jag låta bliva kastade inför edra eländiga avgudar.
Och jag skall låta Israels barns döda kroppar ligga där inför deras eländiga avgudar, och jag skall förströ edra ben runt omkring edra altaren.
Var I än ären bosatta skola städerna bliva öde och offerhöjderna ödelagda, så att edra altaren stå öde och förödda, och edra eländiga avgudar bliva sönderslagna och få en ände, och edra solstoder bliva nedhuggna, och edra verk utplånade.
Dödsslagna män skola då falla bland eder; och I skolen förnimma att jag är HERREN.
Och om jag låter några leva kvar, så att somliga av eder, när I bliven förströdda i länderna, räddas undan svärdet ute bland folken,
så skola dessa edra räddade ute bland folken, där de äro i fångenskap, tänka på mig, när jag har krossat deras trolösa hjärtan, som veko av ifrån mig, och deras ögon, som i trolös avfällighet skådade efter deras eländiga avgudar; och de skola känna leda vid sig själva för det onda som de hava gjort med alla sina styggelser.
Och de skola förnimma att jag är HERREN.
Det är icke ett tomt ord att jag skall låta denna olycka komma över dem.
Så säger Herren, HERREN: Slå dina händer tillsammans, och stampa med dina fötter, och ropa ack och ve över alla de onda styggelserna i Israels hus, ty genom svärd, hunger och pest måste de falla.
Den som är långt borta skall dö av pest, och den som är nära skall falla för svärd, och den som bliver kvar och varder bevarad skall dö av hunger; så skall jag uttömma min vrede på dem.
Och I skolen förnimma att jag är HERREN, när deras slagna män ligga där mitt ibland sina eländiga avgudar, runt omkring sina altaren, på alla höga kullar, på alla bergstoppar, under alla gröna träd och under alla lummiga terebinter, varhelst de hava låtit en välbehaglig lukt uppstiga till alla sina oländiga avgudar.
Och jag skall uträcka min hand mot dem och göra landet mer öde och tomt än öknen vid Dibla, var de än äro bosatta; och de skola förnimma att jag är HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn, så säger Herren, HERREN till Israels land: Änden!
Ja, änden kommer över landets fyra hörn.
Nu kommer änden över dig, ty jag skall sända min vrede mot dig och döma dig efter dina gärningar och låta alla dina styggelser komma över dig.
Jag skall icke visa dig någon skonsamhet och icke hava någon misskund; nej, jag skall låta dina gärningar komma över dig, och dina styggelser skola vila på dig.
Och I skolen förnimma att jag är HERREN.
Så säger Herren, HERREN: Se, en olycka kommer, en olycka ensam i sitt slag!
En ände kommer, ja, änden kommer, den vaknar upp och kommer över dig.
Ja se, det kommer!
Nu kommer ordningen till dig, du folk som bor här i landet; din stund kommer, förvirringens dag är nära, då intet skördeskri mer skall höras på bergen.
Nu skall jag snart utgjuta min förtörnelse över dig och uttömma min vrede på dig, och döma dig efter dina gärningar och låta alla dina styggelser komma över dig.
Jag skall icke visa någon skonsamhet och icke hava någon misskund, jag skall giva dig efter dina gärningar, och dina styggelser skola vila på dig.
Och I skolen förnimma att jag, HERREN, är den som slår.
Se, dagen är inne; se, det kommer!
Ordningen går sin gång, riset blomstrar upp, övermodet grönskar;
våldet reser sig till ett ris för ogudaktigheten.
Då bliver intet kvar av dem, intet av hela deras hop, intet av deras gods, och till intet bliver deras härlighet.
Stunden kommer, dagen nalkas; köparen må icke glädja sig, och säljaren må icke sörja, ty vredesglöd kommer över hela hopen därinne.
Säljaren skall icke få tillbaka vad han har sålt, om han ens får förbliva vid liv.
Ty profetian om hela hopen därinne skall icke ryggas och ingen som lever i missgärning skall kunna hålla stånd.
Man stöter i basun och rustar allt i ordning, men ingen drager ut till strid; ty min vredesglöd går fram över hela hopen därinne.
Ute härjar svärdet och därinne pest och hungersnöd, den som är ute på marken dör genom svärdet, och den som är i staden, honom förtär hungersnöd och pest.
Och om några av dem bliva räddade, så skola de söka sin tillflykt i bergen och vara lika klyftornas duvor, som allasammans klaga.
Så skall det gå var och en genom hans missgärning.
Alla händer skola sjunka ned, och alla knän skola bliva såsom vatten.
Människorna skola kläda sig i sorgdräkt, och förfäran skall övertäcka dem, alla ansikten skola höljas av skam, och alla huvuden skola bliva skalliga.
Man skall kasta sitt silver ut på gatorna och akta sitt guld såsom orenlighet.
Deras silver och guld skall icke kunna rädda dem på HERRENS vredes dag, de skola icke kunna mätta sig därmed eller därmed fylla sin buk; ty det har varit för dem en stötesten till missgärning.
Dess sköna glans brukade man till högfärd, ja, de gjorde därav sina styggeliga bilder, sina skändliga avgudar.
Därför skall jag göra det till orenlighet för dem.
Jag skall giva det såsom byte i främlingars hand och såsom rov åt de ogudaktigaste på jorden, för att de må ohelga det.
Och jag skall vända bort mitt ansikte ifrån dem, så att man får ohelga min klenod; våldsmän skola få draga därin och ohelga den.
Gör kedjorna redo; ty landet är fullt av blodsdomar, och staden är full av orätt.
Och jag skall låta de värsta hednafolk komma och taga deras hus i besittning.
Så skall jag göra slut på de fräckas övermod, och deras helgedomar skola varda oskärade.
Förskräckelse skall komma, och när de söka räddning, skall ingen vara att finna.
Den ena olyckan skall komma efter den andra, det ena sorgebudet skall följa det andra.
Man skall få tigga profeterna om syner, prästerna skola komma till korta med sin undervisning och de äldste med sina råd.
Konungen skall sörja, hövdingarna skola kläda sig i förskräckelse, och folket i landet skall stå där med darrande händer.
Jag skall göra med den efter deras gärningar och skipa rätt åt dem såsom rätt är åt dem; och de skola förnimma att jag är HERREN.
Och i sjätte året, i sjätte månaden, på femte dagen i månaden, när jag satt i mitt hus och de äldste i Juda sutto hos mig, kom Herrens, HERRENS hand där över mig.
Och jag fick se något som till utseendet liknade eld; allt, ända ifrån det som såg ut att vara hans länder och sedan allt nedåt, var eld.
Men från hans länder och sedan allt uppåt syntes något som liknade strålande ljus, och som var såsom glänsande malm.
Och han räckte ut något som var bildat såsom en hand och fattade mig vid en lock av mitt huvudhår; och en andekraft lyfte mig upp mellan himmel och jord och förde mig, i en syn från Gud, till Jerusalem, dit där man går in till den inre förgården genom den port som vetter åt norr, där varest avgudabelätet, det som hade uppväckt Guds nitälskan, hade sin plats.
Och se, där syntes Israels Guds härlighet, alldeles sådan som jag hade sett den på slätten.
Och han sade till mig: »Du människobarn, lyft upp dina ögon mot norr.»
När jag nu lyfte upp mina ögon mot norr, fick jag se avgudabelätet, det som hade uppväckt Guds nitälskan, stå där norr om altarporten, vid själva ingången.
Och han sade till mig: »Du människobarn, ser du vad de göra här?
Stora äro de styggelser som Israels hus här bedriver, så att jag måste draga långt bort ifrån min helgedom; men du skall få se ännu flera, större styggelser.»
Sedan förde han mig till förgårdens ingång, och jag fick där se ett hål i väggen.
Och han sade till mig: »Du människobarn, bryt igenom väggen.»
Då bröt jag igenom väggen och fick nu se en dörr.
Och han sade till mig: »Gå in och se vilka onda styggelser de här bedriva.»
När jag nu kom in, fick jag se allahanda bilder av vederstyggliga kräldjur och fyrfotadjur, så ock Israels hus' alla eländiga avgudar, inristade runt omkring på väggarna.
Och framför dem stodo sjuttio av: de äldste i Israels hus, och Jaasanja, Safans son, stod mitt ibland dem, och var och en av dem hade sitt rökelsekar i handen, och vällukt steg upp från rökelsemolnet.
Och han sade till mig: »Du människobarn, ser du vad de äldste i Israels hus bedriva i mörkret, var och en i sin avgudakammare?
Ty de säga: 'HERREN ser oss icke, HERREN har övergivit landet.'»
Därefter sade han till mig: »Du skall få se ännu flera, större styggelser som dessa bedriva.»
Och han förde mig fram mot ingången till norra porten på HERRENS hus, och se, där sutto kvinnor som begräto Tammus.
Och han sade till mig: »Du människobarn, ser du detta?
Men du skall få se ännu flera styggelser, större än dessa.»
Och han förde mig till den inre förgården till HERRENS hus, och se, vid ingången till HERRENS tempel, mellan förhuset och altaret, stodo vid pass tjugufem män, som vände ryggarna åt HERRENS tempel och ansiktena åt öster, och som tillbådo solen i öster.
Och han sade till mig: »Du människobarn, ser du detta?
Är det icke nog för Juda hus att bedriva de styggelser som de här hava bedrivit, eftersom de nu ock hava uppfyllt landet med orätt och åter hava förtörnat mig?
Se nu huru de sätta vinträdskvisten för näsan!
Därför skall också jag utföra mitt: verk i vrede; jag skall icke visa någon skonsamhet och icke hava någon misskund.
Och om de än ropa med hög röst inför mig, skall jag dock icke höra dem.»
Och jag hörde honom ropa med hög röst och säga: »Kommen hit med hemsökelser över staden, och var och en have sitt mordvapen i handen.»
Och se, då kommo sex män från övre porten, den som vetter åt norr och var och en hade sin stridshammare i handen; och bland dem fanns en man som var klädd i linnekläder och hade ett skrivtyg vid sin länd.
Och de kommo och ställde sig vid sidan av kopparaltaret.
Och Israels Guds härlighet hade lyft sig från keruben, som den vilade på, och hade flyttat sig till tempelhusets tröskel, och ropade nu till mannen som var klädd i linnekläderna och hade skrivtyget vid sin länd;
HERREN sade till honom: »Gå igenom Jerusalems stad, och teckna med ett tecken på pannan de män som sucka och jämra sig över alla styggelser som bedrivas därinne.»
Och till de andra hörde jag honom säga: »Dragen fram i staden efter honom och slån ned folket; visen ingen skonsamhet och haven ingen misskund.
Både åldringar och ynglingar och jungfrur, både barn och kvinnor skolen I dräpa och förgöra, men I mån icke komma vid någon som har tecknet på sig, och I skolen begynna vid min helgedom.»
Och de begynte med de äldste, med de män som stodo framför tempelhuset.
Han sade nämligen till dem: »Orenen tempelhuset, och fyllen upp förgårdarna med slagna; dragen sedan ut.»
Och de drogo ut och slogo ned folket i staden.
Då nu jag blev lämnad kvar, när de så slogo folket, föll jag ned på mitt ansikte och ropade och sade: »Ack, Herre, HERRE, vill du då förgöra hela kvarlevan av Israel, eftersom du så utgjuter din vrede över Jerusalem?»
Han sade till mig: »Israels och Juda hus' missgärning är alltför stor; landet är uppfyllt med orätt, och staden är full av lagvrängning.
Ty de säga: 'HERREN har övergivit landet, HERREN ser det icke.'
Därför skall icke heller jag visa någon skonsamhet eller hava någon misskund, utan skall låta deras gärningar komma över deras huvuden.»
Och mannen som var klädd i linnekläderna och hade skrivtyget vid sin länd kom nu tillbaka och gav besked och sade: »Jag har gjort såsom du bjöd mig.»
Och jag fick se att på fästet, som vilade på kerubernas huvuden, fanns något som tycktes vara av safirsten, något som till utseendet liknade en tron; detta syntes ovanpå dem.
Och han sade till mannen som var klädd i linnekläderna, han sade: »Gå in mellan rundlarna, in under keruben, och tag dina händer fulla med eldsglöd från platsen mellan keruberna, och strö ut dem över staden.»
Och jag såg honom gå.
Och keruberna stodo till höger om huset, när mannen gick ditin, och molnet uppfyllde den inre förgården.
Men HERRENS härlighet höjde sig upp från keruben och flyttade sig till husets tröskel; och huset uppfylldes då av molnet, och förgården blev full av glansen från HERRENS härlighet.
Och dånet av kerubernas vingar hördes ända till den yttre förgården, likt Gud den Allsmäktiges röst, då han talar.
Och när han nu bjöd mannen som var klädd i linnekläderna och sade: »Tag eld från platsen mellan rundlarna, inne mellan keruberna», då gick denne ditin och ställde sig bredvid ett av hjulen.
Då räckte keruben där ut sin hand, mellan de andra keruberna, till elden som brann mellan keruberna, och tog därav och lade i händerna på honom som var klädd i linnekläderna; och denne tog det och gick så ut.
Och under vingarna på keruberna så syntes något som var bildat såsom en människohand.
Och jag fick se fyra hjul stå invid keruberna ett hjul invid var kerub och det såg ut som om hjulen voro av något som liknade krysolitsten.
De sågo alla fyra likadana ut, och ett hjul tycktes vara insatt i ett annat.
När de skulle gå, kunde de gå åt alla fyra sidorna, de behövde icke vända sig, när de gingo.
Ty åt det håll dit den främste begav sig gingo de andra efter, utan att de behövde vända sig, när de gingo.
Och hela deras kropp, deras rygg, deras händer och deras vingar, så ock hjulen, voro fulla med ögon runt omkring; de fyra hade nämligen var sitt hjul.
Och jag hörde att hjulen kallades »rundlar».
Och var och en hade fyra ansikten; det första ansiktet var en kerubs, det andra en människas, det tredje ett lejons, det fjärde en örns.
Och keruberna höjde sig upp; de var samma väsenden som jag hade sett vid strömmen Kebar.
Och när keruberna gingo, gingo ock hjulen invid dem; och när keruberna lyfte sina vingar för att höja sig över jorden, skilde sig hjulen icke ifrån dem.
När de stodo stilla, stodo ock dessa stilla, och när de höjde sig, höjde sig ock dessa med dem, ty väsendenas ande var i dem.
Och HERRENS härlighet flyttade I sig bort ifrån husets tröskel och stannade över keruberna.
Då såg jag huru keruberna lyfte sina vingar och höjde sig från jorden, när de begåvo sig bort, och hjulen jämte dem; och de stannade vid ingången till östra porten på HERRENS hus, och Israels Guds härlighet vilade ovanpå dem.
Det var samma väsenden som jag: hade sett under Israels Gud vid strömmen Kebar, och jag märkte att det var keruber.
Var och en hade fyra ansikten och fyra vingar, och under deras vingar var något som liknade människohänder.
Och deras ansikten voro likadana som de ansikten jag hade sett vid strömmen Kebar, så sågo de ut, och sådana voro de.
Och de gingo alla rakt fram.
Och en andekraft lyfte upp mig och förde mig till östra porten på HERRENS hus, den som vetter åt öster.
Där fick jag se tjugufem män stå vid ingången till porten; och jag såg bland dem Jaasanja, Assurs son, och Pelatja, Benajas son, som voro furstar i folket.
Och han sade till mig: »Du människobarn, det är dessa män som tänka ut vad fördärvligt är och råda till vad ont är, här i staden;
det är de som säga: 'Hus byggas icke upp så snart.
Här är grytan, och vi äro köttet.
Profetera därför mot dem, ja, profetera, du människobarn.»
Då föll HERRENS Ande över mig, han sade till mig: »Säg: Så säger HERREN: Sådant sägen I, I av Israels hus, och edra hjärtans tankar känner jag väl.
Många ligga genom eder slagna här i staden; I haven uppfyllt dess gator med slagna.
Därför säger Herren, HERREN så: De slagna vilkas fall I haven vållat i staden, de äro köttet, och den är grytan; men eder själva skall man föra bort ur den.
I frukten för svärd, och svärd skall jag ock låta komma över eder, säger Herren, HERREN.
Jag skall föra eder bort härifrån och giva eder i främlingars hand; och jag skall hålla dom över eder.
För svärd skolen I falla; vid Israels gräns skall jag döma eder.
Och I skolen förnimma att jag är HERREN.
Staden skall icke vara en gryta för eder, och I skolen icke vara köttet i den; nej, vid Israels gräns skall jag döma eder.
Då skolen I förnimma att jag är HERREN, I som icke haven vandrat efter mina stadgar och icke haven gjort efter mina rätter, utan haven gjort efter de hednafolks rätter, som bo runt omkring eder.»
Medan jag så profeterade, hade Pelatja, Benajas son, uppgivit andan.
Då föll jag ned på mitt ansikte och ropade med hög röst och sade: »Ack, Herre, HERRE, vill du då alldeles göra ände på kvarlevan av Israel?»
Och HERRENS ord kom till mig; han sade:
»Du människobarn, dina bröder, ja, dina bröder dina nära fränder och hela Israels hus, alla de till vilka Jerusalems invånare säga: 'Hållen eder borta från HERREN; det är åt oss som landet har blivit givet till besittning' --
om dem skall du alltså säga: Så säger Herren, HERREN: Ja, väl har jag fört dem långt bort ibland folken och förstrött dem i länderna, och med nöd har jag varit för dem en helgedom i de länder dit de hava kommit;
men därför skall du nu säga: Så säger Herren, HERREN: Jag skall församla eder ifrån folkslagen och hämta eder tillhopa från de länder dit I haven blivit förströdda, och skall giva eder Israels land.
Och när de hava kommit dit, skola de skaffa bort därifrån alla de skändliga och styggeliga avgudar som nu finnas där.
Och jag skall giva dem alla ett och samma hjärta, och en ny ande skall jag låta komma i deras bröst; jag skall taga bort stenhjärtat ur deras kropp och giva dem ett hjärta av kött,
så att de vandra efter mina stadgar och hålla mina rätter och göra efter dem, och de skola vara mitt folk, och jag skall vara deras Gud.
Men de vilkas hjärtan efterfölja de skändliga och styggeliga avgudarnas hjärtan, deras gärningar skall jag låta komma över deras huvuden, säger Herren, HERREN.»
Och keruberna, följda av hjulen, lyfte sina vingar, och Israels Guds härlighet vilade ovanpå dem.
Och HERRENS härlighet höjde sig och lämnade staden och stannade på berget öster om staden.
Men mig hade en andekraft lyft upp och fört bort till de fångna i Kaldeen, så hade skett i synen, genom Guds Ande.
Sedan försvann för mig den syn jag hade fått se.
Och jag talade till de fångna alla de ord som HERREN hade uppenbarat för mig.
Och HERRENS ord kom till mig; han sade;
»Du människobarn, du bor mitt i det gensträviga släktet, bland människor som hava ögon att se med, men dock icke se, och öron att höra med, men dock icke höra, eftersom de äro ett så gensträvigt släkte.
Så red nu till åt dig, du människobarn, vad man behöver, när man skall gå i landsflykt.
Och vandra i deras åsyn åstad på ljusa dagen, ja, vandra i deras åsyn åstad från det ställe där du nu bor bort till en annan ort -- om de till äventyrs ville akta därpå, då de nu äro ett så gensträvigt släkte.
För ut ditt bohag, på ljusa dagen och i deras åsyn, såsom skulle du gå i landsflykt, och vandra så i deras åsyn själv åstad på aftonen, såsom landsflyktiga pläga.
Gör dig i deras åsyn en öppning i väggen, och för bohaget ut genom den.
Lyft det sedan i deras åsyn upp på axeln och för bort det, när det har blivit alldeles mörkt; och betäck ditt ansikte, så att du icke ser landet.
Ty jag gör dig till ett tecken för Israels hus.»
Och jag gjorde såsom han bjöd mig; på ljusa dagen förde jag ut mitt bohag, såsom skulle jag gå i landsflykt.
Sedan, om aftonen, gjorde jag mig med handen en öppning i väggen, och när det hade blivit alldeles mörkt, förde jag det ut genom den och bar det så på axeln, i deras åsyn.
Och HERRENS ord kom till mig den följande morgonen; han sade:
Du människobarn, säkert har Israels hus, det gensträviga släktet, frågat dig: »Vad är det du gör?»
Så svara dem nu: Så säger Herren, HERREN: Denna utsaga gäller fursten i Jerusalem och alla dem av Israels hus, som äro därinne.
Säg: Jag är ett tecken för eder; såsom jag har gjort, så skall det gå dem: de skola vandra bort i landsflykt och fångenskap.
Och fursten som de hava ibland sig skall lyfta upp sin börda på axeln, när det har blivit alldeles mörkt, och skall så draga ut.
Man skall göra en öppning i väggen, så att han genom den kan bära ut sin börda; och han skall betäcka sitt ansikte, så att han icke ser landet med sitt öga.
Och jag skall breda ut mitt nät över honom, och han skall bliva fångad i min snara; och jag skall föra honom till Babel i kaldéernas land, som han dock icke skall se; och där skall han dö.
Och alla som äro omkring honom, till hans hjälp, och alla hans härskaror skall jag förströ åt alla väderstreck, och mitt svärd skall jag draga ut efter dem.
Och de skola förnimma att jag är HERREN, när jag förskingrar dem bland folken och förströr dem i länderna.
Men några få av dem skall jag låta bliva kvar efter svärd, hungersnöd och pest, för att de bland de folk till vilka de komma skola kunna förtälja om alla sina styggelser; och de skola förnimma att jag är HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn, ät nu ditt bröd med bävan, och drick ditt vatten darrande och med oro.
Och säg till folket i landet: Så säger Herren, HERREN om Jerusalems invånare i Israels land: De skola äta sitt bröd med oro och dricka sitt vatten med förfäran; så skall landet bliva ödelagt och plundrat på allt vad däri är, för den orätts skull som alla dess inbyggare hava övat.
Och de städer som nu äro bebodda skola komma att ligga öde, och landet skall bliva en ödemark; och I skolen förnimma att jag är HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn, vad är det för ett ordspråk I haven i Israels land, när I sägen: »Tiden går, och av alla profetsynerna bliver intet»?
Säg nu till dem: Så säger Herren, HERREN: Jag skall göra slut på det ordspråket, så att man icke mer skall bruka det i Israel.
Tala i stället så till dem: »Tiden kommer snart, med alla profetsynernas fullbordan.»
Ty inga falska profetsyner och inga lögnaktiga spådomar skola mer finnas i Israels hus;
nej, jag, HERREN, skall tala det ord som jag vill tala, och det skall fullbordas, utan att länge fördröjas.
Ja, du gensträviga släkte, i edra dagar skall jag tala ett ord och skall ock fullborda det, säger Herren, HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn, se, Israels hus säger: »Den syn som han skådar gäller dagar som icke komma så snart; han profeterar om tider som ännu äro långt borta.»
Säg därför till dem: Så säger Herren, HERREN: Intet av vad jag har talat skall längre fördröjas; vad jag talar, det skall ske, säger Herren, HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn, profetera mot Israels profeterande profeter; säg till dem som profetera efter sina egna hjärtans ingivelser: Hören HERRENS ord.
Så säger Herren, HERREN: Ve eder, I dåraktiga profeter, som följen eder egen ande och syner som I icke haven sett! --
Lika rävar på öde platser äro dina profeter, Israel.
I haven icke trätt fram i gapet eller fört upp någon mur omkring Israels hus, så att det har kunnat bestå i striden på HERRENS dag.
Nej, deras syner voro falskhet och deras spådomar lögn, fastän de sade »Så har HERREN sagt.»
HERREN hade ju icke sänt dem, men de hoppades att deras tal ändå skulle gå i fullbordan.
Ja, förvisso var det falska syner som I skådaden och lögnaktiga spådomar som I uttaladen, fastän I saden: »Så har HERREN sagt.»
Jag hade ju icke talat något sådant.
Därför säger Herren, HERREN så: Eftersom edert tal är falskhet och edra syner äro lögn, se, därför skall jag komma över eder, säger Herren, HERREN.
Och min hand skall drabba profeterna som skåda falska syner och spå lögnaktiga spådomar.
De skola icke få en plats i mitt folks församling och skola icke bliva upptagna i förteckningen på Israels hus, ej heller skola de få komma till Israels land; och I skolen förnimma att jag är Herren, HERREN.
Eftersom, ja, eftersom de förde mitt folk vilse, i det att de sade: »Allt står väl till», och dock stod icke allt väl till, och eftersom de, när folket bygger upp en mur, vitmena den,
därför må du säga till dessa vitmenare att den måste falla.
Ett slagregn skall komma -- ja, I skolen fara ned, I hagelstenar, och du skall bryta ned den, du stormvind!
Och när så väggen faller, då skall man förvisso säga till eder: »Var är nu vitmeningen som I ströken på?»
Därför säger Herren, HERREN så; Jag skall i min förtörnelse låta en stormvind bryta lös, ett slagregn skall komma genom min vrede, och hagelstenar genom min förtörnelse, så att det bliver en ände därpå.
Och jag skall förstöra väggen som I beströken med vitmening, jag skall slå den till jorden, så att dess grundval bliver blottad.
Och när den faller, skolen I förgås därinne; och I skolen förnimma att jag är HERREN.
Och jag skall uttömma min förtörnelse på väggen och på dem som hava bestrukit den med vitmening; och så skall jag säga till eder: Det är ute med väggen, det är ute med dess vitmenare,
med Israels profeter, som profeterade om Jerusalem och skådade syner, det till behag, om att allt stod väl till, och dock stod icke allt väl till, säger Herren, HERREN.
Och du, människobarn, vänd ditt ansikte mot dina landsmaninnor som profetera efter sina egna hjärtans ingivelser; profetera mot dem
och säg: Så säger Herren, HERREN: Ve eder som syn bindlar till alla handleder och gören slöjor till alla huvuden, både ungas och gamlas, för att så fånga själar!
Skullen I få fånga själar bland mitt folk och döma somliga själar till liv, eder till vinning,
I som för några nävar korn och några bitar bröd ohelgen mig hos mitt folk, därmed att I dömen till döden själar som icke skola dö, och dömen till liv själar som icke skola leva, i det att I ljugen för mitt folk, som gärna hör lögn?
Nej, och därför säger Herren, HERREN så: Se, jag skall väl nå edra bindlar, i vilka I fången själarna såsom fåglar, och skall slita dem från edra armar; och jag skall giva själarna fria, de själar som I haven fångat såsom fåglar.
Och jag skall slita sönder edra slöjor och rädda mitt folk ur eder hand, och de skola icke mer vara ett byte i eder hand; och I skolen förnimma att jag är HERREN.
Eftersom I genom lögnaktigt tal haven gjort den rättfärdige försagd i hjärtat, honom som jag ingalunda ville plåga, men däremot haven styrkt den ogudaktiges mod, så att han icke vänder om från sin onda väg och räddar sitt liv,
därför skolen I icke få fortsätta att skåda falska syner och att öva spådom; utan jag skall rädda mitt folk ur eder hand, och I skolen förnimma att jag är HERREN.
Och några av de äldste i Israel kommo till mig och satte sig ned hos mig.
Då kom HERRENS ord till mig; han sade:
Du människobarn, dessa män hava låtit sina eländiga avgudar få insteg i sina hjärtan och hava ställt upp framför sig vad som är dem en stötesten till missgärning.
Skulle jag väl låta fråga mig av sådana?
Nej; tala därför med dem och säg till dem: Så säger Herren, HERREN: Var och en av Israels hus, som låter sina eländiga avgudar få insteg i sitt hjärta och ställer upp framför sig vad som är honom en stötesten till missgärning, och så kommer till profeten, honom skall jag, HERREN, giva svar såsom han har förtjänat genom sina många eländiga avgudar.
Så skall jag gripa Israels barn i hjärtat, därför att de allasammans hava vikit bort ifrån mig genom sina eländiga avgudar.
Säg därför till Israels hus: Så säger Herren, HERREN: Vänden om, ja, vänden eder bort ifrån edra eländiga avgudar, vänden edra ansikten bort ifrån alla edra styggelser.
Ty om någon av Israels hus, eller av främlingarna som bo i Israel, viker bort ifrån mig, och låter sina eländiga avgudar få insteg i sitt hjärta och ställer upp framför sig vad som är honom en stötesten till missgärning, och så kommer till profeten, för att denne skall fråga mig för honom, så vill jag, HERREN, själv giva honom svar:
jag skall vända mitt ansikte mot den mannen och göra honom till ett tecken och till ett ordspråk, och utrota honom ur mitt folk; och I skolen förnimma att jag är HERREN.
Men om profeten låter förföra sig och talar något ord, så har jag, HERREN, låtit den profeten bliva förförd; och jag skall uträcka min hand mot honom och förgöra honom ur mitt folk Israel.
Och de skola båda bära på sin missgärning: profetens missgärning skall räknas lika med den frågandes missgärning --
på det att Israels barn icke mer må gå bort ifrån mig och fara vilse, ej heller mer orena sig med alla sina överträdelser, utan vara mitt folk, såsom jag skall vara deras Gud, säger Herren, HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn, om ett land syndade mot mig och beginge otrohet, så att jag måste uträcka min hand mot det och fördärva dess livsuppehälle och sända hungersnöd över det och utrota därur både människor och djur,
och om då därinne funnes dessa tre män: Noa, Daniel och Job, så skulle de genom sin rättfärdighet rädda allenast sina egna liv, säger Herren, HERREN.
Om jag läte vilddjur draga fram genom landet och göra det folktomt, så att det bleve så öde att ingen vågade draga där fram för djuren skull,
då skulle, så sant jag lever, säger Herren, HERREN, dessa tre män, om de vore därinne, icke kunna rädda vare sig söner eller döttrar; allenast de själva skulle räddas, men landet måste bliva öde.
Eller om jag läte svärd komma över det landet, i det att jag sade: »Svärdet fare fram genom landet!», och jag så utrotade därur både människor och djur,
och om då dessa tre män vore därinne, så skulle de, så sant jag lever, säger Herren, HERREN, icke kunna rädda söner eller döttrar; allenast de själva skulle räddas.
Eller om jag sände pest i det landet och utgöte min vrede däröver i blod, för att utrota därur både människor och djur,
och om då Noa, Daniel och Job vore därinne, så skulle de, så sant jag lever, säger Herren, HERREN, icke kunna rädda vare sig son eller dotter; de skulle genom sin rättfärdighet rädda allenast sina egna liv.
Och så säger Herren, HERREN: Men huru mycket värre bliver det icke, när jag på en gång sänder mina fyra svåra straffdomar: svärd, hungersnöd, vilddjur och pest, över Jerusalem, för att utrota därur både människor och djur!
Likväl skola några räddade bliva kvar där, några söner och döttrar, som skola föras bort.
Och se, dessa skola draga bort till eder; och när I fån se deras vandel och deras gärningar, då skolen I trösta eder för den olycka som jag har låtit komma över Jerusalem, ja, för allt som jag har låtit komma över det.
De skola vara eder till tröst, när I sen deras vandel och deras gärningar; I skolen då förstå att jag icke utan sak har gjort allt vad jag har gjort mot det, säger Herren, HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn, varutinnan är vinstockens trä förmer än annat trä, vinstockens, vars rankor växa upp bland skogens andra träd?
Tager man väl virke därav till att förfärdiga något nyttigt?
Gör man ens därav en plugg för att på den hänga upp någonting?
Och om det nu därtill har varit livet till mat åt elden, så att dess båda ändar hava blivit förtärda av eld, och vad däremellan finnes är svett, duger det då till något nyttigt?
Icke ens medan det ännu var oskadat, kunde man förfärdiga något nyttigt därav; huru mycket mindre kan man förfärdiga något nyttigt därav, sedan det endels har blivit förtärt av elden och endels är svett!
Därför säger Herren, HERREN så: Såsom det händer med vinstockens trä bland annat trä från skogen, att Jag lämnar det till mat åt elden, så skall jag ock göra med Jerusalems invånare.
Jag skall vända mitt ansikte mot dem; ur elden hava de kommit undan, men eld skall dock förtära dem.
Och I skolen förnimma att jag är HERREN, när jag vänder mitt ansikte mot dem.
Och jag skall göra landet till en ödemark, därför att de hava varit otrogna, säger Herren, HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn, förehåll Jerusalem dess styggelser
och säg: Så säger Herren, HERREN till Jerusalem: Från Kanaans land stammar du, och där är du född; din fader var en amoré och din moder en hetitisk kvinna.
Och vid din födelse gick det så till.
När du föddes, skar ingen av din navelsträng, och du blev icke rentvagen med vatten, ej heller ingniden med salt och lindad.
Ingen såg på dig med så mycken ömkan, att han villa göra något sådant med dig eller visa dig någon misskund, utan man kastade ut dig på öppna fältet den dag du föddes; så ringa aktade man ditt liv.
Då gick jag förbi där du låg och fick se dig sprattla i ditt blod, och jag sade till dig: »Du skall få bliva vid liv, du som ligger där i ditt blod.»
Ja, jag sade till dig: »Du skall få bliva vid liv, du som ligger där i ditt blod;
ja, jag skall föröka dig till många tusen, såsom växterna äro på marken.»
Och du sköt upp och blev stor och mycket fager; dina bröst hade höjt sig, och ditt hår hade växt, men du var ännu naken och blottad.
Då gick jag åter förbi där du var och fick se att din tid var inne, din älskogstid; och jag bredde min mantel över dig och betäckte din blygd.
Och så gav jag dig min ed och ingick förbund med dig, säger Herren, HERREN, och du blev min.
Och jag tvådde dig med vatten och sköljde blodet av dig, och smorde dig med olja,
och klädde på dig brokigt vävda kläder och satte på dig skor av tahasskinn och en huvudbindel av fint linne och en slöja av silke.
Och jag prydde dig med smycken: jag satte armband på dina armar och en kedja om din hals,
jag satte en ring i din näsa och örhängen i dina öron och en härlig krona på ditt huvud.
Så blev du prydd med guld och silver, och dina kläder voro av fint linne, av siden och av tyg i brokig vävnad.
Fint mjöl, honung och olja fick du äta.
Du blev övermåttan skön, och så vart du omsider en drottning.
Och ryktet om dig gick ut bland folken för din skönhets skull, ty den var fullkomlig genom de härliga prydnader som jag hade satt på dig, säger Herren, HERREN.
Men du förlitade dig på din skönhet och bedrev otukt, sedan du nu hade fått sådant rykte; du slösade din otukt på var och en som gick där fram: det vore ju något för honom.
Och du tog dina kläder och gjorde dig med dem brokiga offerhöjder och bedrev på dessa otukt, sådana gärningar som eljest aldrig någonsin hava förekommit, ej heller mer skola göras.
Och du tog dina härliga smycken, det guld och silver som jag hade givit dig, och gjorde dig så mansbilder, med vilka du bedrev otukt.
Och du tog dina brokigt vävda kläder och höljde dem i dessa; och min olja och min rökelse satte du fram för dem.
Och det bröd som jag hade givit dig -- ty fint mjöl, olja och honung hade jag ju låtit dig få att äta -- detta satte du fram för dem till en välbehaglig lukt; ja, därhän kom det, säger Herren, HERREN.
Och du tog dina söner och döttrar, dem som du hade fött åt mig, och offrade dessa åt dem till spis.
Var det då icke nog att du bedrev otukt?
Skulle du också slakta mina söner och giva dem till pris såsom offer åt dessa?
Och vid alla dina styggelser och din otukt tänkte du icke på din ungdoms dagar, då du var naken och blottad och låg där sprattlande i ditt blod.
Och sedan du hade bedrivit all denna ondska -- ve, ve dig! säger Herren, HERREN --
byggde du dig kummel och gjorde dig höjdaltaren på alla öppna platser.
I alla gathörn byggde du dig höjd altaren och lät din skönhet skända och spärrade ut benen åt alla som gingo där fram; ja, du bedrev mycken otukt.
Du bedrev otukt med egyptierna, dina grannar med det stora köttet, ja, mycken otukt till att förtörna mig.
Men se, då uträckte jag min hand mot dig och minskade ditt underhåll och gav dig till pris åt dina fiender, filistéernas döttrar, som blygdes över ditt skändliga väsende.
Men sedan bedrev du otukt med assyrierna, ty du hade ännu icke blivit mätt; ja, du bedrev otukt med dem och blev ändå icke mätt.
Du gick med din otukt ända bort till krämarlandet, kaldéernas land; men icke ens så blev du mätt.
Huru älskogskrankt var icke ditt hjärta, säger Herren, HERREN, eftersom du gjorde allt detta, sådana gärningar som allenast den fräckaste sköka kan göra.
Med dina döttrar uppförde du åt dig kummel i alla gathörn och höjdaltaren på alla öppna platser.
Men däri var du olik andra skökor, att du försmådde skökolön,
du äktenskapsbryterska, som i stället för den man du hade tog andra män till dig.
Åt alla andra skökor måste man giva skänker, men här var det du som gav skänker åt alla dina älskare och mutade dem, för att de skulle komma till dig från alla håll och bedriva otukt med dig.
Så gjorde du vid din otukt tvärt emot vad andra kvinnor göra; efter dig lopp ingen för att bedriva otukt, men du gav skökolön, utan att själv få någon skökolön; du gjorde tvärt emot andra.
Hör därför HERRENS ord, du sköka.
Så säger Herren, HERREN: Eftersom du har varit så frikostig med din skam och blottat din blygd i otukt med din älskare, därför, och för alla dina vederstyggliga eländiga avgudars skull och för dina söners blods skull, dina söners, som du gav åt dessa,
se, därför skall jag församla alla dina älskare, dem som du har varit till behag, ja, alla dem som du har älskat mer eller mindre; dem skall jag församla mot dig från alla håll och blotta din blygd inför dem, så att de få se all din blygd.
Och jag skall döma dig efter den lag som gäller för äktenskapsbryterskor och blodsutgjuterskor, och skall låta dig bliva ett blodigt offer för min vrede och nitälskan.
Och jag skall giva dig i deras hand, och de skola slå ned dina kummel och bryta ned dina höjdaltaren, och slita av dig kläderna och taga ifrån dig dina härliga smycken och låta dig ligga naken och blottad.
Och de skola sammankalla en församling mot dig, och man skall stena dig och hugga sönder dig med svärd;
och dina hus skall man bränna upp i eld.
Så skall man hålla dom över dig inför många kvinnors ögon.
Och så skall jag göra slut på din otukt, och du skall icke mer kunna giva någon skökolön.
Och jag skall släcka min vrede på dig, så att min nitälskan kan vika ifrån dig, och så att jag får ro och slipper att mer förtörnas.
Eftersom du icke tänkte på din ungdoms dagar, utan var avog mot mig i allt detta, se, därför skall också jag låta dina gärningar komma över ditt huvud, säger Herren, HERREN, på det att du icke mer må lägga sådan skändlighet till alla dina andra styggelser.
Se, alla som bruka ordspråk skola på dig tillämpa det ordspråket: »Sådan moder, sådan dotter.»
Ja, du är din moders dotter, hennes som övergav sin man och sina barn; du är dina systrars syster deras som övergåvo sina män och sina barn; eder moder var en hetitisk kvinna och eder fader en amoré.
Din större syster var Samaria med sina döttrar, hon som bodde norrut från dig; och din mindre syster, som bodde söderut från dig, var Sodom med sina döttrar.
Men du nöjde dig icke med att vandra på deras vägar och att göra efter deras styggelser; inom kort bedrev du värre ting än de, på alla dina vägar.
Så sant jag lever, säger Herren, HERREN: din syster Sodom och hennes döttrar hava icke gjort vad du och dina döttrar haven gjort.
Se, detta var din syster Sodoms missgärning: fastän höghet, överflöd och tryggad ro hade blivit henne och hennes döttrar beskärd, understödde hon likväl icke den arme och fattige.
Tvärtom blevo de högfärdiga och bedrevo vad styggeligt var inför mig; därför försköt jag dem, när jag såg detta.
Ej heller Samaria har syndat hälften så mycket som du.
Du har gjort så många flera styggelser än dessa, att du genom alla de styggelser du har bedrivit har kommit dina systrar att synas rättfärdiga.
Så må också du nu bara din skam, du som nu kan lända dina systrar till ursäkt; ty därigenom att du har bedrivit ännu vederstyggligare synder än de, stå nu såsom rättfärdiga i jämförelse med dig.
Ja, blygs och bär din skam över att du så har kommit dina systrar att synas rättfärdiga.
Därför skall jag ock åter upp rätta dem, Sodom med hennes döttrar och Samaria med hennes döttrar.
Dig skall jag ock åter upprätta mitt ibland dem,
för att du må bära din skam och skämmas för allt vad du har gjort, och därmed bliva dem till tröst.
Och med dina systrar skall så ske: Sodom och hennes döttrar skola åter bliva vad de fordom voro, och Samaria och hennes döttrar skola åter bliva vad de fordom voro Också du själv och dina döttrar skolen åter bliva vad I fordom voren.
Men om du förr icke ens hördes nämna din syster Sodom, under din höghetstid,
innan ännu din egen ondska hade blivit uppenbarad -- såsom den blev på den tid då du vart till smälek för Arams döttrar och för alla de kringboende filistéernas döttrar, som hånade dig på alla sidor --
Så måste du nu själv bära på din skändlighet och dina styggelser, säger HERREN.
Ty så säger Herren, HERREN: Jag har handlat med dig efter dina gärningar, ty du hade ju föraktat eden och brutit förbundet.
Men jag vill nu tänka på det förbund som jag slöt med dig i din ungdoms dagar, och upprätta med dig ett evigt förbund.
Då skall du tänka tillbaka på dina vägar och skämmas, när du får taga till dig dina systrar, de större jämte de mindre; ty jag skall giva dem åt dig till döttrar, dock icke för din trohet i förbundet.
Men jag skall upprätta mitt förbund med dig, och du skall förnimma att jag är HERREN;
och så skall du tänka därpå och blygas, så att du av skam icke mer kan upplåta din mun, då när jag förlåter dig allt vad du har gjort, säger Herren, HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn, förelägg Israels hus en gåta, och tala till det en liknelse;
säg: Så säger Herren, HERREN: Den stora örnen med de stora vingarna och de långa pennorna, han som är så full med brokiga fjädrar, han kom till Libanon och tog bort toppen på cedern.
Han bröt av dess översta kvist och förde den till krämarlandet och satte den i en köpmansstad.
Sedan tog han en telning som växte i landet och planterade den i fruktbar jordmån; han tog den och satte den bland pilträd, på ett ställe där mycket vatten fanns.
Och den fick växa upp och bliva ett utgrenat vinträd, dock med låg stam, för att dess rankor skulle vända sig till honom och dess rötter vara under honom.
Den blev alltså ett vinträd som bar grenar och sköt skott.
Men där var ock en annan stor örn med stora vingar och fjädrar i mängd; och se, till denne böjde nu vinträdet längtansfullt sina grenar, och från platsen där det var planterat sträckte det sina rankor mot honom, för att han skulle vattna det.
Och dock var det planterat i god jordmån, på ett ställe där mycket vatten fanns, så att det kunde få grenar och bära frukt och bliva ett härligt vinträd.
Säg vidare: Så säger Herren, HERREN: Kan det nu gå det väl?
Skall man icke rycka upp dess rötter och riva av dess frukt, så att det förtorkar, och så att alla blad som hava vuxit ut därpå förtorka?
Och sedan skall varken stor kraft eller mycket folk behövas för att flytta det bort ifrån dess rötter.
Visst står det fast planterat, men kan det gå det väl?
Skall det icke alldeles förtorka, när östanvinden når det, ja, förtorka på den plats där det har vuxit upp?
Och HERRENS ord kom till mig, han sade:
Säg till det gensträviga släktet Förstån I icke vad detta betyder?
Så säg då: Se, konungen i Babel kom till Jerusalem och tog dess konung och dess furstar och hämtade dem till sig i Babel.
Och han tog en ättling av konungahuset och slöt förbund med honom och lät honom anlägga ed.
Men de mäktige i landet hade han fört bort med sig,
för att landet skulle bliva ett oansenligt rike, som icke kunde uppresa sig, och som skulle nödgas hålla förbundet med honom, om det ville bestå.
Men han avföll från honom och skickade sina sändebud till Egypten, för att man där skulle giva honom hästar och mycket folk.
Kan det gå den väl, som så gör?
Kan han undkomma?
Kan den som bryter förbund undkomma?
Så sant jag lever, säger Herren, HERREN: där den konung bor, som gjorde honom till konung, den vilkens ed han likväl föraktade, och vilkens förbund han bröt, där, hos honom i Babel, skall han sannerligen dö.
Och Farao skall icke med stor härsmakt och mycket folk bistå honom i kriget, när en vall kastas upp och en belägringsmur bygges, till undergång för många människor.
Eftersom han föraktade eden och bröt förbundet och gjorde allt detta fastän han hade givit sitt löfte, därför skall han icke undkomma.
Ja, därför säger Herren, HERREN så: Så sant jag lever, jag skall förvisso låta min ed, som han har föraktat, och mitt förbund, som han har brutit, komma över hans huvud.
Och jag skall breda ut mitt nät över honom, och han skall bliva fångad i min snara; och jag skall föra honom till Babel och där hålla dom över honom, för den otrohets skull som han har begått mot mig.
Och alla flyktingar ur alla hans härskaror skola falla för svärd, och om några bliva räddade, så skola de varda förströdda åt alla väderstreck.
Och I skolen förnimma att jag, HERREN, har talat.
Så säger Herren, HERREN: Jag vill ock själv taga en kvist av toppen på den höga cedern och sätta den; av dess översta skott skall jag avbryta en späd kvist och själv plantera den på ett högt och brant berg.
På Israels stolta berg skall jag plantera den, och den skall bära grenar och få frukt och bliva en härlig ceder.
Och allt vad fåglar heter av alla slag skall bo under den; de skola bo i skuggan av dess grenar.
Och alla träd på marken skola förnimma att det är jag, HERREN, som förödmjukar höga träd och upphöjer låga träd, som låter friska träd förtorka och gör torra träd grönskande.
Jag, HERREN, har talat det, och jag fullbordar det också.
Och HERRENS ord kom till mig; han sade:
Vad orsak haven I till att bruka detta ordspråk i Israels land: »Fäderna äta sura druvor, och barnens tänder bliva ömma därav»?
Så sant jag lever, säger Herren, HERREN, I skolen ingen orsak mer hava att bruka detta ordspråk i Israel.
Se, alla själar äro mina, faderns själ såväl som sonens är min; den som syndar, han skall dö.
Om nu en man är rättfärdig och övar rätt och rättfärdighet,
om han icke håller offermåltid på bergen, ej heller upplyfter sina ögon till Israels hus' eländiga avgudar, om han icke skändar sin nästas hustru, ej heller kommer vid en kvinna under hennes orenhets tid,
om han icke förtrycker någon, utan giver tillbaka den pant han har fått för skuld, om han icke tager rov, utan giver sitt bröd åt den hungrige och kläder den nakne,
om han icke ockrar eller tager ränta, om han håller sin hand tillbaka från vad orätt är och fäller rätta domar människor emellan --
ja, om han så vandrar efter mina stadgar och håller mina rätter, i det att han gör vad redligt är, då är han rättfärdig och skall förvisso få leva, säger Herren, HERREN.
Men om han så föder en son som bliver en våldsverkare, vilken utgjuter blod eller gör allenast något av allt detta
som han själv icke gjorde, en som håller offermåltid på bergen, skändar sin nästas hustru,
förtrycker den arme och fattige, tager rov, icke giver pant tillbaka, upplyfter sina ögon till de eländiga avgudarna, bedriver vad styggeligt är,
ockrar och tager ränta -- skulle då denne få leva?
Nej, han skall icke få leva, utan eftersom han bedriver sådana styggelser, skall han straffas med döden; hans blod skall komma över honom.
Och om sedan denne föder en son, vilken ser alla de synder som hans fader begår, och vid åsynen av dem själv tager sig till vara för att göra sådant,
en som icke håller offermåltid på bergen, icke upplyfter sina ögon till Israels hus' eländiga avgudar, icke skändar sin nästas hustru,
en som icke förtrycker någon, icke fordrar pant eller tager rov, utan giver sitt bröd åt den hungrige och kläder den nakne,
en som icke förgriper sig på den arme, ej heller ockrar eller tager ränta, utan gör efter mina rätter och vandrar efter mina stadgar, då skall denne icke dö genom sin faders missgärning, utan skall förvisso få leva.
Hans fader däremot, som begick våldsgärningar och rövade från sin broder och gjorde bland sina fränder det som icke var gott, se, han måste dö genom sin missgärning.
Huru kunnen I nu fråga: »Varför skulle icke sonen bära på sin faders missgärning?»
Jo, sonen övade ju rätt och rättfärdighet och höll alla mina stadgar och gjorde efter dem; därför skall han förvisso få leva.
Den som syndar, han skall dö; en son skall icke bära på sin faders missgärning, och en fader skall icke bära på sin sons missgärning.
Över den rättfärdige skall hans rättfärdighet komma, och över den ogudaktige skall hans ogudaktighet komma.
Men om den ogudaktige omvänder sig från alla de synder som han har begått, och håller alla mina stadgar och övar rätt och rättfärdighet, då skall han förvisso leva och icke dö.
Ingen av de överträdelser han har begått skall du tillräknas honom; genom den rättfärdighet han har övat skall han få leva.
Menar du att jag har lust till den ogudaktiges död, säger Herren, HERREN, och icke fastmer därtill att han vänder om från sin väg och får leva?
Men om den rättfärdige vänder om från sin rättfärdighet och gör vad orätt är, alla sådana styggelser som den ogudaktige gör -- skulle han då få leva, om han gör så?
Nej, intet av all den rättfärdighet han har övat skall då ihågkommas, utan genom den otrohet han har begått och den synd han har övat skall han dö.
Men nu sägen I: »Herrens väg är icke alltid densamma.»
Hören då, I av Israels hus: Skulle verkligen min väg icke alltid vara densamma?
Är det icke fastmer eder väg som icke alltid är densamma?
Om den rättfärdige vänder om från sin rättfärdighet och gör vad orätt är, så måste han dö till straff därför; genom det orätta som han gör måste han dö.
Men om den ogudaktige vänder om från den ogudaktighet som han har övat, och i stället övar rätt och rättfärdighet, då får han behålla sin själ vid liv.
Ja, eftersom han kom till insikt och vände om från alla de överträdelser han hade begått, skall han förvisso leva och icke dö.
Och ändå säga de av Israels hus: »Herrens väg är icke alltid densamma»!
Skulle verkligen mina vägar icke alltid vara desamma, I av Israels hus?
Är det icke fastmer eder väg som icke alltid är densamma?
Alltså: jag skall döma var och en av eder efter hans vägar, I av Israels hus, säger Herren, HERREN.
Vänden om, ja, vänden eder bort ifrån alla edra överträdelser, för att eder missgärning icke må bliva eder till en stötesten.
Kasten bort ifrån eder alla de överträdelser som I haven begått, och skaffen eder ett nytt hjärta och en ny ande; ty icke viljen I väl dö, I av Israels hus?
Jag har ju ingen lust till någons död, säger Herren HERREN.
Omvänden eder därför, så fån I leva.
Men du, stäm upp en klagosång över Israels furstar;
säg: Huru var icke din moder en lejoninna!
Bland lejon låg hon; hon födde upp sina ungar bland kraftiga lejon.
Så födde hon upp en av sina ungar, så att han blev ett kraftigt lejon; han lärde sig att taga rov, människor åt han upp.
Men folken fingo höra om honom och han blev fångad i deras grop; och man förde honom med krok i nosen till Egyptens land.
När hon nu såg att hon fick vänta förgäves, och att hennes hopp blev om intet, då tog hon en annan av sina ungar och gjorde denne till ett kraftigt lejon.
Stolt gick han omkring bland lejonen, ja, han blev ett kraftigt lejon; han lärde sig att taga rov, människor åt han upp.
Han våldförde deras änkor, deras städer förödde han.
Och landet med vad däri var blev förfärat vid dånet av hans rytande.
Då bådade man upp folk mot honom runt omkring från länderna; och de bredde ut sitt nät för honom, och han blev fångad i deras grop
Sedan satte de honom i en bur, med krok i nosen, och förde honom till konungen Babel Där satte man honom in i fasta borgar, för att hans röst ej mer skulle höras bort till Israels berg.
Medan de levde i ro, var din moder såsom ett vinträd, planterat vid vatten.
Och det blev ett fruktsamt träd, rikt på skott, genom det myckna vattnet.
Det fick starka grenar, tjänliga till härskarspiror, och dess stam växte hög, omgiven av lövverk, så att det syntes vida, ty det var högt och rikt på rankor.
Då ryckte man upp det i vrede, och det blev kastat på jorden, och stormen från öster förtorkade dess frukt.
Dess starka grenar brötos av och torkade bort, elden fick förtära dem.
Nu är det utplanterat i öknen, i ett torrt och törstande land.
Och eld har gått ut från dess yppersta gren och har förtärt dess frukt.
Så finnes där nu ingen stark gren kvar, ingen härskarspira!
En klagosång är detta, och den har fått tjäna såsom klagosång.
I sjunde året, på tionde dagen i femte månaden, kommo några av de äldste i Israel för att fråga HERREN; och de satte sig ned hos mig.
Då kom HERRENS ord till mig han sade:
Du människobarn, tala med de äldste i Israel och säg till dem: Så säger Herren, HERREN: Haven I kommit för att fråga mig?
Så sant jag lever, jag låter icke fråga mig av eder, säger Herren, HERREN.
Men vill du döma dem, ja, vill du döma, du människobarn, så förehåll dem deras fäders styggelser
och säg till dem: Så säger Herren, HERREN: På den dag då jag utvalde Israel, då upplyfte jag min hand till ed inför Jakobs hus' barn och gjorde mig känd för dem i Egyptens land; jag upplyfte min hand till ed inför dem och sade: »Jag är HERREN, eder Gud.
På den dagen lovade jag dem med upplyft hand att föra dem ut ur Egyptens land, till det land som jag hade utsett åt dem, ett land som skulle flyta av mjölk och honung, och som vore härligast bland alla länder.
Och jag sade till dem: »Var och en av eder kaste bort sina ögons styggelser, och ingen orene sig på Egyptens eländiga avgudar; jag är HERREN, eder Gud.»
Men de voro gensträviga mot mig och ville icke höra på mig; de kastade icke bort var och en sina ögons styggelser, och de övergåvo icke Egyptens eländiga avgudar.
Då tänkte jag på att utgjuta min förtörnelse över dem och att uttömma min vrede på dem mitt i Egyptens land.
Men vad jag gjorde, det gjorde jag för mitt namns skull, för att detta icke skulle bliva vanärat i de folks ögon, bland vilka de levde, och i vilkas åsyn jag gjorde mig känd för dem, i det jag förde dem ut ur Egyptens land.
Så förde jag dem då ut ur Egyptens land och lät dem komma in i öknen.
Och jag gav dem mina stadgar och kungjorde för dem mina rätter; den människa som gör efter dem får leva genom dem.
Jag gav dem ock mina sabbater, till att vara ett tecken mellan mig och dem, för att man skulle veta att jag är HERREN, som helgar dem.
Men Israels hus var gensträvigt mot mig i öknen; de vandrade icke efter mina stadgar, utan föraktade mina rätter, fastän den människa som gör efter dem får leva genom dem; de ohelgade ock svårt mina sabbater.
Då tänkte jag på att utgjuta min förtörnelse över dem i öknen och så förgöra dem.
Men vad jag gjorde, det gjorde jag för mitt namns skull, för att detta icke skulle bliva vanärat i de folks ögon, i vilkas åsyn jag hade fört dem ut.
Likväl upplyfte jag min hand inför dem i öknen och svor att jag icke skulle låta dem komma in i det land som jag hade givit dem, ett land som skulle flyta av mjölk och honung, och som vore härligast bland alla länder --
detta därför att de föraktade mina rätter och icke vandrade efter mina stadgar, utan ohelgade mina sabbater, i det att deras hjärtan följde efter deras eländiga avgudar.
Men jag visade dem skonsamhet och fördärvade dem icke; jag gjorde icke alldeles ände på dem i öknen.
Och jag sade till deras barn i öknen: »I skolen icke vandra efter edra fäders stadgar och icke hålla deras rätter, ej heller orena eder på deras eländiga avgudar.
Jag är HERREN, eder Gud; vandren efter mina stadgar och håller mina rätter och gören efter dem.
Och helgen mina sabbater, och må de vara ett tecken mellan mig och eder, för att man må veta att jag är HERREN, eder Gud.
Men deras barn voro gensträviga mot mig; de vandrade icke efter mina stadgar och höllo icke mina rätter, så att de gjorde efter dem fastän den människa som gör efter dem får leva genom dem; de ohelgade ock mina sabbater.
Då tänkte jag på att utgjuta min förtörnelse över dem och att uttömma min vrede på dem i öknen.
Men jag drog min hand tillbaka, och vad jag gjorde, det gjorde jag för mitt namns skull, för att detta icke skulle bliva vanärat i de folks ögon, i vilkas åsyn jag hade fört dem ut.
Likväl upplyfte jag min hand inför dem i öknen och svor att förskingra dem bland folken och förströ dem i länderna,
eftersom de icke gjorde efter mina rätter, utan föraktade mina stadgar och ohelgade mina sabbater, och eftersom deras ögon hängde vid deras fäders eländiga avgudar.
Därför gav jag dem ock stadgar som icke voro till deras båtnad, och rätter genom vilka de icke kunde bliva vid liv.
Och jag lät dem orena sig med sina offerskänker, med att låta allt som öppnade moderlivet gå genom eld, ty jag ville slå dem med förfäran, på det att de skulle förstå att jag är HERREN.
Tala därför till Israels hus, du människobarn, och säg till dem: Så säger Herren, HERREN: Också därmed hava edra fäder hädat mig, att de hava begått otrohet mot mig.
När jag hade låtit dem komma in i det land som jag med upplyft hand hade lovat att giva dem, och när de så där fingo se någon hög kulle eller något lummigt träd, då offrade de där sina slaktoffer och framburo där sina offergåvor, mig till förtörnelse, och läto där sina offers välbehagliga lukt uppstiga och utgöto där sina drickoffer.
Då sade jag till dem: »Vad är detta för en offerhöjd, denna som I kommen till?»
Därav fick en sådan plats namnet »offerhöjd», såsom man säger ännu i dag.
Säg därför till Israels hus: Så säger Herren, HERREN: Skolen då I orena eder på samma sätt som edra fäder gjorde, och i trolös avfällighet löpa efter deras styggelser?
I orenen eder ännu i dag på alla edra eländiga avgudar, i det att I frambären åt dem edra offerskänker och låten edra barn gå genom eld.
Skulle jag då låta fråga mig av eder, I av Israels hus?
Nej, så sant jag lever, säger Herren, HERREN, ja låter icke fråga mig av eder.
Och förvisso skall icke det få ske som har kommit eder i sinnet, då I tänken: »Vi vilja bliva såsom hedningarna, såsom folken i andra länder: vi vilja tjäna trä och sten.
Så sant jag lever, säger Herren, HERREN, med stark hand och uträckt arm och utgjuten förtörnelse skall jag sannerligen regera över eder.
Och med stark hand och uträckt arm och utgjuten förtörnelse skall jag föra eder ut ifrån folken och församla eder från de länder i vilka I ären förströdda.
Och jag skall föra eder in i Folkens öken, och där skall jag gå till rätta med eder, ansikte mot ansikte.
Likasom jag gick till rätta med edra fäder i öknen vid Egyptens land, så skall jag ock gå till rätta med eder, säger Herren, HERREN.
Och jag skall låta eder draga fram under staven och tvinga eder in i förbundets band.
Och jag skall rensa bort ifrån eder dem som sätta sig upp emot mig och avfalla från mig, jag skall skaffa bort dem ur det land där de nu bo, men in i Israels land skola de icke få komma; och I skolen förnimma att jag är HERREN.
Men hören nu, I av Israels hus: Så säger Herren, HERREN: Välan, gån åstad och tjänen edra eländiga avgudar, var och en dem han har.
Sedan skolen I förvisso komma att höra på mig, och I skolen då icke mer ohelga mitt heliga namn med edra offerskänker och edra eländiga avgudar.
Ty på mitt heliga berg, på Israels höga berg, säger Herren, HERREN där skall hela Israels hus tjäna mig, så många därav som finnas i landet; där skall jag finna behag i dem, där skall jag hava lust till edra offergärder och till förstlingen av edra gåvor, vadhelst I viljen helga.
Vid den välbehagliga lukten skall jag finna behag i eder, när tiden kommer, att jag för eder ut ifrån folken och församlar eder från de länder i vilka I ären förströdda.
Och jag skall bevisa mig helig på eder inför folkens ögon.
Ja, I skolen förnimma att jag är HERREN, när jag låter eder komma in i Israels land, det land som jag med upplyft hand lovade att giva åt edra fäder.
Och där skolen I tänka tillbaka på edra vägar och på alla de gärningar som I orenaden eder med; och I skolen känna leda vid eder själva för allt det onda som I haven gjort.
Och I skolen förnimma att jag är HERREN, när jag så handlar med eder, för mitt namns skull och icke efter edra onda vägar och edra skändliga gärningar, I av Israels hus, säger Herren, HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn, vänd ditt ansikte söderut och predika mot söder; ja, profetera mot skogslandet söderut;
säg till skogen söderut: Hör HERRENS ord: Så säger Herren, HERREN: Se, jag skall tända upp en eld i dig, och den skall förtära alla träd i dig, både de friska och de torra; den flammande lågan skall icke kunna släckas, och av den skola allas ansikten förbrännas, allas mellan söder och norr.
Och allt kött skall se att jag, HERREN, har upptänt den; den skall icke kunna släckas.
Och jag sade: »Ack, Herre, HERRE!
Dessa säga om mig: 'Denne talar ju gåtor.'»
Och HERRENS ord kom till mig; han sade:
Du människobarn, vänd ditt ansikte mot Jerusalem och predika mot helgedomarna, ja, profetera mot Israels land.
Och säg till Israels land: Så säger HERREN: Se, jag skall vända mig mot dig och draga ut mitt svärd ur skidan och utrota ur dig både rättfärdiga och ogudaktiga.
Ja, eftersom jag skall utrota ur dig både rättfärdiga och ogudaktiga, därför skall mitt svärd fara ut ur skidan och vända sig mot allt kött mellan söder och norr;
och allt kött skall förnimma att jag, HERREN, har dragit ut mitt svärd ur skidan; det skall icke mer stickas in igen.
Men du, människobarn, må sucka, ja, du må sucka inför deras ögon, som om dina länder skulle brista sönder i din bittra smärta.
Och när de fråga dig: »Varför suckar du?», då skall du svara: »För ett olycksbud, som när det kommer, skall göra att alla hjärtan förfäras och alla händer sjunka ned och alla sinnen omtöcknas och alla knän bliva såsom vatten.
Se, det kommer, ja, det fullbordas! säger Herren, HERREN.»
Och HERRENS ord kom till mig; han sade:
Du människobarn, profetera och säg: Så säger HERREN: Säg: Ett svärd, ja, ett svärd har blivit vässt och har blivit fejat.
Det har blivit vässt, för att det skall anställa ett slaktande; det har blivit fejat, för att det skall blixtra.
Eller skola vi få fröjd därav?
Fröjd av det som bliver ett tuktoris för min son, ett för vilket intet trä kan bestå!
Nej, han har lämnat det till att fejas, för att det skall fattas i handen; svärdet har blivit vässt och fejat för att sättas i en dråpares hand.
Ropa och jämra dig, du människobarn, ty det drabbar mitt folk, det drabbar alla Israels hövdingar.
De äro med mitt folk hemfallna åt svärdet; därför må du slå dig på länden.
Ty rannsakning har redan skett; huru skulle det då vara möjligt att riset icke drabbade, det ris för vilket intet kan bestå? säger Herren, HERREN.
Men du, människobarn, profetera och slå händerna tillsammans; må svärdet fördubblas, ja, bliva såsom tre, må det bliva ett mordsvärd, ett mordsvärd jämväl för den störste, svärdet som drabbar dem från alla håll.
Ja, för att deras hjärtan må försmälta av ångest, och för att många må falla, skall jag sända det blänkande svärdet mot alla deras portar.
Ack, det är gjort likt en blixt, det är draget för att slakta!
Hugg lös med all makt åt höger, måtta åt vänster, varthelst din egg kan bliva riktad.
Också jag skall slå mina händer tillsammans och släcka min vrede.
Jag, HERREN, har talat.
Och HERRENS ord kom till mig; han sade:
Du människobarn, märk ut åt dig två vägar på vilka den babyloniske konungens svärd kan gå fram; låt båda gå ut från ett och samma land.
Skär så ut en vägvisare, skär ut den för den plats där stadsvägarna skilja sig.
Märk ut såsom det håll dit svärdet kan gå dels Rabba i Ammons barns land, dels Juda med det befästa Jerusalem.
Ty konungen i Babel står redan vid vägskälet där de båda vägarna begynna; han vill låta spå åt sig, han skakar pilarna, han rådfrågar sina husgudar, han ser på levern.
I sin högra hand får han då ut lotten »Jerusalem», för att han där skall sätta upp murbräckor, öppna sin mun till krigsrop, upphäva sin röst till härskri, för att han där skall sätta upp murbräckor mot portarna, kasta upp en vall och bygga en belägringsmur. --
Detta synes dem vara en falsk spådom: de hava ju heliga eder.
Men han uppväcker minnet av deras missgärning, och så ryckas de bort.
Därför säger Herren, HERREN så: Eftersom I haven uppväckt minnet av eder missgärning i det att edra överträdelser hava blivit uppenbara, så att eder syndfullhet visar sig i allt vad I gören, ja, eftersom minnet av eder har blivit uppväckt, därför skolen I komma att med makt ryckas bort.
Och du, dödsdömde, ogudaktige furste över Israel, du vilkens dag kommer, när din missgärning har nått sin gräns,
så säger Herren, HERREN: Tag av dig huvudbindeln, lyft av dig kronan.
Det som nu är skall icke förbliva vad det är; vad lågt är skall upphöjas, och vad högt är skall förödmjukas.
Omstörtas, omstörtas, omstörtas skall detta av mig; också detta skall vara utan bestånd, till dess han kommer, som har rätt därtill, den som jag har givit det åt.
Och du, människobarn, profetera Och såg: Så säger Herren, HERREN om Ammons barn och om deras smädelser: Säg: Ett svärd, ja, ett svärd är draget, det är fejat för att slakta för att varda mättat och för att blixtra,
mitt under det att man skådar åt dig falska profetsyner och spår åt dig lögnaktiga spådomar om att du skall sättas på de dödsdömda ogudaktigas hals, vilkas dag kommer, när missgärningen har nått sin gräns.
Må det stickas i skidan igen.
I den trakt där du är skapad, i det land varifrån du stammar, där skall jag döma dig.
Jag skall Utgjuta min vrede över dig, jag skall mot dig blåsa upp min förgrymmelses eld; och jag skall giva dig till pris åt vilda människor, åt män som äro mästare i att fördärva.
Du skall bliva till mat åt elden, ditt blod skall flyta i landet; ingen skall mer tänka på dig.
Ty jag, HERREN, har talat.
Och HERRENS ord kom till mig; han sade:
Du människobarn, vill du döma ja, vill du döma blodstaden?
Förehåll henne då alla hennes styggelser
och säg: Så säger Herren, HERREN: Du stad som utgjuter dina invånares blod, så att din stund måste komma, du som gör eländiga avgudar åt dig och så bliver orenad!
Genom det blod som du har utgjutit har du ådragit dig skuld, och genom de eländiga avgudar som du har gjort har du orenat dig; så har du påskyndat dina dagars slut och nu hunnit gränsen för dina år.
Därför skall jag låta dig bliva till smälek för folken och till spott för alla länder.
Ja, både nära och fjärran skall man bespotta dig, du vilkens namn är skändat, du förvirringens stad.
Se, hos dig trotsa Israels hövdingar var och en på sin arm, om det gäller att utgjuta blod.
Över fader och moder uttalar man förbannelser hos dig; mot främlingen övar man våld hos dig; den faderlöse och änkan förtrycker man hos dig.
Mina heliga ting föraktar du, och mina sabbater ohelgar du.
Förtalare finnas hos dig, om det gäller att utgjuta blod.
Man håller hos dig offermåltider på bergen; man bedriver hos dig vad skändligt är.
Man blottar sin faders blygd hos dig; man kränker hos dig kvinnan, när hon har sin orenhets tid.
Man bedriver styggelse, var och en med sin nästas hustru; ja, man orenar i skändlighet sin sons hustru; man kränker hos dig sin syster, sin faders dotter.
Man tager hos dig mutor för att utgjuta blod; ja, du ockrar och tager ränta och skinnar din nästa med våld, och mig förgäter du, säger Herren, HERREN.
Men se, jag slår mina händer tillsammans i harm över det skinneri du övar, och i harm över det blod som du utgjuter hos dig.
Menar du att ditt mod skall bestå, eller att dina händer skola vara starka nog, när tiden kommer, att jag utför mitt verk på dig?
Jag HERREN, har talat, och jag fullbordar det också.
Jag skall förskingra dig bland folken och förströ dig i länderna; så skall jag taga bort ifrån dig all din orenhet.
Du skall bliva vanärad inför folkens ögon, genom din egen skuld; och du skall förnimma att jag är HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn, Israels hus har för mig blivit slagg; de äro allasammans blott koppar, tenn, järn och bly i ugnen; de äro ett silver som kan räknas för slagg.
Därför säger Herren, HERREN så: Eftersom I allasammans haven blivit slagg, se, därför skall jag hopsamla eder i Jerusalem.
Likasom man hopsamlar silver, koppar, järn, bly och tenn i ugnen och där blåser upp eld under det och smälter det, så skall jag i min vrede och förtörnelse hopsamla eder och kasta eder i ugnen och smälta eder.
Ja, jag skall samla eder tillhopa; och blåsa upp min förgrymmelses eld under eder, för att I man smältas däri.
Likasom silver smältes i ugnen, så skolen I smältas däri; och I skolen förnimma att det är jag, HERREN, som utgjuter min förtörnelse över eder.
Och HERRENS ord kom till mig; han sade: Du människobarn, säg till dem:
Du är ett land som icke bliver renat, icke varder sköljt av regn på vredens dag.
De profeter som där finnas hava sammansvurit sig och blivit såsom rytande, rovgiriga lejon; de äta upp själar, de riva till sig gods och dyrbarheter och göra många till änkor därinne.
Prästerna där våldföra min lag och ohelga mina heliga ting; de göra ingen åtskillnad mellan heligt och oheligt och undervisa icke om skillnaden mellan rent och orent.
De tillsluta sina ögon för mina sabbater, och så bliver jag ohelgad mitt ibland dem.
Furstarna därinne äro såsom rovgiriga vargar; de utgjuta blod och förgöra själar för att skaffa sig vinning.
De profeter som de hava tjäna dem såsom vitmenare; de skåda åt dem falska profetsyner och spå åt dem lögnaktiga spådomar; de säga: »Så säger Herren, HERREN», och det fastän HERREN icke har talat.
Folket i landet begår våldsgärningar och tager rov; den arme och fattige förtrycka de, och mot främlingen öva de våld, utan lag och rätt.
Jag söker bland dem efter någon som skulle kunna uppföra en mur och träda fram i gapet inför mig till försvar för landet, på det att jag icke må fördärva det; men jag finner ingen.
Därför utgjuter jag min vrede över dem och gör ände på dem med min förgrymmelses eld.
Deras gärningar skall jag låta komma över deras huvuden, säger Herren, HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn, det var en gång två kvinnor, döttrar till en och samma moder.
Dessa bedrevo otukt i Egypten; de gjorde det redan i sin ungdom.
Där kramades deras bröst, och där smekte man deras jungfruliga barm.
Den äldre hette Ohola, och hennes syster Oholiba.
Därefter blevo de mina, och födde söner och döttrar.
Och om deras namn är att veta att Ohola är Samaria, och Oholiba Jerusalem.
Men Ohola bedrev otukt i stället för att hålla sig till mig; hon upptändes av lusta till sina älskare hennes grannar assyrierna,
där de kommo klädda i mörkblå purpur och voro ståthållare och landshövdingar, vackra unga män allasammans, ryttare som redo på hästar.
Hon gav åt dem sin trolösa älskog, åt Assurs alla yppersta söner; och varhelst hon upptändes av lusta, där orenade hon sig på alla deras eländiga avgudar
Men ändå uppgav hon icke sin otukt med egyptierna, som hade fått ligga hos henne i hennes ungdom, och som hade smekt hennes jungfruliga barm och slösat på henne sin otukt.
Därför gav jag henne till pris åt hennes älskare, åt Assurs söner, till vilka hon var upptänd av lusta.
Och sedan dessa hade blottat hennes blygd, förde de bort hennes söner och döttrar och dräpte henne själv med svärd; så blev hon en varnagel för andra kvinnor, då nu dom blev hållen över henne.
Men fastän hennes syster Oholiba såg detta, upptändes hon av lusta ännu värre och drev sin otukt ännu längre än systern.
Hon upptändes av lusta till Assurs söner; de voro ju ståthållare och landshövdingar och voro hennes grannar, de kommo klädda i präktig dräkt, ryttare som redo på hästar, vackra unga män allasammans.
Och jag såg att också hon orenade sig; båda gingo de samma väg.
Men denna drev sin otukt ännu längre.
Ty när hon fick se mansbilder inristade i väggen, beläten av kaldéer, som man hade inristat och målat röda med dyrbar färg,
framställda med gördlar kring sina länder och med ståtliga huvudbonader, allasammans lika kämpar, ja, när hon fick se dessa bilder av Babels söner, av de män som hade sitt fädernesland i Kaldeen;
då upptändes hon av lusta till dem, strax när hon såg dem för sina ögon.
Och hon sände bud till dem i Kaldeen;
och Babels söner kommo till henne och lågo hos henne i älskog och orenade henne genom sin otukt.
Först sedan hon hade blivit orenad av dem, vände sig hennes själ ifrån dem.
Men när hon så öppet bedrev sin otukt och blottade sin blygd, då vände sig min själ ifrån henne, likasom den hade vänt sig ifrån hennes syster.
Dock drev hon sin otukt ännu längre: hon mindes sin ungdoms dagar, då hon bedrev otukt i Egyptens land;
och så upptändes hon åter av lusta till bolarna där, som hade kött såsom åsnor och flöde såsom hästar.
Ja, din håg stod åter till din ungdoms skändlighet, när egyptierna smekte din barm, därför att du hade så ungdomliga bröst.
Därför, du Oholiba, säger Herren, HERREN så: Se, jag skall uppväcka mot dig dina älskare, dem som din själ har vänt sig ifrån, och jag skall låta dem komma över dig från alla sidor,
Babels söner och alla kaldéer, pekodéer, soéer och koéer och alla Assurs söner med dem, vackra unga män, ståthållare och landshövdingar allasammans, kämpar och berömliga män, som rida på hästar allasammans.
De skola komma över dig med vagnar och hjuldon i mängd och med skaror av folk; rustade med skärmar och sköldar och klädda hjälmar skola de anfalla dig från alla sidor.
Och jag skall överlämna domen åt dem, och de skola döma dig efter sina rätter.
Jag skall låta min nitälskan gå över dig, så att de fara grymt fram mot dig; de skola skära av dig näsa och öron, och de som bliva kvar av dig skola falla för svärd.
Man skall föra bort dina söner och döttrar, och vad som bliver kvar av dig skall förtäras av eld.
Man skall slita av dig dina kläder och taga ifrån dig dina härliga smycken.
Så skall jag göra slut på din skändlighet och på den otukt som du begynte öva i Egyptens land; och du skall icke mer lyfta upp dina ögon till dem och icke mer tänka på Egypten.
Ty så säger Herren, HERREN: Se, jag vill giva dig till pris åt dem som du nu hatar, åt dem som din själ har vänt sig bort ifrån.
Och de skola fara fram mot dig såsom fiender, och skola taga ifrån dig allt vad du har förvärvat och lämna dig naken och blottad; ja, din otuktiga blygd skall varda blottad, med din skändlighet och din otukt.
Detta skall man göra dig, därför att du i otukt lopp efter hedningarna och orenade dig på deras eländiga avgudar.
Du vandrade på din systers väg; därför skall jag sätta i din hand samma kalk som gavs åt henne.
Ja, så säger Herren, HERREN: Du skall nödgas dricka din systers kalk, så djup och så vid som den är, och den skall bringa dig åtlöje och smälek i fullt mått.
Du skall bliva drucken och bliva full av bedrövelse, ty en ödeläggelsens och förödelsens kalk är din syster Samarias kalk.
Du skall nödgas dricka ut den till sista droppen, ja ock slicka dess skärvor, och du skall sarga ditt bröst.
Ty jag har talat, säger Herren, HERREN.
Därför säger Herren, HERREN så: Eftersom du har förgätit mig och kastat mig bakom din rygg, därför måste du ock bära på din skändlighet och din otukt.
Och HERREN sade till mig: Du människobarn, vill du döma Ohola och Oholiba?
Förehåll dem då deras styggelser.
Ty de hava begått äktenskapsbrott, och blod låder vid deras händer.
Ja, med sina eländiga avgudar hava de begått äktenskapsbrott; och till mat åt dem hava de offrat sina barn, dem som de hade fött åt mig.
Därtill gjorde de mig detta: samma dag som de orenade min helgedom ohelgade de ock mina sabbater.
Ty samma dag som de slaktade sina barn åt de eländiga avgudarna gingo de in i min helgedom och ohelgade den.
Se, sådant hava de gjort i mitt hus.
Än mer, de sände bud efter män som skulle komma fjärran ifrån; budbärare skickades till dem, och se, de kommo, de män för vilka du hade tvått dig och sminkat dina ögon och prytt dig med smycken.
Och du satt på en härlig vilobädd, med ett dukat bord framför, och du hade där ställt fram min rökelse och min olja.
Sorglöst larm hördes därinne, och till de män ur hopen, som voro där, hämtade man ytterligare in dryckesbröder från öknen.
Och dessa satte armband på kvinnornas armar och härliga kronor på deras huvuden.
Då sade jag: »Skall hon, den utlevade, få hålla i med att begå äktenskapsbrott?
Skall man alltjämt få bedriva otukt med henne, då hon är en sådan?»
Ty man gick in till henne, såsom man går in till en sköka; ja, så gick man in till Ohola och till Oholiba, de skändliga kvinnorna.
Men rättfärdiga man skola döma dem efter den lag som gäller för äktenskapsbryterskor och blodsutgjuterskor; ty äktenskapsbryterskor äro de, och blod låder vid deras händer.
Ja, så säger Herren, HERREN: Må man sammankalla en församling mot dem och prisgiva dem åt misshandling och plundring.
Och församlingen skall stena dem och hugga dem i stycken med svärd, och dräpa deras söner och döttrar, och bränna upp deras hus i eld.
Så skall jag göra slut på skändligheten i landet, och alla kvinnor må låta varna sig, så att de icke bedriva sådan skändlighet som I.
Och man skall låta eder skändlighet komma över eder, och I skolen få bära på de synder I haven begått med edra eländiga avgudar; och I skolen förnimma att jag är Herren, HERREN.
Och HERRENS ord kom till mig i nionde året, på tionde dagen i tionde månaden; han sade:
Du människobarn, skriv upp åt dig namnet på denna dag, just denna dag; ty konungen i Babel har på just denna dag ryckt fram mot Jerusalem.
Och tala till det gensträviga släktet i en liknelse; säg till dem: Så säger Herren, HERREN: Sätt på grytan, och när du har satt på den, så gjut vatten däri.
Lägg sedan köttstyckena tillhopa däri, allahanda goda stycken, av låret och bogen; och fyll den så med de bästa märgbenen.
Tag härtill det bästa av hjorden; och lägg bränsle under den för att koka benen.
Låt den koka starkt, så att ock benen bliva kokta i den.
Så säger nu Herren, HERREN: Ve över blodstaden, den rostiga grytan, varifrån rosten icke har kunnat tagas bort!
Det ena köttstycket efter det andra har man redan tagit ut därur, utan att kasta lott om ordningen.
Ty det blod hon har utgjutit är ännu kvar därinne; på kala klippan lät hon det rinna ned; hon utgöt det icke på sådan mark att mullen har kunnat skyla det.
För att vreden skulle hava sin gång, och för att jag skulle utkräva hämnd, lät jag det blod hon utgöt komma på kala klippan, där det icke kunde skylas.
Därför säger Herren, HERREN så: Ve över blodstaden!
Jag skall nu ytterligare öka på bränslet därunder.
Ja, lägg på mer ved, tänd upp eld, låt köttet bliva förstört och spadet koka in och benen bliva förbrända.
Och låt den sedan stå tom på eldsglöden, till dess att den bliver så upphettad att dess koppar glödgas och orenligheten smältes bort därur och rosten försvinner.
Tung möda har den kostat, och ändå har dess myckna rost icke gått bort.
Så må nu dess röst komma i elden!
Därför att din orenhet är så skändlig, och därför att du icke blev ren. huru jag än sökte rena dig, därför skall du nu icke mer bliva fri ifrån din orenhet, förrän jag har släckt min vrede på dig.
Jag, HERREN, har talat.
Det kommer!
Jag skall fullborda det!
Jag skall icke släppa efter och icke skona och icke ångra mig.
Efter dina vägar och dina gärningar skall man döma dig, säger Herren, HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn, se, genom en plötslig död skall jag taga ifrån dig den som är dina ögons lust, men du må icke hålla dödsklagan eller gråta eller fälla tårar.
Tyst må du jämra dig; men du skall icke hålla sorgefest såsom efter en död.
Nej, sätt på dig din huvudbindel och tag skor på dina fötter; skyl icke ditt skägg, och ät icke det särskilda bröd som eljest är övligt.
Sedan talade jag nästa morgon till folket, men på aftonen dog min hustru; och följande morgon gjorde jag såsom mig var befallt.
Då sade folket till mig: »Vill du icke omtala för oss vad det betyder att du så gör?»
Jag svarade dem: HERRENS ord kom till mig; han sade:
Säg till Israels hus: Så säger Herren, HERREN: Se, jag vill ohelga min helgedom, eder stolta härlighet, edra ögons lust och eder själs längtan.
Och edra söner och döttrar, som I haven måst övergiva, skola falla för svärd.
Då skolen I komma att göra såsom jag har gjort: I skolen icke skyla skägget och icke äta det övliga brödet.
Och I skolen behålla huvudbindlarna på edra huvuden och skorna på edra fötter; I skolen icke hålla dödsklagan eller gråta, utan skolen sitta där försmäktande genom edra missgärningar och sucka med varandra.
Hesekiel skall vara ett tecken för eder; alldeles såsom han gör skolen I komma att göra.
När detta händer, skolen I förnimma att jag är Herren, HERREN.
Men du, människobarn, må veta att på den tid då jag tager ifrån dem deras värn, deras härliga fröjd, deras ögons lust och deras själs begär, deras söner och döttrar,
på den tiden skall en räddad flykting komma till dig och förkunna detta.
Och då när flyktingen är där, skall din mun upplåtas, och du skall tala och icke mer vara stum; och du skall vara ett tecken för dem, och de skola förnimma att jag är HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn, vänd ditt an- sikte mot Ammons barn och profetera mot dem.
Och säg till Ammons barn: Hören Herrens, HERRENS ord: Så säger Herren, HERREN: Eftersom du ropar: »Rätt så!» över min helgedom, som har blivit oskärad, och över Israels land, som har blivit ödelagt, och över Juda folk, som har måst vandra bort i fångenskap,
se, därför vill jag giva dig till besittning åt österlänningarna, så att de få slå upp sina tältläger i dig och sätta upp sina boningar i dig; de skola få äta din frukt, och de skola dricka din mjölk.
Och jag skall göra Rabba till en betesmark för kameler och Ammons barns land till en lägerplats för får; och I skolen förnimma att Jag är HERREN.
Ty så säger Herren, HERREN: Eftersom du klappar i händerna och stampar med fötterna och i ditt sinnes hela övermod gläder dig vid Israels lands ofärd,
se, därför skall jag uträcka min hand mot dig och giva dig till byte åt hedningarna och utrota dig ifrån folken och utplåna dig ur länderna; jag skall förgöra dig, och du skall förnimma att jag är HERREN.
Så säger Herren, HERREN: Eftersom Moab och Seir säga: »Se, nu är det med Juda hus likasom med alla andra folk»,
se, därför skall jag lägga Moabs bergsluttning öppen och förstöra dess städer, Ja, dess städer så många de äro, vad härligast är i landet, Bet-Hajesimot, Baal-Meon och Kirjatama.
Åt österlänningarna skall jag giva det till besittning, likasom jag skall göra med Ammons barns land, så att man icke mer tänker på Ammons barn ibland folken.
Ja, över Moab skall jag hålla dom, och de skola förnimma att jag är HERREN.
Så säger Herren, HERREN: Eftersom Edom har handlat så hämndgirigt mot Juda hus och ådragit sig svår skuld genom sin hämnd på dem,
därför säger Herren, HERREN så: Jag skall uträcka min hand mot Edom och utrota därur både människor och djur.
Och jag skall göra det till en ödemark ända från Teman, och ända borta i Dedan skola de falla för svärd.
Och jag skall utföra min hämnd på Edom genom mitt folk Israel, och dessa skola göra med Edom efter min vrede och förtörnelse; och det skall så få känna min hämnd, säger Herren, HERREN.
Så säger Herren, HERREN: Eftersom filistéerna hava handlat så hämndgirigt, ja, eftersom de i sitt sinnes övermod hava velat utkräva hämnd och i sin eviga fiendskap hava velat bereda fördärv,
därför säger Herren, HERREN så: Se, jag vill uträcka min hand mot filistéerna och utrota keretéerna och förgöra vad som är kvar av Kustlandet vid havet.
Och jag skall taga stor hämnd på dem och tukta dem i förtörnelse.
Och när jag låter min hämnd drabba dem, då skola de förnimma att jag är HERREN.
Och i elfte året, på första dagen i månaden, kom HERRENS ord till mig; han sade:
Du människobarn, eftersom Tyrus sade om Jerusalem: »Rätt så, uppbruten är nu folkens port, den är öppnad för mig; jag bliver rik, nu då hon är förödd»,
därför säger Herren, HERREN så: Se, jag skall komma över dig, Tyrus, och jag skall upphäva många folk mot dig, likasom havet upphäver sina böljor.
De skola förstöra Tyrus' murar och riva ned dess torn.
Så skall jag sopa bort själva dess grus och förvandla staden till en kal klippa.
En torkplats för fisknät skall den vara ute i havet; ty jag har talat, säger Herren, HERREN.
Ja, den skall bliva ett byte för folken;
och dess döttrar på fastlandet skola dräpas med svärd.
De skola förnimma att jag är HERREN.
Ty så säger Herren, HERREN: Se, jag vill låta Nebukadressar, konungen i Babel, konungarnas konung, komma norrifrån över Tyrus, med hästar och vagnar och ryttare och med en stor hop folk.
Dina döttrar på fastlandet skall han dräpa med svärd; han skall bygga en belägringsmur mot dig och kasta upp mot dig en vall och resa ett sköldtak mot dig.
Sin murbräckas stötar skall han rikta mot dina murar och skall med sina krigsredskap bryta ned dina torn.
Hans hästar äro så många att dammet skall överhölja dig.
Vid dånet av hans ryttare och av hans hjuldon och vagnar skola dina murar darra, när han drager in genom dina portar, såsom man drager in i en erövrad stad.
Med sina hästars hovar skall han trampa sönder alla dina gator; ditt folk skall han dräpa med svärd, och dina stolta stoder skola störta till jorden.
Man skall röva dina skatter och plundra dina handelsvaror; man skall riva dina murar och bryta ned dina sköna hus; och stenarna, trävirket och gruset skall man kasta i havet.
Jag skall göra slut på dina sångers buller, och man skall icke mer höra klangen av dina harpor.
Ja, jag skall göra dig till en kal klippa en torkplats för fisknät skall du bliva; aldrig mer skall du varda uppbyggd.
Ty jag, HERREN, har talat, säger Herren, HERREN.
Så säger Herren, HERREN till Tyrus: Sannerligen, vid dånet av ditt fall, när de slagna jämra sig, vid det att man dräper och mördar i dig, skola havsländerna bäva.
Och alla hövdingar vid havet skola stiga ned från sina troner, de skola lägga bort sina mantlar och taga av sig sina brokigt vävda kläder; förskräckelse bliver deras klädnad, och nere på jorden skola de sitta; deras förskräckelse varder ständigt ny, och de häpna över ditt öde.
De stämma upp en klagosång över dig och säga om dig: Huru har du icke blivit förstörd, du havsfolkens tillhåll, du högtprisade stad, du som var så mäktig på havet, där du låg med dina invånare, vilka fyllde människorna med skräck för alla som bodde i dig!
Nu förskräckas havsländerna på ditt falls dag, och öarna i havet förfäras vid din undergång.
Ty så säger Herren, HERREN: När jag gör dig till en ödelagd stad, lik någon stad som ingen bebor, ja, när jag låter djupet upphäva sig mot dig och de stora vattnen betäcka dig,
då störtar jag dig ned till dem som hava farit ned i graven, till folk som levde för länge sedan; och lik en längesedan ödelagd plats får du ligga där i jordens djup, hos dem som hava farit ned i graven.
Så skall du förbliva obebodd, medan jag gör härliga ting i de levandes land.
Jag skall låta dig taga en ande med förskräckelse, så att man aldrig i evighet skall finna dig, huru man än söker efter dig, säger Herren, HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn, stäm upp en klagosång över Tyrus;
säg till Tyrus: Du som bor vid havets portar och driver köpenskap med folken, hän till många havsländer, så säger Herren, HERREN: O Tyrus, du säger själv: »Jag är skönhetens fullhet.»
Ja, dig som har ditt rike ute i havet, dig gjorde dina byggningsmän fullkomlig i skönhet.
Av cypress från Senir timrade de allt plankverk på dig; de hämtade en ceder från Libanon för att göra din mast.
Av ekar från Basan tillverkade de dina åror.
Ditt däck prydde de med elfenben i ädelt trä från kittéernas öländer.
Ditt segel var av fint linne, med brokig vävnad från Egypten, och det stod såsom ditt baner.
Mörkblått och purpurrött tyg från Elisas öländer hade du till soltält.
Sidons och Arvads invånare voro roddare åt dig; de förfarna män du själv hade, o Tyrus, dem tog du till skeppare.
Gebals äldste och dess förfarnaste män tjänade dig med att bota dina läckor.
Alla havets skepp med sina sjömän tjänade dig vid ditt varubyte.
Perser, ludéer och putéer funnos i din här och voro ditt krigsfolk.
Sköldar och hjälmar hängde de upp i dig; dessa gåvo dig glans.
Arvads söner stodo med din här runt om på dina murar, gamadéer hade sin plats i dina torn.
Sina stora sköldar hängde de upp runt om på dina murar; de gjorde din skönhet fullkomlig.
Tarsis var din handelsvän, ty du var rik på allt slags gods silver, järn, tenn och bly gavs dig såsom betalning.
Javan, Tubal och Mesek, de drevo köpenskap med dig; trälar och kopparkärl gåvo de dig i utbyte.
Vagnshästar, ridhästar och mulåsnor gåvos åt dig såsom betalning från Togarmas land.
Dedans söner drevo köpenskap med dig ja, många havsländer drevo handel i din tjänst; elfenben och ebenholts tillförde de dig såsom hyllningsgåvor.
Aram var din handelsvän, ty du var rik på konstarbeten; karbunkelstenar, purpurrött tyg, brokiga vävnader och fint linne. koraller och rubiner gåvo de dig såsom betalning.
Juda och Israels land drevo köpenskap med dig; vete från Minnit, bakverk och honung, olja och balsam gåvo de dig i utbyte.
Damaskus var din handelsvän, ty du var rik på konstarbeten, ja, på allt slags gods; de kommo med vin från Helbon och med ull från Sahar.
Vedan och Javan gåvo dig spånad såsom betalning; konstsmitt järn och kassia och kalmus fick du i utbyte.
Dedan drev köpenskap hos dig med sadeltäcken att rida på.
Araberna och Kedars alla furstar, de drevo handel i din tjänst; med lamm och vädurar och bockar drevo de handel hos dig.
Sabas och Raemas köpmän drevo köpenskap med dig; kryddor av allra yppersta slag och alla slags ädla stenar och guld gåvo de dig såsom betalning.
Haran, Kanne och Eden, Sabas köpmän, Assur och Kilmad drevo köpenskap med dig.
De drevo köpenskap hos dig med sköna kläder, med mörkblå, brokigt vävda mantlar, med mångfärgade täcken, med välspunna, starka tåg, på din marknad.
Tarsis-skepp foro åstad med dina bytesvaror.
Så fylldes du med gods och blev tungt lastad, där du låg i havet.
Och dina roddare förde dig åstad, ut på de vida vattnen.
Då kom östanvinden och krossade dig. där du låg i havet.
Ditt gods, dina handels- och bytesvaror, dina sjömän och skeppare, dina läckors botare och dina bytesmäklare, allt krigsfolk på dig, allt manskap som fanns ombord på dig, de sjunka nu ned i havet, på ditt falls dag.
Vid dina skeppares klagorop bäva markerna,
och alla som ro med åror övergiva sina skepp; sjömän och alla skeppare på havet begiva sig i land.
De ropa högt över ditt öde och klaga bittert; de strö stoft på sina huvuden och vältra sig i aska.
De raka sig skalliga för din skull och hölja sig i sorgdräkt; de gråta över dig i bitter sorg, under bitter klagan.
Med jämmer stämma de upp en klagosång om dig, en klagosång över ditt öde: »Vem var såsom Tyrus, hon som nu ligger i det tysta ute i havet?»
Där dina handelsvaror sattes i land från havet mättade du många folk; med ditt myckna gods och dina många bytesvaror riktade du jordens konungar.
Men nu, då du har förlist och försvunnit ifrån havet, ned i vattnens djup, nu hava dina bytesvaror och allt ditt manskap sjunkit med dig.
Havsländernas alla inbyggare häpna över ditt öde, deras konungar stå rysande, med förfäran i sina ansikten.
Köpmännen ute bland folken vissla åt dig; du har tagit en ände med förskräckelse till evig tid.
Och HERRENS ord kom till mig; han sade:
Du människobarn, säg till fursten i Tyrus: Så säger Herren, HERREN: Eftersom ditt hjärta är så högmodigt och du säger: »Jag är en gud, ja, på ett gudasäte tronar jag mitt ute i havet», du som dock är en människa och icke en gud, huru mycket du än i ditt hjärta tycker dig vara en gud --
och sant är att du är visare än Daniel; ingen hemlighet är förborgad för dig;
genom din vishet och ditt förstånd har du skaffat dig rikedom, guld och silver har du skaffat dig i dina förrådshus;
och genom den stora vishet varmed du drev din köpenskap har du ökat din rikedom, och så har ditt hjärta blivit högmodigt för din rikedoms skull --
därför säger Herren, HERREN så: Eftersom du i ditt hjärta tycker dig vara en gud,
se, därför skall jag låta främlingar komma över dig, de grymmaste folk; och de skola draga ut sina svärd mot din visdoms skönhet och skola oskära din glans.
De skola störta dig ned i graven, och du skall dö såsom en dödsslagen man, mitt ute i havet.
Månne du då skall säga till din dråpare: »Jag är en gud», du som ej är en gud, utan en människa, i dens våld, som slår dig till döds?
Såsom de oomskurna dö, så skall du dö, för främlingars hand.
Ty jag har talat, säger Herren, HERREN.
Och HERRENS ord kom till mig han sade:
Du människobarn, stäm upp en klagosång över konungen i Tyrus och säg till honom: Så säger Herren, HERREN: Du var ypperst bland härliga skapelser, full med vishet och fullkomlig i skönhet.
I Eden, Guds lustgård, bodde du, höljd i alla slags ädla stenar: karneol, topas och kalcedon, krysolit, onyx och jaspis, safir, karbunkel och smaragd, jämte guld; du var prydd med smycken och klenoder, beredda den dag då du skapades.
Du var en kerub, som skuggade vida, och jag hade satt dig att vara på det heliga gudaberget, du fick där gå omkring bland gnistrande stenar.
Lyckosam var du på dina vägar från den dag då du skapades, till dess att orättfärdighet blev funnen hos dig.
Men under din myckna köpenskap blev ditt inre fyllt med orätt, och du föll i synd.
Då förvisade jag dig från gudaberget och förgjorde dig, du vittskuggande kerub; du fick ej stanna bland de gnistrande stenarna.
Eftersom ditt hjärta högmodades över din skönhet och du förspillde din vishet för ditt pråls skull, därför slog jag dig ned till jorden och gav dig till pris åt konungarna, så att de fingo se sin lust på dig.
Genom dina många missgärningar vid din orättrådiga köpenskap ohelgade du dina helgedomar.
Därför lät jag eld gå ut ifrån dig, och av den blev du förtärd.
Jag lät dig ligga såsom aska på jorden inför alla som besökte dig.
Alla som kände dig bland folken häpnade över ditt öde.
Du tog en ände med förskräckelse för evig tid.
Och HERRENS ord kom till mig; han sade:
Du människobarn, vänd ditt ansikte mot Sidon och profetera mot det
och säg: Så säger Herren, HERREN: Se, jag skall komma över dig, Sidon, och förhärliga mig i dig.
Ja, att jag är HERREN, det skall man förnimma, när jag håller dom över henne och bevisar mig helig på henne.
Och jag skall sända över henne pest och blod på hennes gator, och dödsslagna män skola falla därinne för ett svärd som skall drabba henne från alla sidor; och man skall förnimma att jag är HERREN.
Sedan skall för Israels hus icke mer finnas någon stingande tagg eller något sårande törne bland alla de grannfolk som nu håna dem; och man skall förnimma att jag är Herren, HERREN.
Ja, så säger Herren, HERREN: När jag församlar Israels barn från de folk bland vilka de äro förströdda, då skall jag bevisa mig helig på dem inför folkens ögon, och de skola sedan få bo i sitt land, det som jag har givit åt min tjänare Jakob.
De skola bo där i trygghet och bygga hus och plantera vingårdar ja, de skola bo i trygghet, när jag håller dom över alla som håna dem på alla sidor; och de skola förnimma att jag är HERREN, deras Gud.
I tionde året, på tolfte dagen i tionde månaden, kom HERRENS ord till mig; han sade:
Du människobarn, vänd ditt ansikte mot Farao, konungen i Egypten, och profetera mot honom och mot hela Egypten.
Tala och säg: Så säger Herren, HERREN: Se, jag skall komma över dig, Farao, du Egyptens konung, du stora drake, som ligger där i dina strömmar och säger: »Min Nilflod är min; själv har jag gjort mig.»
Jag skall sätta krokar i dina käftar och låta fiskarna i dina strömmar fastna vid dina fjäll, och så skall jag draga dig upp ur dina strömmar med alla de fiskar i dina strömmar, som hänga fast vid dina fjäll.
Och jag skall kasta dig ut i öknen med alla fiskarna ifrån dina strömmar; du skall falla på marken och ej tagas bort därifrån eller upphämtas, ty åt markens djur och himmelens fåglar vill jag giva dig till mat;
och alla Egyptens inbyggare skola förnimma att jag är HERREN.
Ty de äro en rörstav för Israels barn;
ja, när dessa fatta i dig med handen, går du sönder och sårar envar av dem i sidan; och när de stödja sig på dig, brytes du av och lämnar dem alla med vacklande länder.
Därför säger Herren, HERREN så: Se, jag vill låta svärd komma över dig, och jag skall utrota ur dig både människor och djur.
Och Egyptens land skall bliva förött och ödelagt, och man skall förnimma att jag är HERREN.
Detta därför att han sade: »Nilfloden är min; själv har jag gjort den.
Ja, därför skall jag komma över dig och dina strömmar, och göra Egyptens land till en ödemark, ett ödelagt land, från Migdol till Sevene, fram till Etiopiens gräns.
Ingen människofot skall gå där fram, och ingen fot av något boskapsdjur skall gå där fram; och det skall ligga obebott i fyrtio år.
Och jag skall göra Egyptens land till en ödemark bland ödelagda länder, och dess städer skola ligga öde bland förhärjade städer i fyrtio år; och jag skall förskingra egyptierna bland folken och förströ dem i länderna.
Ty så säger Herren, HERREN: När fyrtio år äro förlidna, skall jag församla egyptierna från de folk bland vilka de äro förskingrade.
Och jag skall åter upprätta Egypten och låta egyptierna komma tillbaka till Patros' land, varifrån de stamma.
Där skola de bliva ett oansenligt rike,
ja, ett rike oansenligare än andra riken, så att det icke mer skall kunna upphäva sig över folken; jag skall låta dem bliva så få att de icke kunna råda över folken.
Och Israels barn skola icke mer sätta sitt hopp till dem som allenast uppväcka minnet av deras missgärning, när de vända sig till dem; och de skola förnimma att jag är Herren, HERREN.
I tjugusjunde året, på första dagen i första månaden, kom HERRENS ord till mig; han sade:
Du människobarn, Nebukadressar konungen i Babel, har låtit sin här förrätta ett svårt arbete mot Tyrus; alla huvuden hava blivit skalliga och alla skuldror sönderskavda.
Men han och hans här hava icke fått någon lön från Tyrus för det arbete som han har förrättat mot det.
Därför säger Herren, HERREN så: Se, jag vill giva Egyptens land åt Nebukadressar, konungen i Babel; och han skall föra bort dess rikedomar och taga rov därifrån och göra byte där, och detta skall hans här få till lön.
Såsom en vedergällning för hans arbete giver jag honom Egyptens land; ty för min räkning hava de utfört sitt verk, säger Herren, HERREN.
På den tiden skall jag låta ett horn växa upp åt Israels hus, och du skall få upplåta din mun mitt ibland dem; och de skola förnimma att jag är HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn, profetera och säg: Så säger Herren, HERREN: Jämren eder: »Ack ve, vilken dag!»
Ty dagen är nära, HERRENS dag är nära; en molnhöljd dag är det, hednafolkens stund är inne.
Ett svärd kommer över Egypten, och Etiopien fattas av ångest, när de slagna falla i Egypten och dess rikedomar föras bort och dess grundvalar upprivas.
Etiopier, putéer och ludéer, och hela hopen av främmande folk, och kubéer och förbundslandets söner skola med dem falla för svärd.
Så säger HERREN: Ja, Egyptens försvarare skola falla, och dess stolta makt skall störtas ned; från Migdol till Sevene skola de som bo där falla för svärd, säger Herren, HERREN.
Och deras land skall ligga öde bland ödelagda länder, och städerna där skola vara bland förhärjade städer.
Och man skall förnimma att jag är HERREN, när jag tänder eld på Egypten och låter alla dess hjälpare varda krossade.
På den dagen skola sändebud draga ut från mig på skepp, för att injaga skräck hos Etiopien mitt i dess trygghet; och man skall där fattas av ångest på Egyptens dag; ty se, det kommer!
Så säger Herren, HERREN: Ja, jag skall göra slut på Egyptens rikedomar genom Nebukadressar, konungen i Babel.
Han och hans folk med honom, de grymmaste hedningar, skola hämtas dit till att fördärva landet; de skola draga sina svärd mot Egypten och uppfylla landet med slagna.
Och jag skall göra strömmarna till torr mark och sälja landet i onda mäns hand.
Jag skall ödelägga landet med allt vad däri är, genom främmande män.
Jag, HERREN, har talat.
Så säger Herren, HERREN: Jag skall ock förstöra de eländiga avgudarna och göra slut på avgudarna i Nof, och ur Egyptens land skall ingen furste mer uppstå; och jag skall låta fruktan komma över Egyptens land.
Jag skall ödelägga Patros och tända eld på Soan och hålla dom över No.
Och jag skall utgjuta min vrede över Sin, Egyptens värn, och utrota den larmande hopen i No.
Ja, jag skall tända eld på Egypten, Sin skall gripas av ångest, No skall bliva intaget och Nof överfallas på ljusa dagen.
Avens och Pi-Besets unga män skola falla för svärd, och själva skola de vandra bort i fångenskap.
I Tehafnehes bliver dagen mörk, när jag där bryter sönder Egyptens ok och dess stolta makt där får en ände; ja, ett moln skall övertäcka det, och dess döttrar skola vandra bort i fångenskap.
Jag skall hålla dom över Egypten, och man skall förnimma att jag är HERREN.
I elfte året, på sjunde dagen i första månaden, kom HERRENS ord till mig; han sade:
Du människobarn, jag har brutit sönder Faraos, den egyptiske konungens, arm; och se, den har icke blivit förbunden, man har icke brukat läkemedel, icke lindat den, icke lagt på den förband, för att åter göra den stark nog till att föra svärdet.
Därför säger Herren, HERREN så: Se, jag skall komma över Farao, konungen i Egypten, och bryta sönder hans armar, både den som ännu är stark och den som redan är sönderbruten, och skall låta svärdet falla ur hans hand.
Och jag skall förskingra egyptierna bland folken och förströ dem i länderna.
Den babyloniske konungens armar skall jag stärka, och jag skall sätta milt svärd i hans hand; men Faraos armar skall jag bryta sönder, så att han upphäver jämmerrop inför honom, såsom en dödsslagen kämpe gör.
Ja, jag skall stärka den babyloniske konungens armar, men Faraos armar skola sjunka ned; och man skall förnimma att jag är HERREN, när jag sätter mitt svärd i den babyloniske konungens hand, för att han skall svänga det mot Egyptens land.
Och jag skall förskingra egyptierna bland folken och förströ dem i länderna; och de skola förnimma att jag är HERREN.
I elfte året, på första dagen i tredje månaden, kom HERRENS ord till mig; han sade:
Du människobarn, säg till Farao, konungen i Egypten, och till hans larmande hop: Vem kan förliknas med dig i din storhet?
Se, du är ett ädelt träd, en ceder på Libanon, med sköna grenar och skuggrik krona och hög stam, en som med sin topp räcker upp bland molnen.
Vatten gåvo den växt, djupets källor gjorde den hög.
Ty med sina strömmar omflöto de platsen där den var planterad; först sedan sände de sina flöden till alla andra träd på marken.
Så fick den högre stam än alla träd på marken, den fick talrika kvistar och långa grenar, genom det myckna vatten den hade, när den sköt skott.
Alla himmelens fåglar byggde sig nästen bland dess kvistar, under dess grenar födde alla markens djur sina ungar, och i dess skugga bodde allahanda stora folk.
Och den blev skön genom sin storhet och genom sina grenars längd, där den stod med sin rot invid stora vatten.
Ingen ceder i Guds lustgård gick upp emot denna, ingen cypress hade kvistar som kunde förliknas med dennas, ingen lönn bar grenar, jämförliga med dennas; nej, intet träd i Guds lustgård liknade den i skönhet
Så skön hade jag låtit den bliva, i dess rikedom på grenar, att alla Edens träd i Guds lustgård måste avundas den.
Därför säger Herren, HERREN så Eftersom du växte så hög, ja, eftersom ditt träd sträckte sin topp upp bland molnen och förhävde sig i sitt hjärta över att det var så högt,
därför skall jag prisgiva det åt en som är väldig bland folken.
Han skall förvisso utföra sitt verk därpå, ty för dess ogudaktighets skull har jag förkastat det.
Ja, främlingar hava fått hugga ned det, de grymmaste folk, och hava låtit det ligga.
Dess kvistar hava nu fallit på bergen och i alla dalar; dess grenar hava blivit avbrutna och kastade i alla landets bäckar, och alla folk på jorden hava måst draga bort därifrån och försaka dess skugga och låta det ligga.
På dess kullfallna stam bo alla himmelens fåglar, och på dess grenar lägra sig alla markens djur.
Så sker, för att ett träd som växer vid vatten aldrig skall yvas över sin höjd och sträcka sin topp upp bland molnen; ja, för att icke ens de väldigaste av dem skola stå och yvas, intet träd som har haft vatten att dricka.
Ty de äro allasammans hemfallna åt döden och måste ned i jordens djup, till att vara där bland människors barn, hos dem som hava farit ned i graven.
Så säger Herren, HERREN: På den dag då det for ned till dödsriket lät jag djupet för dess skull hölja sig i sorgdräkt; jag hämmade strömmarna där, och de stora vattnen höllos tillbaka.
Jag lät Libanon för dess skull kläda sig i svart, och alla träd på marken förtvinade i sorg över det.
Genom dånet av dess fall kom jag folken att bäva, när jag störtade det ned i dödsriket, till dem som hade farit ned i graven.
Men då tröstade sig i jordens djup alla Edens träd, de yppersta och bästa på Libanon, alla de som hade haft vatten att dricka.
Också de hade, såsom det trädet, måst fara ned till dödsriket, till dem som voro slagna med svärd; dit foro ock de som hade varit dess stöd och hade bott i dess skugga bland folken.
Kan nu något bland Edens träd förliknas med dig i härlighet och storhet?
Och dock skall du, såsom Edens träd, störtas ned i jordens djup och ligga där bland oomskurna, hos dem som äro slagna med svärd.
Så skall det gå Farao och hela hans larmande hop, säger Herren, HERREN.
I tolfte året, på första dagen i tolfte månaden, kom HERRENS ord till mig; han sade:
Du människobarn, stäm upp en klagosång över Farao, konungen i Egypten, och säg till honom: Det är förbi med dig, du lejon bland folken!
Och du var dock lik draken i havet, där du for fram i dina strömmar och rörde upp vattnet med dina fötter och grumlade dess strömmar.
Så säger nu Herren, HERREN: Jag skall breda ut mitt nät över dig genom skaror av många folk, och de skola draga upp dig i mitt garn.
Jag skall kasta dig upp på jorden, jag skall slunga dig bort på marken och låta alla himmelens fåglar slå ned på dig och låta de vilda djuren på hela jorden mätta sig med dig.
Jag skall kasta ditt kött på bergen och fylla dalarna med ditt stora skrov.
Och landet som du har nedsölat skall jag vattna med ditt blod ända upp till bergen, och bäckarna skola bliva fulla av dig.
Och när jag utsläcker dig, skall jag övertäcka himmelen och förmörka dess stjärnor; jag skall övertäcka solen med moln, och månens ljus skall icke lysa mer.
Alla ljus på himmelen skall jag förmörka för din skull och låta mörker komma över ditt land, säger Herren, HERREN.
Och många folks hjärtan skall jag slå med skräck, när jag gör din undergång bekant bland folkslagen, ja, i länder som du icke känner.
Jag skall komma många folk att häpna för din skull, och deras konungar skola för din skull gripas av bävan, när jag i deras åsyn svänger mitt svärd; vart ögonblick skola de frukta, envar för sitt liv, på ditt falls dag.
Ty så säger Herren, HERREN: Den babyloniske konungens svärd skall komma över dig.
Jag skall låta din larmande hop falla för hjältars svärd, grymmast bland hedningar äro de alla.
De skola föröda Egyptens härlighet, och hela dess larmande hop skall förgöras;
jag skall utrota all dess boskap, den som betar vid det myckna vattnet.
Av människofot skall det icke mer röras upp, ej heller röras upp av boskapsklövar.
Sedan skall jag låta deras vatten sjunka undan och deras strömmar flyta bort såsom olja, säger Herren, HERREN,
i det jag gör Egyptens land till en ödslig ödemark och berövar landet allt vad däri är, när jag nu slår alla dess inbyggare, så att man förnimmer att jag är HERREN.
Detta är en klagosång som man skall sjunga, ja, folkens döttrar skola sjunga den; de skola sjunga den över Egypten med hela dess larmande hop, säger Herren, HERREN.
I tolfte året, på femtonde dagen i månaden, kom HERRENS ord till mig; han sade:
Du människobarn, sjung sorgesång över Egyptens larmande hop.
Bjud henne att såsom döttrarna av de väldigaste folk fara ned i jordens djup, till dem som redan hava farit ned i graven.
Finnes någon så ringa att du är förmer än hon?
Nej, far du ned och låt dig bäddas bland de oomskurna.
Bland män som äro slagna med svärd skola ock dina falla.
Svärdet är redo; släpen bort henne med hela hennes larmande hop.
Mäktiga hjältar skola tala till Farao ur dödsriket, till honom och till hans hjälpare: »Ja, de hava måst fara hitned, och nu ligga de där, de oomskurna, slagna med svärd.»
Där ligger redan Assur med hela sin skara; runt omkring honom har denna sin gravplats.
Allasammans ligga de där slagna, fallna för svärd.
Sin grav har han fått längst ned i underjorden, och runt omkring honom ligger hans skara begraven.
Allasammans ligga de slagna, fallna för svärd, de man som en gång utbredde skräck i de levandes land.
Där ligger Elam med hela sin larmande hop, vilande runt omkring hans grav.
Allasammans ligga de slagna, männen som föllo för svärd, och som oomskurna måste fara, ned i jordens djup, desamma som en gång utbredde skräck omkring sig i de levandes land; nu måste de bära sin skam bland de andra som hava farit ned i graven.
Ja, bland slagna har han fått sitt läger med hela sin larmande hop; runt omkring honom har denna sin gravplats.
Allasammans ligga de där oomskurna, slagna med svärd; en gång utbredde sig ju skräck omkring dem i de levandes land, men de måste nu bära sin skam bland dem som hava farit ned i graven.
Ja, bland slagna har han fått sin plats.
Där ligger Mesek-Tubal med hela sin larmande hop; runt omkring honom har denna sin gravplats.
Allasammans ligga de där oomskurna, slagna med svärd; en gång utbredde de ju skräck omkring sig i de levandes land.
Men dessa fallna män ur de oomskurnas hop, de få icke vila bland hjältarna, bland dem som hava farit ned till dödsriket i sin krigiska rustning och fått sina svärd lagda under sina huvuden.
Nej, deras missgärningar hava kommit över deras ben.
De utbredde ju skräck i de levandes land, såsom hjältar göra.
Ja, också du skall bliva krossad bland de oomskurna och få ligga bland dem som äro slagna med svärd.
Där ligger Edom med sina konungar och alla sina hövdingar; huru mäktiga de än voro, hava de nu fått sin plats bland dem som äro slagna med svärd; de måste ligga bland de oomskurna, bland dem som hava farit ned i graven.
Där ligga Nordlandets furstar allasammans, med alla sidonier, ty de hava måst fara ned till de slagna, de hava kommit på skam, trots den skräck de utbredde genom sina väldiga gärningar.
Och de ligga där oomskurna bland dem som hava blivit slagna med svärd; de måste bära sin skam bland dem som hava farit ned i graven.
Dem skall nu Farao få se, och han skall så trösta sig över hela sin larmande hop.
Ja, Farao och hela hans har äro slagna med svärd, säger Herren, HERREN.
Ty väl utbredde jag skräck för honom i de levandes land, men nu måste han, Farao, med hela sin larmande hop, låta sig bäddas bland de oomskurna, hos dem som äro slagna med svärd, säger Herren, HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn, tala till dina landsmän och säg till dem: Om jag vill låta svärdet komma över ett land, och folket i landet har utsett bland sig en man som det har gjort till sin väktare,
och denne ser svärdet komma över landet och stöter i basunen och varnar folket,
men den som får höra basunljudet ända icke låter varna sig, och svärdet sedan kommer och tager honom bort, då kommer hans blod över hans eget huvud.
Ty han hörde ju basunljudet, men lät icke varna sig; därför kommer hans blod över honom själv.
Om han hade låtit varna sig, så hade han räddat sitt liv. --
Men om väktaren ser svärdet komma och icke stöter i basunen och folket så icke bliver varnat, och svärdet sedan kommer och tager bort någon bland dem, då bliver visserligen denne borttagen genom sin egen missgärning, men hans blod skall jag utkräva av väktarens hand.
Dig, du människobarn, har jag satt till en väktare för Israels hus, för att du å mina vägnar skall varna dem, när du hör ett ord från min mun.
Om jag säger till den ogudaktige: »Du ogudaktige, du måste dö», och du då icke säger något till att varna den ogudaktige för hans väg, så skall väl den ogudaktige dö genom sin missgärning, men hans blod skall jag utkräva av din hand.
Men om du varnar den ogudaktige för hans väg, på det att han må vända om ifrån den, och han likväl icke vänder om ifrån sin väg, då skall visserligen han dö genom sin missgärning, men du själv har räddat din själ.
Och du, människobarn, säg till Israels hus: I sägen så: »Våra överträdelser och synder tynga på oss och vi försmäkta genom dem.
Huru kunna vi då bliva vid liv?»
Men svara dem: Så sant jag lever, säger Herren, HERREN, jag har ingen lust till den ogudaktiges död, utan fastmer därtill att den ogudaktige vänder om från sin väg och får leva.
Så vänden då om, ja, vänden om från edra onda vägar; ty icke viljen I väl dö, I av Israels hus?
Men du, människobarn, säg till dina landsmän: Den rättfärdiges rättfärdighet skall icke rädda honom, när han begår överträdelser; och den ogudaktige skall icke komma på fall genom sin ogudaktighet, när han vänder om från sin ogudaktighet, lika litet som den rättfärdige skall kunna leva genom sin rättfärdighet, när han syndar.
Om jag säger till den rättfärdige att han skall få leva, och han sedan i förlitande på sin rättfärdighet gör vad orätt är, så skall intet ihågkommas av all hans rättfärdighet, utan genom det orätta som han gör skall han dö.
Och om jag säger till den ogudaktige: »Du måste dö», och han sedan vänder om från sin synd och övar rätt och rättfärdighet,
så att han, den ogudaktige, give tillbaka den pant han har fått och ersätter vad han har rövat och vandrar efter livets stadgar, så att han icke gör vad orätt är, då skall han förvisso leva och icke dö.
Ingen av de synder han har begått skall då tillräknas honom; han har övat rätt och rättfärdighet, därför skall han förvisso få leva. --
Men nu säga dina landsmän: »Herrens väg är icke alltid densamma», då det fastmer är deras egen väg som icke alltid är densamma.
Om den rättfärdige vänder om från sin rättfärdighet och gör vad orätt är, så måste han just därför dö.
Men om den ogudaktige vänder om från sin ogudaktighet och övar rätt och rättfärdighet, då skall han just därför få leva.
Och ändå sägen I: »Herrens väg är icke alltid densamma.»
Jo, jag skall döma var och en av eder efter hans vägar, I av Israels hus.
I det tolfte året sedan vi hade blivit bortförda i fångenskap, på femte dagen i tionde månaden, kom en flykting ifrån Jerusalem till mig med budskapet: »Staden är intagen.»
Nu hade på aftonen före flyktingens ankomst HERRENS hand kommit över mig; men på morgonen öppnade han åter min mun, just före mannens ankomst, så att jag, då nu min mun blev öppnad, upphörde att vara stum.
Och HERRENS ord kom till mig; han sade:
Du människobarn, de som bo ibland ruinerna där borta i Israels land säga »Abraham var en ensam man, och han fick dock landet till besittning.
Vi äro många, oss måste väl landet då vara givet till besittning!»
Säg därför till dem: Så säger Herren, HERREN: I äten kött med blodet i, I upplyften edra ögon till edra eländiga avgudar, och I utgjuten blod; och likväl skullen I få hava landet till besittning!
I trotsen på edra svärd, I bedriven vad styggeligt är, I skänden varandras hustrur; och likväl skullen I få hava landet till besittning!
Nej; så skall du säga till dem: Så säger Herren, HERREN: Så sant jag lever, de som bo där bland ruinerna skola falla för svärd; och dem som bo på landsbygden skall jag giva till mat åt de vilda djuren, och de som bo i bergfästen eller i grottor skola dö genom pest.
Jag skall göra landet öde och tomt, och dess stolta makt skall få en ände; och Israels berg skola ödeläggas, så att ingen går där fram.
Och de skola förnimma att jag är HERREN, när jag gör landet öde och tomt, för alla de styggelsers skull som de hava bedrivit.
Men du, människobarn, dina landsmän, som orda om dig invid väggarna och i ingångarna till husen, de tala sinsemellan, den ene med den andre, och säga: »Kom, låt oss höra vad det är för ett ord som nu utgår från HERREN.»
Och de komma till dig, såsom gällde det en folkförsamling, och sätta sig hos dig såsom mitt folk; och de höra dina ord, men göra icke efter dem.
Ty väl hopgöra de med munnen ljuvliga ord, men deras hjärtan stå blott efter egen vinning.
Och se, du är för dem, såsom när någon som har vacker röst och spelar väl sjunger en kärleksvisa; de höra väl dina ord, men göra icke efter dem.
Men när det kommer -- ty se det kommer! -- då skola de förnimma att en profet har varit ibland dem.
Och HERRENS ord kom till mig; han sade:
Du människobarn, profetera mot Israels herdar, profetera och säg till dem, till herdarna: Så säger Herren, HERREN: Ve eder, I Israels herdar, som haven sörjt allenast för eder själva!
Var det då icke för hjorden som herdarna borde sörja?
I stället åten I upp det feta, med ullen klädden I eder, det gödda slaktaden I; men om hjorden vårdaden I eder icke.
De svaga stärkten I icke, det sjuka heladen I icke, det sargade förbunden I icke, det fördrivna förden I icke tillbaka, det förlorade uppsökten I icke, utan med förtryck och hårdhet fören I fram mot dem.
Så blevo de förskingrade, därför att de icke hade någon herde, de blevo till mat åt alla markens djur, ja, de blevo förskingrade.
Mina får gå nu vilse på alla berg och alla höga kullar; över hela jorden äro mina får förskingrade, utan att någon frågar efter dem eller uppsöker dem.
Hören därför HERRENS ord, I herdar:
Så sant jag lever, säger Herren, HERREN, sannerligen, eftersom mina får hava lämnats till rov, ja, eftersom mina får hava blivit till mat åt alla markens djur, då de nu icke hava någon herde, och eftersom mina herdar icke fråga efter mina får ja, eftersom herdarna sörja för sig själva och icke sörja för mina får,
därför, I herdar: Hören HERRENS ord:
Så säger Herren, HERREN: Se, jag skall komma över herdarna och utkräva mina får ur deras hand och göra slut på deras herdetjänst; och herdarna skola då icke mer kunna sörja för sig själva, ty jag skall rädda mina får ur deras gap, så att de icke bliva till mat åt dem.
Ty så säger Herren, HERREN: Se, jag skall själv taga mig an mina får och leta dem tillsammans.
Likasom en herde letar tillsammans sin hjord, när hans får äro förströdda omkring honom, så skall ock jag leta tillsammans mina får och rädda dem från alla de orter till vilka de förskingrades på en dag av moln och töcken.
Och jag skall föra dem ut ifrån folken och församla dem ur länderna, och skall låta dem komma till sitt eget land och föra dem i bet på Israels berg, vid bäckarna och var man eljest kan bo i landet.
På goda betesplatser skall jag föra dem i bet, på Israels höga berg skola de få sina betesmarker; där skola de lägra sig på goda betesmarker, och fett bete skola de hava på Israels berg.
Jag skall själv föra mina får i bet och själv utse lägerplatser åt dem, säger Herren, HERREN.
Det förlorade skall jag uppsöka, det fördrivna skall jag föra tillbaka, det sargade skall jag förbinda, och det svaga skall jag stärka.
Men det feta och det starka skall jag förgöra; ja, jag skall sköta det såsom rätt är.
Men I, mina får, så säger Herren, HERREN: Se, jag vill döma mellan får och får, mellan vädurar och bockar.
Är det eder icke nog att I fån beta på den bästa betesplatsen, eftersom I med edra fötter trampen ned vad som är kvar på eder betesplats?
Och är det eder icke nog att I fån dricka det klaraste vattnet, eftersom I med edra fötter grumlen vad som har lämnats kvar?
Skola mina får beta av det som edra fötter hava trampat ned, och dricka vad edra fötter hava grumlat?
Nej; därför säger Herren, HERREN så till dem: Se, jag skall själv döma mellan de feta fåren och de magra fåren.
Eftersom I med sida och bog stöten undan alla de svaga och med edra horn stången dem, till dess att I haven drivit dem ut och förskingrat dem,
därför skall jag frälsa mina får, så att de icke mer bliva till rov, och skall döma mellan får och får.
Och jag skall låta en herde uppstå, gemensam för dem alla, och han skall föra dem i bet, nämligen min tjänare David; ja, han skall föra dem i bet, han skall vara deras herde.
Jag, HERREN, skall vara deras Gud, men min tjänare David skall vara hövding bland dem.
Jag, HERREN, har talat.
Och jag skall med dem sluta ett fridsförbund; jag skall göra ände på vilddjuren i landet, så att man i trygghet kan bo mitt i öknen och sova i skogarna.
Och jag skall låta dem själva och landet runt omkring min höjd bliva till välsignelse.
Jag skall låta regn falla i rätt tid; regnskurar till välsignelse skall det bliva.
Träden på marken skola bära sin frukt, och jorden skall giva sin gröda, och själva skola de bo i sitt land i trygghet; och de skola förnimma att jag är HERREN, när jag bryter sönder deras ok och räddar dem från de människors hand, som hava hållit dem i träldom.
De skola sedan icke mer bliva ett byte för folken, och markens djur skola ej äta upp dem, utan de skola bo i trygghet, och ingen skall förskräcka dem.
Och jag skall åt dem låta en plantering växa upp, som skall bliva dem till berömmelse; och de som bo i landet skola icke mer ryckas bort av hunger, ej heller skola de mer lida smälek av folken.
Och de skola förnimma att jag, HERREN, deras Gud, är med dem, och att de, Israels hus, äro mitt folk, säger Herren, HERREN.
Ja, I ären mina får, I ären får i min hjord, människor som I ären, och jag är eder Gud, säger Herren, HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn, vänd ditt ansikte mot Seirs berg och profetera mot det;
säg till det: Så säger Herren, HERREN: Se, jag skall komma över dig, du Seirs berg, och uträcka min hand mot dig och göra dig öde och tomt.
Jag skall göra dina städer till ruiner, och självt skall du bliva öde; och du skall förnimma att jag är HERREN.
Eftersom du har hyst en evig fiendskap mot Israels barn och givit dem till pris åt svärdet under deras ofärds tid, den tid då missgärningen hade nått sin gräns,
därför, så sant jag lever, säger Herren, HERREN, skall jag förvandla dig till blod, och blod skall förfölja dig; eftersom du icke har hatat blod, skall blod förfölja dig.
Ja, jag skall göra Seirs berg tomt och öde och utrota därifrån envar som färdas där, fram eller tillbaka.
Och jag skall uppfylla dess berg med dess slagna män; ja, på dina höjder, i dina dalar och vid alla dina bäckar skola svärdsslagna män falla.
Jag skall göra dig till en ödemark för evärdlig tid, och dina städer skola icke mer bliva bebodda; och I skolen förnimma att jag är HERREN.
Eftersom du sade: »De båda folken och de båda länderna skola bliva mina, vi skola taga dem i besittning» -- detta fastän HERREN bodde där --
därför, så sant jag lever, säger Herren, HERREN, skall jag utföra mitt verk med samma vrede och nitälskan varmed du i din hätskhet har utfört ditt verk mot dem; och jag skall göra mig känd bland dem, när jag dömer dig.
Och du skall förnimma att jag är HERREN.
Jag har hört alla de smädelser som du har talat mot Israels berg, i det du har sagt: »Det är en ödemark; de äro givna åt oss till mat.»
Ja, I spärraden upp munnen mot mig och togen den full av ord mot mig; jag har väl hört det.
Så säger Herren, HERREN: Till hela jordens glädje skall jag göra dig till en ödemark.
Därför att du gladde dig åt att Israels hus' arvedel blev ödelagd, därför skall jag göra likaså med dig.
Du skall bliva en ödemark, du Seirs berg, du hela Edom, så långt du sträcker dig; och man skall förnimma att jag är HERREN.
Och du, människobarn, profetera om Israels berg och säg: I Israels berg, hören HERRENS ord.
Så säger Herren, HERREN: Eftersom fienden säger om eder: »Rätt så, de urgamla offerhöjderna hava nu blivit vår besittning»,
därför må du profetera och säga: Så säger Herren, HERREN: Eftersom, ja, eftersom man har förött eder och fikar efter eder från alla sidor, för att I måtten tillfalla de övriga folken såsom deras besittning och eftersom I ären så utsatta för onda tungors hån och folks förtal,
därför, I Israels berg, mån I nu höra Herrens, HERRENS ord: Så säger Herren, HERREN till bergen och höjderna, till bäckarna och dalarna, till de förödda ruinerna och de övergivna städerna, som hava lämnats till rov och spott åt de övriga folken runt omkring,
ja, därför säger Herren, HERREN så: Sannerligen, i brinnande nitälskan talar jag mot de övriga folken och mot Edom, så långt det sträcker sig, ja, mot dessa som med hela sitt hjärtas glädje och i sitt sinnes övermod hava tillägnat sig mitt land såsom besittning, för att driva ut dess inbyggare och göra det till sitt byte.
Profetera alltså om Israels land och säg till bergen och höjderna, till bäckarna och dalarna: Så säger Herren, HERREN: Se, i nitälskan och vrede är det som jag talar, eftersom I liden sådan smälek av folken.
Därför säger Herren, HERREN så Jag upplyfter min hand och betygar: Sannerligen, folken runt omkring eder skola själva få lida smälek.
Men I, Israels berg, I skolen åter grönska och bära frukt åt mitt folk Israel, ty snart skola de komma åter.
Ty se, jag skall komma till eder, jag skall vända mig till eder, och I skolen bliva brukade och besådda.
Och jag skall församla på eder människor i myckenhet, alla Israels barn, så många de äro; och städerna skola ånyo bliva bebodda och ruinerna åter byggas upp.
Ja, jag skall församla på eder människor och boskap i myckenhet, och de skola föröka sig och bliva fruktsamma.
Jag skall låta eder bliva bebodda, alldeles såsom I fordom voren; ja, jag skall göra eder ännu mer gott, än I förut fingen röna; och I skolen förnimma att jag är HERREN.
Jag skall låta människor åter vandra fram över eder, nämligen mitt folk Israel; de skola hava dig till besittning, och du skall vara deras arvedel; och du skall icke vidare döda deras barn.
Så säger Herren, HERREN: Eftersom man säger till dig: »Du är en människoäterska, du har dödat ditt eget folks barn»,
därför skall du nu icke mer få äta upp människor och icke mer få döda ditt folks barn, säger Herren, HERREN.
Jag skall icke mer låta dig höra smälek av folken, och du skall icke mer nödgas bära folkslagens förakt; ej heller skall du mer bringa ditt folk på fall, säger Herren, HERREN.
Och HERRENS ord kom till mig; han sade:
Du människobarn när Israels barn ännu bodde i sitt land, då orenade de det genom sitt väsende och sina gärningar; såsom en kvinnas orenhet var deras väsende för mig.
Då utgöt jag min vrede över dem, för det blods skull som de hade utgjutit över landet, och därför att de hade orenat det med sina eländiga avgudar.
Jag förskingrade dem bland folken, och de blevo förströdda i länderna; efter deras väsende och deras gärningar dömde jag dem.
Men till vilka folk de än kommo vanärade de mitt heliga namn, i det att man sade om dem: »Detta är HERRENS folk, och de hava likväl måst draga ut ur sitt land.
Då ville jag skona mitt heliga namn, som Israels barn vanärade bland de folk till vilka de kommo.
Säg därför till Israels barn: Så säger Herren, HERREN: Icke för eder skull gör jag detta, I Israels barn, utan för mitt heliga namns skull, som I haven vanärat bland de folk till vilka I haven kommit.
Jag vill nu helga mitt stora namn, som har blivit vanärat bland folken, i det att I haven vanärat det bland dem; och folken skola förnimma att jag är HERREN, säger Herren, HERREN, när jag bevisar mig helig på eder inför deras ögon.
Ty jag skall hämta eder ifrån folken och församla eder ifrån alla länder och föra eder till edert land.
Och jag skall stänka rent vatten på eder, så att I bliven rena; jag skall rena eder från all eder orenhet och från alla edra eländiga avgudar.
Och jag skall giva eder ett nytt hjärta och låta en ny ande komma i edert bröst; jag skall taga bort stenhjärtat ur eder kropp och giva eder ett hjärta av kött.
Jag skall låta min Ande komma i edert bröst och så göra, att I vandren efter mina stadgar och hållen mina rätter och gören efter dem.
Så skolen I få bo i det land som jag gav åt edra fäder, och I skolen vara mitt folk, och jag skall vara eder Gud.
Och jag skall frälsa eder från all eder orenhet.
Och jag skall kalla fram säden och låta den bliva ymnig och skall icke mer låta någon hungersnöd komma över eder.
Ja, ymnig skall jag låta trädens frukt och markens gröda bliva, för att I icke mer skolen lida hungersnödens smälek bland folken.
Då skolen I tänka på edra onda vägar och på edra gärningar, som icke voro goda; och I skolen känna leda vid eder själva för edra missgärningars och styggelsers skull.
Men icke för eder skull gör jag detta, säger Herren, HERREN; det vare eder kunnigt.
I mån skämmas och blygas för edra vägar, I Israels barn.
Så säger Herren, HERREN: När jag har renat eder från alla edra missgärningar, då skall jag låta städerna ånyo bliva bebodda, och då skola ruinerna åter byggas upp,
och det förödda landet skall åter bliva brukat, i stället för att det har legat såsom en ödemark inför var man som har gått där fram.
Och då skall man säga: »Det landet som var så förött har nu blivit såsom Edens lustgård, och städerna som voro så ödelagda, förödda och förstörda, de äro nu bebodda och befästa.»
Då skola de folk som äro kvar runt omkring eder förnimma att jag, HERREN, nu åter har byggt upp det som var förstört och ånyo planterat det som var förött.
Jag, HERREN, har talat det, och jag fullbordar det också.
Så säger Herren, HERREN; Också på detta sätt vill jag bönhöra Israels barn, så vill jag handla med dem: jag skall där föröka människorna, så att de bliva såsom fårhjordar.
Såsom hjordar av offerdjur, såsom fårhjordar i Jerusalem vid dess högtider, så skola de hjordar av människor vara, som skola uppfylla de ödelagda städerna.
Och man skall förnimma att jag är HERREN.
HERRENS hand kom över mig, och genom HERRENS Ande fördes jag åstad och sattes ned mitt på slätten, som nu låg full med ben.
Och han förde mig fram runt omkring dem, och jag såg att de lågo där i stor myckenhet utöver dalen och jag såg att de voro alldeles förtorkade.
Och han sade till mig: »Du människobarn, kunna väl dessa ben åter bliva levande?»
Jag svarade: »Herre, HERRE, du vet det.»
Då sade han till mig: »Profetera över dessa ben och säg till dem: I förtorkade ben, hören HERRENS ord;
Så säger Herren, HERREN till dessa ben: Se, jag skall låta ande komma in i eder, så att I åter bliven levande.
Jag skall fästa senor vid eder och låta kött växa på eder och övertäcka eder med hud och giva eder ande, så att I åter bliven levande; och I skolen förnimma att jag är HERREN.»
Och jag profeterade, såsom det hade blivit mig bjudet.
Och när jag nu profeterade, hördes ett rassel, och där blev ett gny, och benen kommo åter tillhopa, så att det ena benet fogades till det andra.
Och jag såg huru senor och kött växte på dem, och huru de övertäcktes med hud därovanpå; men ingen ande var ännu i dem.
Då sade han till mig: »Profetera och tala till anden, ja, profetera, du människobarn, och säg till anden: Så säger Herren, HERREN: Kom, du ande, från de fyra väderstrecken och blås på dessa dräpta, så att de åter bliva levande.»
Och jag profeterade, såsom han hade bjudit mig.
Då kom anden in i dem, och de blevo åter levande och reste sig upp på sina fötter, en övermåttan stor skara.
Och han sade till mig: »Du människobarn, dessa ben, de äro alla Israels barn.
Se, de säga: 'Våra ben äro förtorkade, vårt hopp har blivit om intet, det är ute med oss.'
Profetera därför och säg till dem: Så säger Herren, HERREN: Se, jag vill öppna edra gravar och hämta eder, mitt folk, upp ur edra gravar och låta eder komma till Israels land.
Och I skolen förnimma att jag är HERREN, när jag öppnar edra gravar och hämtar eder, mitt folk, upp ur edra gravar.
Och jag skall låta min ande komma in i eder, så att I åter bliven levande, och jag skall låta eder få bo i edert land; och I skolen förnimma att jag, HERREN, har tala det, och att jag också har fullborda det, säger HERREN.»
Och HERRENS ord kom till mig han sade:
Du människobarn, tag dig en trästav och skriv på den: »För Juda och hans fränder bland Israels barn.»
Tag sedan en annan trästav och skriv på den: »En stav för Josef, Efraim, och för hans fränder av hela Israels hus.»
Foga dem sedan tillhopa med varandra till en enda stav, så att de bliva förenade till ett i din hand.
När då dina landsmän säga till dig: »Förklara för oss vad du menar härmed»,
så svara dem: »Så säger Herren, HERREN: Se, jag vill taga Josefs stav, den som är i Efraims hand, vilken stav ock gäller för de stammar av Israel, som äro hans fränder, och intill denna vill jag lägga Judas stav, båda tillhopa, och så göra dem till en enda stav, så att de bliva ett i min hand.»
Och stavarna som du har skrivit på skall du hålla i din hand inför deras ögon.
Och du skall tala till dem: Så säger Herren, HERREN: Se, jag skall hämta Israels barn ut ifrån de folk till vilka de hava måst vandra bort; jag skall samla dem tillhopa från alla håll och föra dem in i deras land.
Och jag skall göra dem till ett enda folk i landet, på Israels berg; en och samma konung skola de alla hava; de skola icke mer vara två folk och icke mer vara delade i två riken.
Sedan skola de icke mer orena sig med sina eländiga avgudar och styggelser och med alla slags överträdelser.
Och jag skall frälsa dem och hämta dem från alla orter där de hava syndat, och skall rena dem, så att de bliva mitt folk, och jag skall vara deras Gud.
Och min tjänare David skall vara konung över dem, och de skola så alla hava en och samma herde; och de skola vandra efter mina rätter och hålla mina stadgar och göra efter dem.
Så skola de få bo i det land som jag gav åt min tjänare Jakob, det vari edra fäder bodde.
De skola själva få bo där, så ock deras barn och deras barnbarn till evig tid; och min tjänare David skall vara deras hövding evinnerligen.
Och jag skall med dem sluta ett fridsförbund; ett evigt förbund med dem skall det vara.
Jag skall insätta dem och föröka dem och låta min helgedom stå bland dem evinnerligen.
Ja, min boning skall vara hos dem, och jag skall vara deras Gud, och de skola vara mitt folk.
Så skola folken förnimma att jag är HERREN, som helgar Israel, då nu min helgedom förbliver ibland dem evinnerligen.
Och HERRENS ord kom till mig; han sade:
Du människobarn, vänd ditt ansikte mot Gog i Magogs land, mot hövdingen över Ros, Mesek och Tubal, och profetera mot honom
och säg: Så säger Herren, HERREN: Se, jag skall komma över dig, Gog, du hövding över Ros, Mesek och Tubal.
Jag skall locka dig åstad, jag skall sätta krokar i dina käftar och föra dig ut med hela din här, hästar och ryttare, allasammans i präktig rustning, en stor skara, väpnad med skärmar och sköldar, och allasammans med svärd i hand.
Perser, etiopier och putéer är, med dem, allasammans med sköld och hjälm,
Gomer och alla dess härskaror, Togarmas folk ifrån den yttersta norden och alla dess härskaror; ja, många folk har du med dig.
Rusta dig och gör dig redo med alla de skaror som hava församlat sig till dig; och bliv du deras hövitsman.
När lång tid har gått, skall du bliva uppbådad; i kommande år skall du få tåga in i ett land som då har fått ro efter svärdet, och vart folk då har blivit hopsamlat från många andra folk, ja, upp till Israels berg, som så länge lågo öde, men vilkas folk då har blivit hämtat fram ifrån de andra folken, så att alla nu bo där i trygghet.
Dit skall du draga upp, du skall komma såsom ett oväder och vara såsom ett moln som övertäcker landet, du med alla dina härskaror och med många folk som följa dig.
Så säger Herren, HERREN: På den tiden skola planer uppstå i ditt hjärta, och du skall tänka ut onda anslag.
Du skall säga: »Jag vill draga upp mot det obefästa landet, jag vill komma över dessa säkra, som bo där i trygghet, ja, som allasammans bo där utan murar och varken hava bommar eller portar.»
Ty du vill taga rov och göra byte och vända din hand mot ödemarker som nu åter äro bebyggda, och mot ett folk som har blivit hopsamlat från hedningarna, och som nu förvärvar sig boskap och gods, där det bor på jordens mittelhöjd.
Saba och Dedan och Tarsis' köpmän och alla dess unga lejon skola då utfråga dig: »Har du kommit för att taga rov, har du församlat dina skaror till att göra byte till att föra bort silver och guld, till att taga boskap och gods, ja, till att taga stort rov?»
Profetera därför, du människobarn och säg till Gog: Så säger Herren HERREN: Se, på den tiden, när mitt folk Israel åter bor i trygghet, då skall du förnimma det.
Du skall då komma från ditt land längst uppe i norr, du själv och många folk med dig, allasammans ridande på hästar, en stor skara, en talrik här.
Du skall draga upp mot mitt folk Israel och komma såsom ett moln för att övertäcka landet.
I kommande dagar skall detta ske; jag skall då låta dig komma över mitt land, för att folken skola lära känna mig, när jag inför deras ögon bevisar mig helig på dig, du Gog.
Så säger Herren, HERREN: Du är ju den om vilken jag i forna tider talade genom mina tjänare, Israels profeter, som i de tiderna, år efter år, profeterade om att jag skulle låta dig komma över dem.
Men på den dagen, den dag då Gog kommer över Israels land, säger Herren, HERREN, då skall jag giva luft åt min vrede.
Ja, i min nitälskan och min vredes eld betygar jag det: på den dagen skall det förvisso bliva en stor jordbävning i Israels land.
Då skola de bäva för mig, både fiskarna i havet och fåglarna under himmelen och djuren på marken och alla kräldjur som röra sig på jorden och alla människor på jordens yta.
Och bergen skola slås ned och klipporna störta omkull och alla murar falla till jorden.
Och jag skall båda upp svärd mot honom på alla mina berg, säger Herren, HERREN; den enes svärd skall vara vänt mot den andres.
Och jag skall gå till rätta med honom medelst pest och blod; och slagregn och hagelstenar, eld och svavel skall jag låta regna över honom och hans härskaror och över de många folk som följa honom.
Så skall jag bevisa mig stor och helig och göra mig känd inför många folks ögon; och de skola förnimma att jag är HERREN.
Och du, människobarn, profetera mot Gog och säg: Så säger Herren, HERREN: Se, jag skall komma över dig, Gog, du hövding över Ros, Mesek och Tubal.
Jag skall locka dig åstad och leda dig fram och föra dig från landet längst uppe i norr och låta dig komma till Israels berg.
Där skall jag slå bågen ur din vänstra hand och låta pilarna falla ur din högra hand.
På Israels berg skall du falla, med alla dina härskaror och med de folk som följa dig; jag skall giva dig till mat åt rovfåglar av alla slag och åt markens djur.
Ute på marken skall du falla.
Ty jag har talat, säger Herren, HERREN.
Och jag skall sända eld över Magog och över dem som bo trygga i havsländerna; och de skola förnimma att jag är HERREN.
Och jag skall göra mitt heliga namn kunnigt bland mitt folk Israel, jag skall icke mer låta mitt heliga namn bliva ohelgat; och folken skola förnimma att jag är HERREN, helig i Israel.
Se, det kommer, ja, det fullbordas! säger Herren, HERREN.
Detta är den dag om vilken jag har talat.
Sedan skola invånarna i Israels städer gå ditut och taga rustningar, sköldar och skärmar, bågar och pilar, handpåkar och spjut såsom bränsle till att elda med, och de skola elda därmed i sju år.
De skola icke behöva hämta trä från marken eller hugga ved i skogarna, ty de skola elda med rustningarna.
Så skola de taga rov av sina rövare och plundra sina plundrare, säger Herren, HERREN.
På den tiden skall jag där i Israel giva åt Gog en plats till grav, nämligen »De framtågandes dal» öster om havet, och den skall stänga vägen för andra som vilja tåga där fram.
Där skall man begrava Gog och hela hans larmande hop, och man skall kalla den »Gogs larmande hops dal».
Och i sju månader skola Israels barn hålla på med att begrava dem, för att rena landet.
Allt folket i landet skall hålla på med begravandet, och detta skall lända dem till berömmelse.
Så skall ske på den tid då jag förhärligar mig, säger Herren, HERREN.
Och man skall avskilja män som beständigt skola genomvandra landet och begrava dem som tågade där fram, och som ännu ligga kvar ovan jord, och de skola så rena landet; efter sju månaders förlopp skola dessa begynna sitt letande.
När så någon av dessa män, som genomvandra landet, på sin färd får se människoben, då skall han sätta upp en vård därbredvid, till dess att dödgrävarna hinna begrava dem i »Gogs larmande hops dal».
Där skall ock finnas en stad med namnet Hamona.
På detta sätt skola de rena landet.
Du människobarn, så säger Herren, HERREN: Säg till alla slags fåglar och till alla markens djur: Församlen eder och kommen hit; samlen eder tillhopa från alla håll till mitt slaktoffer, till ett stort slaktoffer som jag vill anställa åt eder på Israels berg; I skolen få äta kött och dricka blod.
I skolen få äta kött av hjältar och dricka blod av jordens hövdingar: av vädurar och lamm och bockar och tjurar, allasammans gödda i Basan.
I skolen få äta eder mätta av fett och dricka eder druckna av blod från det slaktoffer som jag anställer åt eder.
Ja, mätten eder vid mitt bord av ridhästar och vagnshästar, av hjältar och allt slags krigsfolk, säger Herren, HERREN.
Och jag skall uppenbara min härlighet bland folken, så att alla folk skola se den dom som jag har utfört, och se huru jag har låtit min hand drabba dem.
Och Israels barn skola förnimma att jag, HERREN, är deras Gud, från den dagen och allt framgent.
Och folken skola förnimma att Israels barn blevo bortförda i fångenskap för sin missgärnings skull, eftersom de voro trolösa mot mig, så att jag måste fördölja mitt ansikte för dem; och jag gav dem då i deras ovänners hand, så att de allasammans föllo för svärd.
Efter deras orenhet och deras överträdelser handlade jag med dem och fördolde mitt ansikte för dem.
Därför säger Herren, HERREN så: Nu skall jag åter upprätta Jakob och förbarma mig över hela Israels hus och nitälska för mitt heliga namn.
Och de skola förgäta sin skam och all den otrohet som de hava begått mot mig, då de nu få bo i trygghet i sitt land, utan att någon förskräcker dem.
Ja, när jag låter dem vända tillbaka ifrån folkslagen och församlar dem från deras fienders länder, då skall jag bevisa mig helig på dem inför många folks ögon.
Och de skola förnimma att jag är HERREN, deras Gud, ty om jag än drev dem bort i fångenskap bland folken, så samlade jag dem sedan tillhopa till deras land och lät ingen enda av dem bliva kvar därute;
och jag skall därefter icke mer fördölja mitt ansikte för dem, ty jag skall utgjuta min Ande över Israels hus, säger Herren, HERREN'.
I det tjugufemte året sedan vi hade blivit bortförda i fångenskap, vid årets begynnelse, på tionde dagen i månaden, i det fjortonde året sedan staden hade blivit intagen, på just den dagen kom HERRENS hand över mig, och han förde mig ditbort.
I en syn från Gud förde han mig till Israels land och satte mig ned på ett mycket högt berg, och på detta var likasom en stad byggd söderut.
Och dit förde han mig, och se, där stod en man vilkens utseende var såsom koppar; han hade ett linnesnöre i sin hand, så ock en mätstång; och han stod vid porten.
Och mannen talade till mig: »Du människobarn, se med dina ögon och hör med dina öron, och akta på allt som jag kommer att visa dig, ty du har blivit förd hit, för att jag skall visa dig det; förkunna för Israels hus allt vad du får se.»
Och jag såg att en mur gick utomkring huset, runt omkring det.
Och mätstången som mannen hade i sin hand var sex alnar lång, var aln en handsbredd längre än en vanlig aln.
Och han mätte murbyggnadens bredd: den var en stång, och dess höjd: den var en stång.
Därefter gick han till en port som låg mot öster och steg uppför dess trappsteg; och han mätte portens ena tröskel: den var en stång bred och sedan den andra tröskeln: den var en stång bred.
Och var vaktkammare var en stång lång och en stång bred, och avståndet mellan vaktkamrarna var fem alnar; och porttröskeln invid portens förhus på inre sidan mätte en stång.
Och han mätte upp portens förhus på inre sidan: det mätte en stång.
Han mätte upp portens förhus det höll åtta alnar, och dess murpelare: de höllo två alnar.
Och portens förhus låg på inre sidan.
Och vaktkamrarna i porten mot öster voro tre på var sida, alla tre lika stora; och murpelarna på båda sidorna voro lika stora.
Och han mätte portöppningens bredd: den var tio alnar, och portens längd: den var tretton alnar.
Och framför vaktkamrarna var en avskrankning, som höll en aln; en aln höll ock avskrankningen på motsatta sidan; och var vaktkammare, på vardera sidan, höll sex alnar.
Och han mätte porten från den ena vaktkammarens tak till den andras: den var tjugufem alnar bred; och dörr låg mot dörr.
Och han tog upp murpelarna till sextio alnar; och intill förgårdens murpelare sträckte sig porten runt omkring.
Och avståndet mellan ingångsportens framsida och förhusets framsida vid den inre portöppningen var femtio alnar.
Och slutna fönster funnos till vaktkamrarna och till deras murpelare invändigt i porten runt omkring, och likaledes i förhusen; fönstren sutto runt omkring invändigt, och murpelarna voro prydda med palmer.
Och han förde mig till den yttre förgården, och jag såg att där voro tempelkamrar och ett stengolv, anlagt runt omkring förgården; trettio tempelkamrar voro uppbyggda på stengolvet.
Och stengolvet gick utefter portarnas sidoväggar, så att det motsvarade portarnas längd; detta var det nedre stengolvet.
Och han mätte avståndet från den nedre portens framsida till den inre förgårdens yttre framsida: det var hundra alnar, både på östra sidan och på norra.
Sedan mätte han ock längden och bredden på den port som låg mot norr på den yttre förgården.
Också den hade tre vaktkamrar på var sida och likaledes murpelare och förhus, lika stora som den förra portens; den var femtio alnar lång och tjugufem alnar bred.
Och fönstren, förhuset och palmerna däri voro lika stora som i den port som låg mot öster; och man steg upp till den på sju trappsteg, och dess förhus låg framför dessa.
Och en port till den inre förgården fanns mitt emot denna port, det var i norr såsom i öster; och han mätte avståndet från den ena porten till den andra: det var hundra alnar.
Därefter lät han mig gå till södra sidan, och jag såg att också på södra sidan fanns en port.
Och han mätte dess murpelare och förhus; de voro lika stora som de andra.
Och fönster funnos på den och på dess förhus runt omkring, likadana som de andra fönstren.
Den var femtio alnar lång och tjugufem alnar bred.
Och trappan ditupp utgjordes av sju trappsteg, och dess förhus låg framför dessa; och den var prydd med palmer på sina murpelare, på båda sidor.
Och en port till den inre förgården fanns ock på södra sidan; och han mätte avståndet från den ena porten till den andra på södra sidan: det var hundra alnar.
Därefter förde han mig till den inre förgården genom södra porten.
Och han mätte den södra porten den var lika stor som de andra
Och dess vaktkamrar, murpelare och förhus voro lika stora som de andra, och fönster funnos på den och på dess förhus runt omkring.
Den var femtio alnar lång och tjugu fem alnar bred.
Och förhus funnos runt omkring tjugufem alnar långa och fem alnar breda.
Och dess förhus låg utåt den yttre förgården, och dess murpelare voro prydda med palmer; och uppgången därtill utgjordes av åtta trappsteg.
Sedan förde han mig till den inre förgårdens östra sida och mätte porten där; den var lika stor som de andra.
Och dess vaktkamrar, murpelare och förhus voro lika stora som de andra, och fönster funnos på den och på dess förhus runt omkring.
Den var femtio alnar lång och tjugufem alnar bred.
Och dess förhus låg mot den yttre förgården, och dess murpelare voro prydda med palmer på båda sidor; och uppgången därtill utgjordes av åtta trappsteg.
Därefter förde han mig till den norra porten och mätte den; den var lika stor som de andra.
Så ock dess vaktkamrar, murpelare och förhus, och fönster funnos på den runt omkring.
Den var femtio alnar lång och tjugufem alnar bred.
Och dess murpelare stodo vid den yttre förgården, och dess murpelare voro prydda med palmer på båda sidor; och uppgången därtill utgjordes av åtta trappsteg.
Och en tempelkammare med sin ingång fanns vid murpelarna, i portarna; där skulle man skölja brännoffren.
Och i portens förhus stodo två bord på var sida, och på dem skulle man slakta brännoffers-, syndoffers- och skuldoffersdjuren.
Och vid den yttre sidovägg som låg norrut, när man steg upp till portens ingång, stodo två bord; och vid den andra sidoväggen på porten förhus stodo ock två bord.
Alltså stodo vid portens sidoväggar fyra bord på var sida, eller tillsammans åtta bord, på vilka man skulle slakta.
Och för brännoffret stodo där fyra bord av huggna stenar, en och en halv aln långa, en och en halv aln breda och en aln höga; på dessa skulle man lägga de redskap som man slaktade brännoffers- och slaktoffersdjuren med.
Och dubbelkrokar, en handsbredd långa, voro fästa innantill runt om kring; och på borden skulle offerköttet läggas.
Och utanför den inre porten funnos för sångarna, på den inre gården, tempelkamrar, som lågo vid den norra portens sidovägg, med sin framsida åt söder; och en annan låg vid den östra portens sidovägg med sin framsida åt norr.
Och han talade till mig: »Denna tempelkammare, vars framsida ligger mot söder, är för de präster som förrätta tjänsten inne i huset.
Och den tempelkammare vars framsida ligger mot norr är för de präster som förrätta tjänsten vid altaret, alltså för Sadoks söner, vilka äro de av Levi barn, som få träda fram till HERREN för att göra tjänst inför honom.»
Och han mätte förgården; den var hundra alnar lång och hundra alnar bred, en liksidig fyrkant; och altaret stod framför huset.
Sedan förde han mig till huset förhus.
Och han mätte för husets murpelare: de höllo fem alnar var på sin sida, så ock porten bredd: den var på var sida tre alnar.
Förhuset var tjugu alnar lång och elva alnar brett, nämligen vid trappstegen på vilka man steg ditupp.
Och vid murpelarna stodo pelare, en på var sida.
Därefter förde han mig till tempelsalen.
Och han mätte murpelarna de voro sex alnar breda, var på sin sida -- tabernaklets bredd.
Och ingången var tio alnar bred, och sidoväggarna vid ingången voro på var sida fem alnar.
Sedan mätte han salens längd: den var fyrtio alnar, och dess bredd: den var tjugu alnar.
Därefter gick han in i det innersta rummet.
Och han mätte murpelarna vid ingången: de höllo två alnar, och ingången: den höll sex alnar, och ingångens bredd: den var sju alnar.
Och han mätte dess längd: den var tjugu alnar, och dess bredd: den var tjugu alnar, framför tempelsalen.
Och han sade till mig: »Detta är det allraheligaste.»
Därefter mätte han husets mur: den höll sex alnar, och sidokamrarnas bredd: den var fyra alnar, runt omkring hela huset.
Och sidokamrarna lågo den ena ovanför den andra, i trettiotre omgångar; och på den mur som sträckte sig innanför sidokamrarna runt omkring funnos avsatser, på vilka de skulle hava sitt fäste; ty i själva husväggen skulle de icke vara infästa.
Härigenom blevo sidokamrarna, där de lågo kring huset, bredare alltefter som de lågo högre upp.
Ty husets kringbyggnad sträckte sig med övervåning ovanpå övervåning runt omkring huset.
Därför växte bredden inåt, alltefter som våningen låg högre upp.
Och från den nedersta våningen steg man så upp i den översta genom den mellersta.
Och jag såg att huset låg på en upphöjd fot, som sträckte sig runt däromkring; sidokamrarnas grundvalar voro nämligen en hel stång höga, sex alnar till kanten.
Sidokamrarnas yttermur var fem alnar tjock; och den plats som blev fri tillhörde husets sidokamrar.
Och mellanrummet bort till tempelkamrarna var tjugu alnar brett runt omkring hela huset.
Och ingångarna till sidokamrarna lågo utåt den fria platsen, en ingång mot norr och en ingång åt söder; den fria platsen var fem alnar bred, runt omkring.
Och den byggnad som låg invid den avsöndrade platsen på västra sidan var sjuttio alnar bred, och byggnadens mur var fem alnar tjock runt omkring och nittio alnar lång.
Och han mätte huset: det var hundra alnar långt.
Och den avsöndrade platsen jämte byggnaden med dess murar utgjorde en längd av hundra alnar.
Och bredden på husets framsida jämte den avsöndrade platsen åt öster utgjorde en längd av hundra alnar.
Och han mätte längden på den byggnad som låg invid den avsöndrade platsen, på dennas baksida, och mätte avsatserna på dess framvägg åt båda sidor -- de höllo hundra alnar -- vidare det inre tempelrummet och förgårdsförhusen,
trösklarna och de slutna fönstren, avsatserna på framväggen runt omkring, i deras tre våningar, platsen invid tröskeln -- som var av polerat trä -- runt omkring,
så ock avståndet från marken upp till fönstren.
Och fönstren voro täckta.
Men ovanför dörren, både in emot det inre rummet och utåt, och eljest utefter hela väggen runt omkring, innantill och utantill, funnos avmätta fält,
på vilka framställdes keruber och palmer, var palm mellan två keruber.
Och var kerub hade två ansikten:
ett människoansikte åt palmen på ena sidan, och ett lejonansikte åt palmen på andra sidan; så var gjort på hela huset runt omkring.
Från marken ända upp över ingången funnos keruber och palmer framställda, så ock på tempelsalens väggar.
Tempelsalens dörröppning var fyrkantig, och framsidan av det heligaste hade sitt givna utseende.
Altaret var av trä, tre alnar högt och två alnar långt, och det hade hörn; och dess långsidor och väggar voro av trä.
Och han talade till mig: »Detta är det bord som skall stå inför HERRENS ansikte.»
Och både tempelsalen och det heligaste hade dubbeldörrar.
Och var dörr hade två dörrskivor, två vridbara dörrskivor: den ena dörren hade två dörrskivor, och likaledes den andra två.
Och på dem, på dörrarna till tempelsalen, funnos framställda keruber och palmer, likasom på väggarna; och på förhusets framsida, utantill, var ett trapphus av trä.
Och slutna fönster och palmer funnos på förhusets sidoväggar, på båda sidor, så ock i husets sidokamrar och i trapphusen.
Och han lät mig gå ut på den yttre förgården den väg som gick åt norr, och förde mig därefter till den byggnad med tempelkamrar, som låg invid den avsöndrade platsen och tillika invid murbyggnaden norrut,
till långsidan, som mätte hundra alnar, med sin ingång i norr; men bredden var femtio alnar.
Ut emot den tjugu alnar breda platsen på den inre förgården och ut emot stengolvet på den yttre förgården lågo avsatserna på det ena husets framvägg mitt emot avsatserna på det andra husets framvägg, i tre våningar.
Och framför tempelkamrarna gick en tio alnar bred gång till den inre förgården, en alnsbred väg; och ingångarna lågo mot norr.
Men de översta tempelkamrarna voro mindre än de andra, ty avsatserna på framväggen togo bort mer rum från dem än från de nedersta och mellersta kamrarna i byggnaden.
Ty kamrarna lågo i tre våningar och hade inga pelare, såsom förgårdarna hade; därför blevo de översta våningens kamrar mer indragna än den nedersta och den mellersta våningens.
Och en yttre skiljemur gick utmed tempelkamrarna åt den yttre förgården till, framför tempelkamrarna, och den var femtio alnar lång.
Ty längden på tempelkammarbyggnaden utåt den yttre förgården var femtio alnar, men åt templet till hundra alnar.
Och nedanför dessa tempelkamrar var ingången från öster, när man ville komma till dem från den yttre förgården.
Där förgårdens skiljemur var som tjockast, lågo ock på östra sidan tempelkamrar invid den avsöndrade platsen och tillika invid murbyggnaden.
Och en väg gick framför dem, likadan som vägen framför tempelkamrarna på norra sidan; och de hade samma längd och bredd.
Och alla utgångar här voro såsom där, både i fråga om övriga anordningar och i fråga om själva dörröppningarna.
Och såsom det var med dörröppningarna på tempelkamrarna vid södra sidan, så fanns också har en dörröppning, vid vilken en väg begynte, en väg som gick utefter den behöriga skiljemuren, och som låg österut, när man gick in i tempelkamrarna.
Och han sade till mig: »De norra och södra tempelkamrarna invid den avsöndrade platsen skola vara de heliga tempelkamrar i vilka prästerna, som få träda fram inför HERREN, skola äta det högheliga; där skola de förvara det högheliga, såväl spisoffer som syndoffer och skuldoffer ty det är en helig plats.
När prästerna -- som från helgedomen icke strax få begiva sig till den yttre förgården -- hava kommit ditin, skola de där lämna kvar de kläder i vilka de hava gjort tjänst, ty dessa äro heliga; först när de hava iklätt sig andra kläder, få de träda ut på den plats som är för folket.»
När han nu hade slutat uppmätningen av det inre huset, lät han mig gå ut till den port som låg mot öster.
Och han mätte platsen runt omkring.
Han mätte med sin mätstång åt östra sidan: den höll efter mätstången fem hundra stänger runt omkring.
Han mätte åt norra sidan: den höll efter mätstången fem hundra stänger runt omkring.
Han mätte ock åt södra sidan: den höll efter mätstången fem hundra stänger.
Han vände sig mot västra sidan och mätte med mätstången fem hundra stänger.
Åt alla fyra sidorna mätte han platsen.
Den var omgiven av en mur, som utefter platsens längd höll fem hundra stänger och utefter dess bredd fem hundra stänger.
Och den skulle skilja det heliga från det som icke var heligt.
Och han lät mig gå åstad till porten, den port som vette åt öster.
Då såg jag Israels Guds härlighet komma österifrån, och dånet därvid var såsom dånet av stora vatten, och jorden lyste av hans härlighet.
Och den syn som jag då såg var likadan som den jag såg, när jag kom för att fördärva staden; det var en syn likadan som den jag såg vid strömmen Kebar.
Och jag föll ned på mitt ansikte.
Och HERRENS härlighet kom in i huset genom den port som låg mot öster.
Och en andekraft lyfte upp mig och förde mig in på den inre förgården, och jag såg att HERRENS härlighet uppfyllde huset.
Då hörde jag en röst tala till mig från huset, under det att en man stod bredvid mig.
Den sade till mig: Du människobarn, detta är den plats där min tron är, den plats där mina fötter skola stå, där jag vill bo ibland Israels barn evinnerligen.
Och Israels hus skall icke mer orena mitt eviga namn, varken de själva eller deras konungar, med sin trolösa avfällighet, med sina konungars döda kroppar och med sina offerhöjder:
de som satte sin tröskel invid min tröskel, och sin dörrpost vid sidan av min dörrpost, så att allenast muren var mellan mig och dem, och som så orenade mitt heliga namn med de styggelser de bedrevo, varför jag ock förgjorde dem i min vrede.
Men nu skola de skaffa sin trolösa avfällighet och sina konungars döda kroppar långt bort ifrån mig, så att jag kan bo ibland dem evinnerligen.
Men du, människobarn, förkunna nu för Israels barn om detta hus, på det att de må blygas för sina missgärningar.
Må de mäta det härliga byggnadsverket.
Om de då blygas för allt vad de hava gjort, så kungör för dem och teckna för deras ögon upp husets form och inredning, dess utgångar och ingångar, alla dess former och alla stadgar därom, alla dess former och alla lagar därom, så att de akta på hela dess form och alla stadgar därom och göra efter dem.
Detta är lagen om huset: på toppen av berget skall hela dess område runt omkring vara högheligt.
Ja, detta är lagen om huset.
Men dessa voro måtten på altaret i alnar, var aln en handsbredd längre an en vanlig aln: Dess bottenram var en aln hög och en aln bred, och kanten på ramen, runt omkring utmed randen, var ett kvarter hög; detta var altarets underlag.
Avståndet från bottenramen vid marken upp till den nedre avsatsen var två alnar, och bredden var en aln.
Avståndet från den mindre avsatsen upp till den större var fyra alnar, och bredden var en aln.
Altarhärden höll fyra alnar; och från altarhärden stodo de fyra hornen uppåt.
Och altarhärden var tolv alnar lång och tolv alnar bred, så att dess fyra sidor bildade en liksidig fyrkant.
Och avsatsen var fjorton alnar lång och fjorton alnar bred, utefter sina fyra sidor.
Kanten runt omkring den höll en halv aln, och dess bottenram sträckte sig en aln runt omkring.
Och altarets trappsteg vette åt öster.
Och han sade till mig: »Du människobarn, så säger Herren, HERREN: Dessa äro stadgarna om altaret för den dag då det bliver färdigt, så att man kan offra brännoffer och stänka blod därpå.
Då skall du åt de levitiska prästerna giva en ungtjur till syndoffer, åt dem som äro av Sadoks säd, och som få träda fram till mig, säger Herren, HERREN, för att göra tjänst inför mig.
Och du skall taga något av dess blod och stryka på altarets fyra hörn och på avsatsens fyra hörn och på kanten runt omkring; så skall du rena det och bringa försoning för det.
Sedan skall du taga syndofferstjuren, och utanför helgedomen skall den brännas upp på en därtill bestämd plats, som hör till huset.
Och nästa dag skall du föra fram en felfri bock till syndoffer; och man skall rena altaret med den, på samma sätt som man renade det med tjuren.
När du så har fullbordat reningen, skall du föra fram en felfri ungtjur och en felfri vädur av småboskapen.
Dem skall du föra fram inför HERREN, och prästerna skola strö salt på dem och offra dem såsom brännoffer åt HERREN.
Under sju dagar skall du dagligen offra en syndoffersbock; och en ungtjur och en vädur av småboskapen, båda felfria, skall man likaledes offra.
Under sju dagar skall man sålunda bringa försoning för altaret och rena det och inviga det.
Men sedan dessa dagar hava gått till ända, skola prästerna på åttonde dagen och allt framgent offra på altaret edra brännoffer och tackoffer; och jag skall då hava behag till eder, säger Herren, HERREN».
Därefter förde han mig tillbaka mot helgedomens yttre port, den kom vette åt öster; den var nu stängd.
Och HERREN sade till mig: »Denna port skall förbliva stängd och icke mer öppnas, och ingen skall gå in genom den, ty HERREN, Israels Gud, har gått in genom den; därför skall den vara stängd.
Dock skall fursten, eftersom han är furste, få sitta där och hålla måltid inför HERRENS ansikte; han skall då gå in genom portens förhus, och samma väg skall han gå ut igen.»
Därefter förde han mig genom norra porten till platsen framför huset; och jag fick se huru HERRENS härlighet uppfyllde HERRENS hus.
Då föll jag ned på mitt ansikte.
och HERREN sade till mig: Du människobarn, akta på och se med dina ögon, och hör med dina öron allt vad jag nu talar med dig om alla stadgar angående HERRENS hus och om alla lagar som röra det; och giv akt på huru man går in i huset genom alla helgedomens utgångar.
Och säg till Israels hus, det gensträviga: Så säger Herren, HERREN: Nu må det vara nog med alla de styggelser I haven bedrivit, I av Israels hus,
I som haven låtit främlingar med oomskuret hjärta och oomskuret kött komma in i min helgedom och vara där, så att mitt hus har blivit ohelgat, under det att I framburen min spis, fett och blod.
Så har mitt förbund blivit brutet, för att icke nämna alla edra andra styggelser.
I haven icke själva förrättat tjänsten vid mina heliga föremål, utan haven satt andra till att åt eder förrätta tjänsten i min helgedom.
Så säger Herren, HERREN: Ingen främling med oomskuret hjärta och oomskuret kött får komma in i min helgedom, ingen av de främlingar som finnas bland Israels barn.
Utan de leviter som gingo bort ifrån mig, när Israel for vilse de som då själva foro vilse och gingo bort ifrån mig och följde sina eländiga avgudar, de skola bära på sin missgärning
och skola i min helgedom bestrida vakttjänstgöringen vid husets portar och annan tjänstgöring i huset; de skola slakta brännoffer och slaktoffer åt folket, och skola stå inför dem till att betjäna dem.
Eftersom de betjänade dem inför deras eländiga avgudar och så blevo för Israels hus en stötesten till missgärning, därför betygar jag om dem med upplyft hand, säger Herren, HERREN, att de skola få bära på sin missgärning.
De skola icke få nalkas mig, till att förrätta prästerlig tjänst inför mig, eller till att nalkas något av mina heliga föremål, nämligen de högheliga, utan de skola bära på sin skam och på de styggeliga synder som de hava bedrivit.
Och jag skall sätta dem till att förrätta tjänsten i huset vid allt tjänararbete där, allt som där skall utföras.
Men de levitiska präster, nämligen Sadoks söner, som förrättade tjänsten vid min helgedom, när de övriga israeliterna foro vilse och gingo bort ifrån mig, de skola få träda fram till mig för att göra tjänst inför mig; de skola stå inför mitt ansikte för att offra åt mig fett och blod, säger Herren, HERREN.
De skola gå in i min helgedom, och de skola träda fram till mitt bord för att göra tjänst inför mig och förrätta vad som är att förrätta åt mig.
Och när de komma in i den inre förgårdens portar, skola de ikläda sig linnekläder; de få icke hava på sig något av ylle, när de göra tjänst i den inre förgårdens portar och inne i huset.
De skola hava huvudbonader av linne på sina huvuden, och benkläder av linne omkring sina länder; de skola icke omgjorda sig med något som framkallar svett.
Och när de sedan gå ut på den yttre förgården, till folket på den yttre förgården, skola de taga av sig de kläder i vilka de hava gjort tjänst, och skola lämna dem kvar i helgedomens tempelkamrar och ikläda sig andra kläder, för att de icke må göra folket heligt med sina kläder.
De skola icke raka huvudet, men skola icke heller låta håret växa fritt, utan skola klippa sitt huvudhår kort.
Och vin får ingen präst dricka, när han har kommit in på den inre förgården.
En änka eller en frånskild kvinna får han icke taga till hustru åt sig, utan allenast en jungfru av Israels barns släkt; dock får han taga en änka, om hon är änka efter en präst.
Och de skola lära mitt folk att skilja mellan heligt och oheligt och undervisa dem om skillnaden mellan orent och rent.
Och i rättssaker skola de uppträda såsom domare och skola avdöma dem efter mina rätter.
Och mina lagar och stadgar skola de iakttaga vid alla mina högtider, och mina sabbater skola de hålla heliga.
Ingen av dem får orena sig genom att gå in till någon död människa; allenast genom fader eller moder eller son eller dotter eller broder, eller genom en syster som icke har tillhört någon man må han ådraga sig orenhet.
Men när han därefter har blivit ren, skall man räkna för honom ytterligare sju dagar;
och på den dag då han går in i- helgedomen, på den inre förgården, för att göra tjänst i helgedomen, då skall han bära fram ett syndoffer för sig, säger Herren, HERREN.
Och deras arvedel skall bestå däri att jag själv skall vara deras arvedel.
Och I skolen icke giva dem någon besittning i Israel, ty jag själv är deras besittning.
Spisoffret och syndoffret och skuldoffret få de äta, och allt tillspillogivet i Israel skall höra dem till.
Och det första av alla förstlingsfrukter av alla slag, och alla offergärder av alla slag, vadhelst I frambären såsom offergärd, detta skall höra prästerna till; och förstlingen av edert mjöl skolen I giva åt prästen, för att du må bringa välsignelse över ditt hus.
Intet självdött eller ihjälrivet djur, vare sig fågel eller boskapsdjur, få prästerna äta.
Och när I genom lottkastning fördelen landet till arvedel, då skolen I åt HERREN giva en offergärd, en helig del av landet, i längd tjugufem tusen alnar och i bredd tio tusen; detta stycke skall vara heligt till hela sitt omfång runt omkring.
Härav skall tagas till helgedomen en liksidig fyrkant, fem hundra alnar i längd och fem hundra i bredd, runt omkring, och till utmark där runt omkring femtio alnar.
Av det tillmätta stycket skall du alltså avmäta ett område, tjugufem tusen alnar i längd och tio tusen i bredd; där skall helgedomen, det högheliga, ligga.
Detta skall vara en helig del av landet, och det skall tillhöra prästerna, som göra tjänst i helgedomen, dem som få träda fram till att göra tjänst inför HERREN; detta skall vara en plats åt dem för deras hus, så ock en helig plats för helgedomen.
Och ett stycke, tjugufem tusen alnar i längd och tio tusen i bredd, skall tillhöra leviterna, som göra tjänst i huset, såsom deras besittning, med tjugu tempelkamrar.
Och åt staden skolen I giva till besittning ett område, fem tusen alnar i bredd och tjugufem tusen i längd, motsvarande det heliga offergärdsområdet; det skall höra hela Israels hus till.
Och fursten skall på båda sidor om det heliga offergärdsområdet och stadens besittning få ett område, beläget invid det heliga offergärdsområdet och stadens besittning, dels på västra sidan, västerut, dels ock på östra sidan, österut, och I längd motsvarande en stamlotts utsträckning från västra gränsen till östra.
Detta skall han hava till sitt land, till besittning i Israel.
Och mina furstar skola då icke mer förtrycka mitt folk, utan skola låta Israels hus få behålla sitt land efter sina stammar.
Så säger Herren, HERREN: Nu må det vara nog, I Israels furstar.
Skaffen bort våld och förtryck, och öven rätt och rättfärdighet; hören upp att driva mitt folk ifrån hus och hem, säger Herren, HERREN.
Riktig våg, riktig efa, riktigt bat-mått skolen I hava.
Efan och bat-måttet skola hålla samma mått, så att bat-måttet rymmer tiondedelen av en homer, och likaledes efan tiondedelen av en homer; ty efter homern skall man bestämma måtten.
Sikeln skall innehålla tjugu gera; tjugu siklar, tjugufem siklar, femton siklar skall minan innehålla hos eder.
Detta är den offergärd I skolen giva: en sjättedels efa av var homer vete och en sjättedels efa av var homer korn;
vidare den stadgade gärden av olja, räknat efter bat av olja: en tiondedels bat av var kor (som är ett mått på tio bat och lika med en homer, ty tio bat utgöra en homer);
vidare av småboskapen från Israels betesmarker ett djur på vart tvåhundratal, till spisoffer, brännoffer och tackoffer, för att bringa försoning för folket, säger Herren, HERREN.
Allt folket i landet skall vara förpliktat till denna offergärd åt fursten i Israel.
Men fursten skall det åligga att frambära brännoffer, spisoffer och drickoffer på festerna, nymånaderna och sabbaterna, vid alla Israels hus' högtider.
Han skall anskaffa syndoffer, spisoffer, brännoffer och tackoffer till att bringa försoning för Israels hus.
Så säger Herren, HERREN: På första dagen i första månaden skall du taga en felfri ungtjur och rena helgedomen.
Och prästen skall taga något av syndoffrets blod och stryka på husets dörrpost och på altaravsatsens fyra hörn och på dörrposten till den inre förgårdens port.
Så skall du ock göra på sjunde dagen i månaden, om så är, att någon har syndat ouppsåtligen och av fåkunnighet; på detta sätt skolen I bringa försoning för huset.
På fjortonde dagen i första månaden skolen I fira påskhögtid; i sju dagar skolen I hålla högtid, och man skall då äta osyrat bröd.
På den dagen skall fursten för sig själv och för allt folket i landet offra en tjur till syndoffer.
Men sedan, under högtidens sju dagar, skall han dagligen under de sju dagarna offra såsom brännoffer åt HERREN sju tjurar och sju vädurar, alla felfria, och såsom syndoffer en bock dagligen.
Och såsom spisoffer skall han offra en efa till var tjur och en efa till var vädur, jämte en hin olja till var efa.
På femtonde dagen i sjunde månaden skall han vid högtiden frambära likadana offer under de sju dagarna, likadana syndoffer, brännoffer och spisoffer och lika mycket olja.
Så säger Herren, HERREN: Den inre förgårdens port, den som vetter åt öster, skall vara stängd under de sex arbetsdagarna, men på sabbatsdagen skall den öppnas; likaledes skall den öppnas på nymånadsdagen.
Och då skall fursten utifrån gå in genom portens förhus och ställa sig vid portens dörrpost; och när prästerna offra hans brännoffer och hans tackoffer, skall han tillbedja på portens tröskel och därefter gå ut.
Men porten skall icke stängas förren om aftonen.
Och folket i landet skall på sabbater och nymånader tillbedja inför HERREN vid ingången till samma port.
Och brännoffret som fursten skall frambära åt HERREN skall på sabbatsdagen utgöras av sex felfria lamm och en felfri vädur.
Och såsom spisoffer skall han frambära en efa till väduren, men till lammen såsom spisoffer så mycket han vill giva, jämte en hin olja till var efa.
Men på nymånadsdagen skall han frambära en felfri ungtjur, sex lamm och en vädur, allasammans felfria.
Och såsom spisoffer skall han offra en efa till tjuren och en efa till väduren, och till lammen så mycket han vill anskaffa, jämte en hin olja till var efa.
Och när fursten vill gå in, skall han gå in genom portens förhus, och samma väg skall han gå ut igen.
Men när folket i landet kommer inför HERRENS ansikte vid högtiderna, då skall den som har gått in genom norra porten för att tillbedja gå ut genom södra porten, och den som har gått in genom södra porten skall gå ut genom norra porten; ingen skall gå tillbaka genom samma port som han har kommit in igenom, utan man skall gå ut genom den motsatta.
Och fursten skall gå in tillsammans med de andra, när de gå in; och när de gå ut, skola de gå ut tillsammans.
Men vid fester och högtider skall spisoffret utgöras av en efa till var tjur och en efa till var vädur, och till lammen av så mycket han vill giva, jämte en hin olja till var efa.
Och när fursten vill offra ett frivilligt offer, vare sig ett brännoffer eller ett tackoffer såsom frivilligt offer åt HERREN, då skall man öppna åt honom den port som vetter åt öster, och han skall offra sitt brännoffer och sitt tackoffer alldeles så, som han plägar offra på sabbatsdagen; och därefter skall han gå ut och sedan han har gått ut, skall man stänga porten.
Du skall dagligen offra såsom brännoffer åt HERREN ett felfritt årsgammalt lamm; var morgon skall du offra ett sådant.
Och såsom spisoffer skall du därtill offra var morgon en sjättedels efa, så ock en tredjedels hin olja för att fukta mjölet -- detta såsom spisoffer åt HERREN, såsom evärdlig rätt för beständigt.
I skolen offra lammet och spisoffret och oljan var morgon såsom dagligt brännoffer.
Så säger Herren, HERREN: Om fursten giver någon av sina söner en gåva, så bliver det dennes arvedel, det skall höra hans söner till; de skola besitta det såsom arv.
Men om han av sin arvedel giver något såsom gåva åt någon av sina tjänare, så skall detta tillhöra denne intill friåret; då skall det återgå till fursten.
Hans arvedel är det ju, och hans söner skall det tillfalla.
Fursten må icke taga något av folkets arvedel och så kränka den i deras besittningsrätt; allenast av sin egen besittning må han giva arvedelar åt sina söner, för att ingen av mitt folk skall bliva undanträngd från sin särskilda besittning.
Och han förde mig genom den ingång som låg vid sidan av porten till de heliga tempelkamrar som voro bestämda för prästerna, och som vette åt norr; och jag såg att där var en plats längst uppe i väster.
Och han sade till mig: »Detta är den plats där prästerna skola koka skuldoffret och syndoffret, och där de skola baka spisoffret, för att icke behöva bära ut det på den yttre förgården och så göra folket heligt.»
Därefter lät han mig gå ut på den yttre förgården och förde mig omkring till förgårdens fyra hörn; och jag såg då att i vart och ett av förgårdens hörn fanns en gård.
I förgårdens fyra hörn funnos kringstängda gårdar, fyrtio alnar långa och trettio alnar breda; dessa fyra hörngårdar voro lika stora.
Och runt omkring inuti dem gick en mur, runt omkring i alla fyra; och nedtill vid muren runt omkring hade man inrättat eldstäder till kokning.
Och han sade till mig: »Detta är de kök i vilka husets tjänare skola koka folkets slaktoffer.»
Därefter förde han mig tillbaka till husets ingång, och där fick jag se vatten rinna fram under husets tröskel på östra sidan, ty husets framsida låg mot öster; och vattnet flöt ned under husets södra sidovägg, söder om altaret.
Sedan lät han mig gå ut genom norra porten och förde mig omkring på en yttre väg till den yttre porten, den som vette åt öster.
Där fick jag se vatten välla fram på södra sidan.
Sedan gick mannen, med ett mätsnöre i handen, ett stycke mot öster och mätte därvid upp tusen alnar och lät mig så gå över vattnet, och vattnet räckte mig där till fotknölarna.
Åter mätte han upp tusen alnar och lät mig så gå över vattnet, och vattnet räckte mig där till knäna.
Åter mätte han upp tusen alnar och lät mig så gå över vattnet, som där räckte mig upp till länderna.
Ännu en gång mätte han upp tusen alnar, och nu var det en ström som jag icke kunde gå över.
Ty vattnet gick så högt att man måste simma; det var en ström som man icke kunde gå över.
Och han sade till mig: »Nu har du ju sett det, du människobarn?»
Sedan förde han mig tillbaka upp på strömmens strand.
Och när han hade fört mig dit tillbaka, fick jag se träd i stor myckenhet stå på strömmens strand, på båda sidor.
Och han sade till mig: »Detta vatten rinner fram mot Östra kretsen och flyter ned på Hedmarken och faller därefter ut i havet.
Vattnet som fick bryta fram går alltså till havet, och så bliver vattnet där sunt.
Och överallt dit den dubbla strömmen kommer, där upplivas alla levande varelser som röra sig i stim, och fiskarna bliva där mycket talrika; ty när detta vatten kommer dit, bliver havsvattnet sunt, och allt får liv, där strömmen kommer.
Och fiskare skola stå utmed den från En-Gedi ända till En-Eglaim, och såsom ett enda fiskeläge skall den sträckan vara.
Där skola finnas fiskar av olika slag i stor myckenhet, alldeles såsom i Stora havet.
Men gölar och dammar där skola icke bliva sunda, utan skola tjäna till saltberedning.
Och vid strömmen, på dess båda stränder, skola allahanda fruktträd växa upp, vilkas löv icke skola vissna, och vilkas frukt icke skall taga slut, utan var månad skola träden bara ny frukt, ty deras vatten kommer från helgedomen.
Och deras frukter skola tjäna till föda och deras löv till läkedom.»
Så säger Herren, HERREN: Dessa äro de gränser efter vilka I skolen utskifta landet såsom arvedel åt Israels tolv stammar (varvid Josef får mer än en lott).
I skolen få det till arvedel, den ene såväl som den andre, därför att jag med upplyft hand har lovat att giva det åt edra fader; så skall nu detta land tillfalla eder såsom arvsegendom.
Detta skall vara landets gräns på norra sidan: från Stora havet längs Hetlonsvägen, dit fram där vägen går till Sedad,
Hamat, Berota, Sibraim, som ligger mellan Damaskus' och Hamat områden, det mellersta Haser, som ligger invid Haurans område.
Så skall gränsen gå från havet till Hasar-Enon vid Damaskus' område och vidare allt längre norrut och upp mot Hamats område.
Detta är norra sidan.
Och på östra sidan skall gränsen begynna mellan Hauran och Damaskus och gå mellan Gilead och Israels land och utgöras av Jordan; från nordgränsen nedåt, utmed Östra havet, skolen I mäta ut den.
Detta är östra sidan.
Och på sydsidan, söderut, skall gränsen gå från Tamar till Meribots vatten vid Kades, till bäcken, fram till Stora havet.
Detta är sydsidan, söderut.
Och på västra sidan skall gränsen utgöras av Stora havet och gå från sydgränsen till en punkt mitt emot det ställe där vägen går till Hamat.
Detta är västra sidan.
Och I skolen utskifta detta land åt eder efter Israels stammar.
I skolen utdela det genom lottkastning till arvedel åt eder själva och åt främlingarna som bo ibland eder och hava fött barn ibland eder.
Ty de skola av eder hållas lika med infödda israeliter; de skola tillfalla eder såsom en arvedel bland Israels stammar.
I den stam där främlingen bor, där skolen I giva honom hans arvedel, säger Herren, HERREN.
Och dessa äro namnen på stammarna.
Vid norra gränsen längs efter Hetlonsvägen, dit fram där vägen går till Hamat, vidare bort mot Hasar-Enan -- med Damaskus' område jämte Hamat i norr -- där skall Dan hava en lott, så att hela sträckan från östra sidan till västra tillhör honom.
Och närmast Dans område skall Aser hava en lott, från östra sidan till västra.
Och närmast Asers område skall Naftali hava en lott, från östra sidan till västra.
Och närmast Naftalis område skall Manasse hava en lott, från östra sidan till västra.
Och närmast Manasses område skall Efraim hava en lott, från östra sidan till västra.
Och närmast Efraims område skall Ruben hava en lott, från östra sidan till västra.
Och närmast Rubens område skall Juda hava en lott, från östra sidan till västra.
Och närmast Juda område skall från östra sidan till västra sträcka sig det offergärdsområde som I skolen giva såsom gärd, tjugufem tusen alnar i bredd, och i längd lika med en stamlotts längd från östra sidan till västra; och helgedomen skall ligga där i mitten.
Det offergärdsområde som I skolen giva såsom gärd åt HERREN skall vara i längd tjugufem tusen alnar och i bredd tio tusen.
Och av detta heliga offergärdsområde skall ett stycke tillhöra prästerna, i norr tjugufem tusen alnar, i väster tio tusen i bredd, i öster likaledes tio tusen i bredd och i söder tjugufem tusen i längd; och HERRENS helgedom skall ligga där i mitten.
Det skall tillhöra prästerna, dem som hava blivit helgade bland Sadoks söner, dem som hava förrättat tjänsten åt mig, och som icke, såsom leviterna gjorde, foro vilse, när de övriga israeliterna foro vilse.
Därför skall en särskild offergärdsdel av den från landet avtagna offergärden tillhöra dem såsom ett högheligt område invid leviternas.
Men leviterna skola få ett område motsvarande prästernas, i längd tjugufem tusen alnar och i bredd tiotusen -- längden överallt tjugufem tusen och bredden tio tusen.
Och de få icke sälja något därav; det bästa landet må man icke byta bort eller eljest överlåta åt någon annan, ty det är helgat åt HERREN.
Men de fem tusen alnar som bliva över på bredden invid de tjugufem tusen skola utgöra ett icke heligt område för staden, dels till att bo på, dels såsom utmark; och staden skall ligga där i mitten.
Och detta är måttet på den: norra sidan fyra tusen fem hundra alnar, södra sidan fyra tusen fem hundra, på östra sidan fyra tusen fem hundra, och västra sidan fyra tusen fem hundra.
Och staden skall hava en utmark, som norrut är två hundra femtio alnar, söderut två hundra femtio, österut två hundra femtio och västerut två hundra femtio.
Och vad som bliver över på långsidan utmed det heliga offergärdsområdet, nämligen tio tusen alnar österut och tio tusen västerut -- ty det skall sträcka sig utmed det heliga offergärdsområdet -- av detta skall avkastningen tjäna till föda åt stadens bebyggare.
Alla stadens bebyggare från alla Israels stammar skola bruka det.
Hela offergärdsområdet skall alltså vara tjugufem tusen alnar i längd och tjugufem tusen i bredd; det heliga offergärdsområde som I given såsom gärd skall bilda en fyrkant, stadens besittning inberäknad.
Och fursten skall få vad som bliver över på båda sidor om det heliga offergärdsområdet och stadens besittning, nämligen landet invid det tjugufem tusen alnar breda offergärdsområdet, ända till östra gränsen, och likaledes västerut landet utefter det tjugufem tusen alnar breda området, ända till västra gränsen.
Dessa områden, motsvarande stamlotterna, skola tillhöra fursten.
Och det heliga offergärdsområdet med det heliga huset skall ligga mitt emellan dem.
Med sin gräns å ena sidan mot leviternas besittning, å andra sidan mot stadens, skall detta område ligga mitt emellan furstens besittningar.
Och furstens besittningar skola ligga mellan Juda område och Benjamins område.
Därefter skola de återstående stammarna komma.
Först skall Benjamin hava en lott från östra sidan till västra.
Och närmast Benjamins område skall Simeon hava en lott, från östra sidan till västra.
Och närmast Simeons område skall Isaskar hava en lott, från östra sidan till västra.
Och närmast Isaskars område skall Sebulon hava en lott, från östra sidan till västra.
Och närmast Sebulons område skall Gad hava en lott, från östra sida till västra.
Och närmast Gads område, på dess sydsida, söderut, skall gränser gå från Tamar över Meribas vatten vid Kades till bäcken, fram emot Stora havet.
Detta är det land som I genom lottkastning skolen utdela åt Israels stammar till arvedel; och detta skall vara deras stamlotter, säger Herren, HERREN.
Och följande utgångar skall staden hava: På norra sidan skall den hålla ett mått av fyra tusen fem hundra alnar,
och av stadens portar, uppkallade efter Israels stammars namn, skola tre ligga i norr: den första Rubens port, den andra Juda port, den tredje Levi port.
Och på östra sidan skall den ock. hålla fyra tusen fem hundra alnar och hava tre portar: den första Josefs port, den andra Benjamins port, den tredje Dans port.
Sammalunda skall ock södra sidan hålla ett mått av fyra tusen fem hundra alnar och hava tre portar: den första Simeons port, den andra Isaskars port, den tredje Sebulons port.
Västra sidan skall hålla fyra tusen fem hundra alnar och hava tre portar: den första Gads port, den andra Asers port, den tredje Naftali port.
Runt omkring skall den hålla aderton tusen alnar.
Och stadens namn skall allt framgent vara: Här är HERREN.
I Jojakims, Juda konungs, tredje regeringsår kom Nebukadnessar, konungen i Babel, mot Jerusalem och belägrade det.
Och Herren gav Jojakim, Juda konung, i hans hand, så ock en del av kärlen i Guds hus; och han förde dem till Sinears land, in i sin guds hus.
Och kärlen förde han in i sin guds skattkammare.
Och konungen befallde Aspenas, sin överste hovman, att han skulle av Israels barn taga till sig ynglingar av konungslig släkt eller av förnäm börd,
sådana som icke hade något lyte, utan voro fagra att skåda och utrustade med förstånd till att inhämta allt slags visdom, kloka och läraktiga ynglingar, som kunde bliva dugliga att tjäna i konungens palats; dem skulle han låta undervisa i kaldéernas skrift och tungomål.
Och konungen bestämde åt dem ett visst underhåll för var dag, av konungens egen mat och av det vin han själv drack, och befallde att man skulle uppfostra dem i tre år; när den tiden vore förliden, skulle de få göra tjänst hos konungen.
Bland dessa voro nu Daniel, Hananja, Misael och Asarja, av Juda barn.
Men överste hovmannen gav dem andra namn: Daniel kallade han Beltesassar, Hananja Sadrak, Misael Mesak och Asarja Abed-Nego.
Men Daniel lät sig angeläget vara att icke orena sig med konungens mat eller med vinet som denne drack av; och han bad överste hovmannen att han icke skulle nödgas orena sig.
Och Gud lät Daniel finna nåd och barmhärtighet inför överste hovmannen.
Men överste hovmannen sade till Daniel: »Jag fruktar att min herre, konungen, som har beställt om eder mat och dryck, då skall finna edra ansikten magrare än de ynglingars som äro jämnåriga med eder, och att I så skolen draga skuld över mitt huvud inför konungen.»
Då sade Daniel till hovmästaren som av överste hovmannen hade blivit satt till att hava uppsikt över Daniel, Hananja, Misael och Asarja:
»Gör ett försök med dina tjänare i tio dagar, och låt giva oss grönsaker att äta och vatten att dricka.
Sedan må du jämföra vårt utseende med de ynglingars som hava ätit av konungens mat; och efter vad du då anser må du göra med dina tjänare.»
Och han lyssnade till denna deras begäran och gjorde ett försök med dem i tio dagar.
Och efter de tio dagarnas förlopp befunnos de vara fagrare att skåda och stadda vid bättre hull än alla de ynglingar som hade ätit av konungens mat.
Då lät hovmästaren dem allt fortfarande slippa den mat som hade varit bestämd för dem och det vin som de skulle hava druckit, och gav dem grönsaker.
Åt dessa fyra ynglingar gav nu Gud kunskap och insikt i allt slags skrift och visdom; och Daniel fick förstånd på alla slags syner och drömmar.
Och när den tid var förliden, efter vilken de, enligt konungens befallning, skulle föras fram för honom, blevo de av överste hovmannen förda inför Nebukadnessar
När då konungen talade med dem, fanns bland dem alla ingen som kunde förliknas med Daniel, Hananja, Misael och Asarja; och de fingo så göra tjänst hos konungen.
Och närhelst konungen tillfrågade dem i en sak som fordrade vishet i förståndet, fann han dem vara tio gånger klokare än någon av de spåmän och besvärjare som funnos i hela hans rike.
Och Daniel fortfor så intill konung Kores' första regeringsår.
I sitt andra regeringsår hade Nebukadnessar drömmar av vilka han blev orolig till sinnes, och sömnen vek bort ifrån honom.
Då lät konungen tillkalla sina spåmän, besvärjare, trollkarlar och kaldéer, för att de skulle giva konungen till känna vad han hade drömt, och de kommo och trädde fram för konungen.
Och konungen sade till dem: »Jag har haft en dröm, och jag är orolig till sinnes och ville veta vad jag har drömt.»
Då talade kaldéerna till konungen på arameiska: »Må du leva evinnerligen, o konung!
Förtälj drömmen för dina tjänare, så skola vi meddela uttydningen.»
Konungen svarade och sade till kaldéerna: »Nej, mitt oryggliga beslut är, att om I icke sägen mig drömmen och dess uttydning, skolen I huggas i stycken, och edra hus skola göras till platser för orenlighet.
Men om I meddelen drömmen och dess uttydning, så skolen I få gåvor och skänker och stor ära av mig.
Meddelen mig alltså nu drömmen och dess uttydning.»
De svarade för andra gången och sade: »Konungen må förtälja drömmen för sina tjänare, så skola vi meddela uttydningen.»
Konungen svarade och sade: »Jag märker nogsamt att I viljen vinna tid, eftersom I sen att mitt beslut är oryggligt,
att om I icke sägen mig drömmen, domen över eder icke kan bliva annat än en.
Ja, I haven kommit överens om att inför mig föra lögnaktigt och bedrägligt tal, i hopp att tiderna skola förändra sig.
Sägen mig alltså nu vad jag har drömt, så märker jag att I ock kunnen meddela mig uttydningen därpå.»
Då svarade kaldéerna konungen och sade: »Det finnes ingen människa på jorden, som förmår meddela konungen det som han vill veta; aldrig har ju heller någon konung, huru stor och mäktig han än var, begärt sådant som detta av någon spåman eller besvärjare eller kaldé.
Ty det som konungen begär är alltför svårt, och ingen finnes, som kan meddela konungen det, förutom gudarna; och de hava icke sin boning ibland de dödliga.
Då blev konungen vred och mycket förtörnad och befallde att man skulle förgöra alla de vise i Babel.
När alltså påbudet härom hade blivit utfärdat och man skulle döda de vise, sökte man ock efter Daniel och hans medbröder för att döda dem.
Då vände sig Daniel med kloka och förståndiga ord till Arjok, översten för konungens drabanter, vilken hade dragit ut för att döda de vise i Babel.
Han tog till orda och frågade Arjok, konungens hövitsman: »Varför har detta stränga påbud blivit utfärdat av konungen?»
Då omtalade Arjok för Daniel vad som var på färde.
Och Daniel gick in och bad konungen att tid måtte beviljas honom, så skulle han meddela konungen uttydningen.
Därefter gick Daniel hem och omtalade för Hananja, Misael och Asarja, sina medbröder, vad som var på färde,
och han uppmanade dem att bedja himmelens Gud om förbarmande, så att denna hemlighet bleve uppenbarad, på det att icke Daniel och hans medbröder måtte förgöras tillika med de övriga vise Babel.
Då blev hemligheten uppenbarad för Daniel i en syn om natten.
Och Daniel lovade himmelens Gud därför;
Daniel hov upp sin röst och sade: »Lovat vare Guds namn från evighet till evighet!
Ty vishet och makt höra honom till.
Han låter tider och stunder omskifta, han avsätter konungar och tillsätter konungar, han giver åt de visa deras vishet och åt de förståndiga deras förstånd.
Han uppenbarar det som är djupt och förborgat, han vet vad i mörkret är, och hos honom bor ljuset.
Dig, mina fäders Gud, tackar och prisar jag för att du har givit mig vishet och förmåga, och för att du nu har uppenbarat för mig det vi bådo dig om; ty det som konungen ville veta har du uppenbarat för oss.»
I följd härav gick Daniel in till Arjok, som av konungen hade fått befallning att förgöra de vise i Babel; han gick åstad och sade till honom så: »De vise i Babel må du icke förgöra.
För mig in till konungen, så skall jag meddela konungen uttydningen.»
Då förde Arjok med hast Daniel inför konungen och sade till honom så: »Jag har bland de judiska fångarna funnit en man som kan säga konungen uttydningen.»
Konungen svarade och sade till Daniel, som hade fått namnet Beltesassar: »Förmår du säga mig den dröm som jag har haft och dess uttydning?»
Daniel svarade konungen och sade: »Den hemlighet som konungen begär att få veta kunna inga vise, besvärjare, spåmän eller stjärntydare meddela konungen.
Men det finnes en Gud i himmelen, som kan uppenbara hemligheter, och han har låtit konung Nebukadnessar veta vad som skall ske i kommande dagar.
Detta var din dröm och den syn du hade på ditt läger:
När du, o konung, låg på ditt läger, uppstego hos dig tankar på vad som skall ske i framtiden; och han som uppenbarar hemligheter lät dig veta vad som skall ske.
Och för mig har denna hemlighet blivit uppenbarad, icke i kraft av någon vishet som jag äger framför alla andra levande varelser, utan på det att uttydningen må bliva kungjord för konungen, så att du förstår ditt hjärtas tankar.
Du, o konung, såg i din syn en stor bildstod stå framför dig, och den stoden var hög och dess glans övermåttan stor, och den var förskräcklig att skåda.
Bildstodens huvud var av bästa guld, dess bröst och armar voro av silver, dess buk och länder av koppar; dess ben voro av järn,
dess fötter delvis av järn och delvis av lera.
Medan du nu betraktade den, blev en sten lösriven, dock icke genom människohänder, och den träffade bildstoden på fötterna, som voro av järn och lera, och krossade dem.
Då blev på en gång alltsammans krossat, järnet, leran, kopparen, silvret och guldet, och det blev såsom agnar på en tröskloge om sommaren, och vinden förde bort det, så att man icke mer kunde finna något spår därav.
Men av stenen som hade träffat bildstoden blev ett stort berg, som uppfyllde hela jorden.
Detta var drömmen; och vi vilja nu säga konungen uttydningen:
Du, o konung, konungarnas konung, åt vilken himmelens Gud har givit rike, väldighet, makt och ära,
och i vilkens hand han har givit människors barn och djuren på marken och fåglarna under himmelen, varhelst varelser bo, och som han har satt till herre över allasammans, du är det gyllene huvudet.
Men efter dig skall uppstå ett annat rike, ringare än ditt, och därefter ännu ett tredje rike, ett som är av koppar, och det skall råda över hela jorden.
Ett fjärde rike skall ock uppstå och vara starkt såsom järn, ty järnet krossar och sönderslår ju allt; och såsom järnet förstör allt annat, så skall ock detta krossa och förstöra.
Men att du såg fötterna och tårna vara delvis av krukmakarlera och delvis av järn, det betyder att det skall vara ett söndrat rike, dock så att det har något av järnets fasthet, ty du såg ju järn vara där, blandat med lerjord.
Och att tårna på fötterna voro delvis av järn och delvis av lera, det betyder att riket skall vara delvis starkt och delvis svagt.
Och att du såg järnet vara blandat med lerjord, det betyder att väl en beblandning där skall äga rum genom människosäd, men att delarna likväl icke skola hålla ihop med varandra, lika litet som järn kan förbinda sig med lera.
Men i de konungarnas dagar skall himmelens Gud upprätta ett rike som aldrig i evighet skall förstöras och vars makt icke skall bliva överlämnad åt något annat folk.
Det skall krossa och göra en ände på alla dessa andra riken, men självt skall det bestå evinnerligen;
ty du såg ju att en sten blev lösriven från berget, dock icke genom människohänder, och att den krossade järnet, kopparen, leran, silvret och guldet.
Så har en stor Gud uppenbarat för konungen vad som skall ske i framtiden, och drömmen är viss, och dess uttydning är tillförlitlig.»
Då föll konung Nebukadnessar på sitt ansikte och tillbad inför Daniel, och befallde att man skulle offra åt honom spisoffer och rökoffer.
Och konungen svarade Daniel och sade: »I sanning, eder Gud är en Gud över andra gudar och en herre över konungar och en uppenbarare av hemligheter, eftersom du har kunnat uppenbara denna hemlighet.»
Därefter upphöjde konungen Daniel och gav honom många stora skänker och satte honom till herre över hela Babels hövdingdöme och till högste föreståndare för alla de vise i Babel.
Och på Daniels bön förordnade konungen Sadrak, Mesak och Abed-Nego att förvalta Babels hövdingdöme; men Daniel själv stannade vid konungens hov.
Konung Nebukadnessar lät göra en gyllene bildstod, sextio alnar hög och sex alnar bred; den lät han ställa upp på Duraslätten i Babels hövdingdöme.
Och konung Nebukadnessar sände åstad och lät församla satraper, landshövdingar och ståthållare, fogdar, skattmästare, domare, lagtolkare och alla andra makthavande i hövdingdömena, för att de skulle komma till invigningen av den bildstod som konung Nebukadnessar hade låtit ställa upp.
Då församlade sig satraperna, landshövdingarna och ståthållarna, fogdarna, skattmästarna, domarna, lagtolkarna och alla andra makthavande i hövdingdömena till invigningen av den bildstod som konung Nebukadnessar hade låtit ställa upp och när de så stodo framför den bildstod som Nebukadnessar hade låtit ställa upp,
utropade en härold med hög röst: »Detta vare eder befallt, I folk och stammar och tungomål:
När I hören ljudet av horn, pipor, cittror, sambukor, psaltare, säckpipor och allahanda andra instrumenter, skolen I falla ned och tillbedja den gyllene bildstod som konung Nebukadnessar har låtit ställa upp.
Men den som icke faller ned och tillbeder, han skall i samma stund kastas i den brinnande ugnen.»
Så snart nu allt folket hörde ljudet av horn, pipor, cittror, sambukor, psaltare och allahanda andra instrumenter, föllo de alltså ned, alla folk och stammar och tungomål, och tillbådo den gyllene bildstod som konung Nebukadnessar hade låtit ställa upp.
Men strax därefter kommo några kaldeiska män fram och anklagade judarna.
De togo till orda och sade till konung Nebukadnessar: Må du leva evinnerligen, o konung!
Du, o konung, har givit befallning att alla människor, när de hörde ljudet av horn, pipor, cittror, sambukor, psaltare, säckpipor och allahanda andra instrumenter, skulle falla ned och tillbedja den gyllene bildstoden,
och att var och en som icke fölle ned och tillbåde skulle kastas i den brinnande ugnen.
Men nu äro här några judiska män, Sadrak, Mesak och Abed-Nego, vilka du har förordnat att förvalta Babels hövdingdöme.
Dessa män hava icke aktat på dig, o konung.
De dyrka icke dina gudar; och den gyllene bildstod som du har låtit ställa upp tillbedja de icke.»
Då befallde Nebukadnessar i vrede och förbittring att man skulle föra fram Sadrak, Mesak och Abed-Nego.
Och när man hade fört fram männen inför konungen,
talade Nebukadnessar till dem och sade: »Är det av förakt som I, Sadrak, Mesak och Abed-Nego, icke dyrken mina gudar och icke tillbedjen den gyllene bildstod som jag har låtit ställa upp?
Välan, allt må vara gott, om I ären redo, att när I hören ljudet av horn, pipor, cittror, sambukor, psaltare, säckpipor och allahanda andra instrumenter, falla ned och tillbedja den bildstod som jag har låtit göra.
Men om I icke tillbedjen, då skolen I i samma stund bliva kastade i den brinnande ugnen; och vilken är väl den gud som då kan rädda eder ur min hand?»
Då svarade Sadrak, Mesak och Abed-Nego och sade till konungen: »O Nebukadnessar, vi behöva icke giva dig något svar på detta.
Om vår Gud, den som vi dyrka, förmår rädda oss, så skall han ock rädda oss ur den brinnande ugnen och ur din hand, o konung.
Men om han icke vill det, så må du veta, o konung, att vi ändå icke dyrka dina gudar, och att vi icke vilja tillbedja den gyllene bildstod som du har låtit ställa upp.»
Då uppfylldes Nebukadnessar av vrede mot Sadrak, Mesak och Abed-Nego, så att hans ansikte förvandlades.
Och han hov upp sin röst och befallde att man skulle göra ugnen sju gånger hetare, än man någonsin hade sett den vara.
Och några handfasta män i hans här fingo befallning att binda Sadrak, Mesak och Abed-Nego och kasta dem i den brinnande ugnen.
Så blevo dessa med sina underkläder, livrockar, mössor och andra kläder bundna och kastade i den brinnande ugnen.
Men eftersom konungens befallning hade varit så sträng, och ugnen därför hade blivit så övermåttan starkt upphettad, blevo de män som förde Sadrak, Mesak och Abed-Nego ditupp själva dödade av eldslågorna,
vid det att de tre männen Sadrak, Mesak och Abed-Nego bundna kastades ned i den brinnande ugnen.
Då blev konung Nebukadnessar förskräckt och stod upp med hast och frågade sina rådsherrar och sade: »Var det icke tre män som vi läto kasta bundna i elden?
De svarade och sade till konungen: »Jo förvisso, o konung.»
Han fortfor och sade: »Och ändå ser jag nu fyra män, som gå lösa och lediga inne i elden, och ingen skada har skett dem; och den fjärde ser så ut, som vore han en gudason.»
Därefter trädde Nebukadnessar fram till öppningen på den brinnande ugnen och hov upp sin röst och sade: »Sadrak, Mesak och Abed-Nego, I den högste Gudens tjänare kommen hitut.»
Då gingo Sadrak, Mesak och Abed-Nego ut ur elden.
Och satraperna, landshövdingarna och ståthållarna och konungens rådsherrar församlade sig där, och fingo då se att elden icke hade haft någon makt över männens kroppar, och att håret på deras huvuden icke var svett, och att deras kläder icke hade blivit skadade; ja, man kunde icke ens känna lukten av något bränt på dem.
Då hov Nebukadnessar upp sin röst och sade: »Lovad vare Sadraks, Mesaks och Abed-Negos Gud, som sände sin ängel och räddade sina tjänare, vilka så förtröstade på honom, att de överträdde konungens befallning och vågade sina liv för att icke nödgas dyrka eller tillbedja någon annan gud än sin egen Gud!
Och härmed giver jag nu befallning att vilken som helst av alla folk och stammar och tungomål, som säger något otillbörligt om Sadraks, Mesaks och Abed-Negos Gud, han skall huggas i stycken, och hans hus skall göras till en plats för orenlighet; ty ingen gud finnes, som så kan hjälpa som denne.
Därefter lät konungen Sadrak, Mesak och Abed-Nego komma till stor ära och makt i Babels hövdingdöme.
Konung Nebukadnessar till alla folk och stammar och tungomål som finnas på hela jorden.
Mycken frid vare med eder!
Jag har funnit för gott att härmed kungöra de tecken och under som den högste Guden har gjort med mig.
Ty stora äro förvisso hans tecken, och mäktiga äro hans under.
Hans rike är ett evigt rike, och hans välde varar från släkte till släkte.
Jag, Nebukadnessar, satt i god ro i mitt hus och levde lycklig i mitt palats.
Då hade jag en dröm som förskräckte mig; jag ängslades genom drömbilder på mitt läger och genom en syn som jag såg.
Därför gav jag befallning att man skulle hämta alla de vise i Babel till mig, för att de skulle säga mig drömmens uttydning.
Så kommo nu spåmännen, besvärjarna, kaldéerna och stjärntydarna, och jag förtäljde drömmen för dem, men de kunde icke säga mig dess uttydning.
Slutligen kom ock Daniel inför mig, han som hade fått namnet Beltesassar efter min guds namn, och i vilken heliga gudars ande är; och jag förtäljde drömmen för honom sålunda:
»Beltesassar, du som är den överste bland spåmännen, du om vilken jag vet att heliga gudars ande är i dig, och att ingen hemlighet är dig för svår, säg mig vad jag såg i min dröm, och vad den betyder.
Detta var den syn jag hade på mitt läger: Jag såg i min syn ett träd stå mitt på jorden, och det var mycket högt.
Ja, stort och väldigt var trädet, och så högt att det räckte upp till himmelen och syntes allt intill jordens ända.
Dess lövverk var skönt, och de bar mycken frukt, så att det hade föda åt alla.
Markens djur funno skugga därunder, och himmelens fåglar bodde på dess grenar, och allt kött hade sin föda därav.
Vidare såg jag, i den syn jag hade på mitt läger, huru en helig ängel steg ned från himmelen.
Han ropade med hög röst och sade: 'Huggen ned trädet och skären av dess grenar, riven bort dess lövverk och förströn dess frukt, så att djuren som ligga därunder fara sin väg och fåglarna flyga bort ifrån dess grenar.
Dock må stubben med rötterna lämnas kvar i jorden, bunden med kedjor av järn och koppar, bland markens gräs; av himmelens dagg skall han vätas och hava sin lott med djuren bland markens örter.
Hans hjärta skall förvandlas, så att det icke mer är en människas, och ett djurs hjärta skall givas åt honom, och sju tider skola så gå fram över honom.
Så är det förordnat genom änglarnas rådslut, och så är det befallt om denna sak av de heliga, för att de levande skola besinna att den Högste råder över människors riken och giver dem åt vem han vill, ja, upphöjer den lägste bland människor till att härska över dem.'
Sådan var den dröm som jag, konung Nebukadnessar, hade.
Och du, Beltesassar, må nu säga uttydningen; ty ingen av de vise i mitt rike kan säga mig uttydningen, men du kan det väl, ty heliga gudars ande är i dig.»
Då stod Daniel, som också hade namnet Beltesassar, en stund häpen, uppfylld av oroliga tankar.
Men konungen tog åter till orda och sade: »Beltesassar, låt icke drömmen och vad den betyder förskräcka dig.
Beltesassar svarade och sade: »Min herre, o att drömmen gällde dem som hata dig, och dess betydelse dina fiender!
Trädet som du såg, vilket var så stort och väldigt och så högt att det räckte upp till himmelen och syntes över hela jorden,
och som hade ett så skönt lövverk och bar mycken frukt, så att det hade föda åt alla, trädet under vilket markens djur bodde, och på vars grenar himmelens fåglar hade sina nästen,
det är du själv, o konung, du som har blivit så stor och väldig, du vilkens storhet har vuxit, till dess att den har nått upp till himmelen, och vilkens välde sträcker sig till jordens ända.
Men att konungen såg en helig ängel stiga ned från himmelen, vilken sade: 'Huggen ned trädet och förstören det; dock må stubben med rötterna lämnas kvar i jorden, bunden med kedjor av järn och koppar, bland markens gräs; av himmelens dagg skall han vätas och hava sin lott med markens djur, till dess att sju tider hava gått fram över honom',
detta betyder följande, o konung, och detta är den Högstes rådslut, som har drabbat min herre konungen:
Du skall bliva utstött från människorna och nödgas bo ibland markens djur och äta gräs såsom en oxe och vätas av himmelens dagg; och sju tider skola så gå fram över dig, till dess du besinnar att den Högste råder över människors riken och giver dem åt vem han vill.
Men att det befalldes att trädets stubbe med rötterna skulle lämnas kvar, det betyder att du skall återfå ditt rike, när du har besinnat att det är himmelen som har makten.
Därför, o konung, må du låta mitt råd täckas dig: gör dig fri ifrån dina synder genom att göra gott, och ifrån dina missgärningar genom att öva barmhärtighet mot de fattiga, om till äventyrs din lycka så kunde bliva beståndande.»
Allt detta drabbade också konung Nebukadnessar.
Tolv månader därefter, när konungen en gång gick omkring på taket av det kungliga palatset i Babel,
hov han upp sin röst och sade: »Se, detta är det stora Babel, som jag har byggt upp till ett konungasäte genom min väldiga makt, min härlighet till ära!»
Medan ordet ännu var i konungens mun, kom en röst från himmelen: »Dig, konung Nebukadnessar, vare det sagt: Ditt rike har blivit taget ifrån dig;
du skall bliva utstött från människorna och nödgas bo ibland markens djur och äta gräs såsom en oxe; och sju tider skola så gå fram över dig, till dess du besinnar att den Högste råder över människors riken och giver dem åt vem han vill.»
I samma stund gick det ordet i fullbordan på Nebukadnessar; han blev utstött från människorna och måste äta gräs såsom en oxe, och av himmelens dagg vättes hans kropp, till dess att hans hår växte och blev såsom örnfjädrar, och till dess att hans naglar blevo såsom fågelklor.
Men när tiden var förliden, upplyfte jag, Nebukadnessar, mina ögon till himmelen och fick åter mitt förstånd.
Då lovade jag den Högste, jag prisade och ärade honom som lever evinnerligen, honom vilkens välde är ett evigt välde, och vilkens rike varar från släkte till släkte,
honom mot vilken alla som bo på jorden äro att akta såsom intet, ty han gör vad han vill både med himmelens här och med dem som bo på jorden, och ingen kan stå emot hans hand eller säga till honom: »Vad gör du?»
Så fick jag då på den tiden åter mitt förstånd, och jag fick tillbaka min härlighet och glans, mitt rike till ära; och mina rådsherrar och stormän sökte upp mig.
Och jag blev åter insatt i mitt rike, och ännu större makt blev mig given.
Därför prisar nu jag, Nebukadnessar, och upphöjer och ärar himmelens konung, ty alla hans gärningar äro sanning, och hans vägar äro rätta, och dem som vandra i högmod kan han ödmjuka.
Konung Belsassar gjorde ett stort gästabud för sina tusen stormän och höll dryckeslag med de tusen.
Medan nu Belsassar var under vinets välde, befallde han att man skulle bära fram de kärl av guld och silver, som hans fader Nebukadnessar hade tagit ur templet i Jerusalem; ur dem skulle så konungen och hans stormän, hans gemåler och bihustrur dricka.
Då bar man fram de gyllene kärl som hade blivit tagna ur tempelsalen i Guds hus i Jerusalem; och konungen och hans stormän, hans gemåler och bihustrur drucko ur dem.
Medan de så drucko vin, prisade de sina gudar av guld och silver, av koppar, järn, trä och sten.
Då visade sig i samma stund fingrar såsom av en människohand, vilka mitt emot den stora ljusstaken skrevo på den vitmenade väggen i konungens palats; och konungen såg handen som skrev.
Då vek färgen bort ifrån konungens ansikte, och han uppfylldes av oroliga tankar, så att hans länder skälvde och hans knän slogo emot varandra.
Och konungen ropade med hög röst och befallde att man skulle hämta besvärjarna, kaldéerna ock stjärntydarna.
Och konungen lät säga så till de vise i Babel: »Vemhelst som kan läsa denna skrift och meddela mig dess uttydning, han skall bliva klädd i purpur, och den gyllene kedjan skall hängas om hans hals, och han skall bliva den tredje herren i riket.»
Då kommo alla konungens vise tillstädes, men de kunde icke läsa skriften eller säga konungen dess uttydning.
Då blev konung Belsassar ännu mer förskräckt, och färgen vek bort ifrån hans ansikte, och hans stormän stodo bestörta.
Men när konungens och hans stormäns tal kom för konungamodern, begav hon sig till gästabudssalen; där tog hon till orda och sade: »Må du leva evinnerligen, o konung!
Låt icke oroliga tankar uppfylla dig, och må färgen icke vika bort ifrån ditt ansikte.
I ditt rike finnes en man i vilken heliga gudars ande är.
I din faders dagar befanns han hava insikt och förstånd och vishet, lik gudars vishet; och din fader, konung Nebukadnessar, satte honom till den överste bland spåmännen, besvärjarna, kaldéerna och stjärntydarna; ja, detta gjorde din fader konungen,
eftersom en övermåttan hög ande och klokhet och förstånd och skicklighet att uttyda drömmar och lösa gåtor och reda ut invecklade ting fanns hos denne Daniel, åt vilken konungen hade givit namnet Beltesassar.
Låt därför nu tillkalla Daniel; han skall meddela uttydningen.»
När så Daniel hade blivit hämtad till konungen, talade denne till Daniel och sade: »Du är ju Daniel, en av de judiska fångar som min fader konungen förde hit från Juda?
Jag har hört sägas om dig att gudars ande är i dig, och att du har befunnits hava insikt och förstånd och övermåttan stor vishet.
Nu är det så, att de vise och besvärjarna hava blivit hämtade hit till mig för att läsa denna skrift och säga mig dess uttydning; men de kunna icke meddela mig någon uttydning därpå.
Men om dig har jag hört att du kan giva uttydningar och reda ut invecklade ting.
Om du alltså nu kan läsa skriften och säga mig dess uttydning, så skall du bliva klädd i purpur, och den gyllene kedjan skall hängas om din hals, och du skall bliva den tredje herren i riket.»
Då svarade Daniel och sade till konungen: »Dina gåvor må du själv behålla, och dina skänker må du giva åt en annan; dem förutan skall jag läsa skriften för konungen och säga honom uttydningen:
Åt din fader Nebukadnessar, o konung, gav den högste Guden rike, storhet, ära och härlighet;
och för den storhets skull som han hade givit honom darrade alla folk och stammar och tungomål, i förskräckelse för honom.
Vem han ville dödade han, och vem han ville lät han leva; vem han ville upphöjde han, och vem han ville ödmjukade han.
Men när hans hjärta förhävde sig och hans ande blev stolt och övermodig, då störtades han från sin konungatron, och hans ära togs ifrån honom.
Han blev utstött från människors barn, och hans hjärta blev likt ett djurs, och han måste bo ibland vildåsnor och äta gräs såsom en oxe, och av himmelens dagg vättes hans kropp -- detta till dess han besinnade att den högste Guden råder över människors riken och upphöjer vem han vill till att härska över dem.
Men du, Belsassar, hans son, som har vetat allt detta, har ändå icke ödmjukat ditt hjärta,
utan förhävt dig mot himmelens Herre och låtit bära fram inför dig kärlen från hans hus; och du och dina stormän, dina gemåler och bihustrur haven druckit vin ur dem och du har därunder prisat dina gudar av silver och guld, av koppar, järn, trä och sten, som varken se eller höra eller veta något.
Men den Gud som har i sitt våld din ande och alla dina vägar, honom har du icke ärat.
Därför har nu av honom denna hand blivit sänd och denna skrift blivit tecknad.
Och så lyder den skrift som här är tecknad: Mene mene tekel u-farsin.
Och detta är uttydningen därpå: Mene, det betyder: Gud har räknat ditt rikes dagar och gjort ände på det
Tekel, det betyder: du är vägd på en våg och befunnen för lätt.
Peres, det betyder: ditt rike har blivit styckat och givet åt meder och perser.»
Då befallde Belsassar att man skulle kläda Daniel i purpur, och att den gyllene kedjan skulle hängas om hans hals, och att man skulle utropa om honom att han skulle vara den tredje herren i riket.
Samma natt blev Belsassar, kaldéernas konung, dödad.
Och Darejaves av Medien mottog riket, när han var sextiotvå år gammal.
Darejaves fann för gott att sätta över riket ett hundra tjugu satraper, för att sådana skulle finnas överallt i riket.
Och över dem satte han tre furstar, av vilka Daniel var en; inför dessa skulle satraperna avlägga räkenskap, så att konungen icke lede något men.
Men Daniel gjorde sig bemärkt framför de andra furstarna och satraperna, ty en övermåttan hög ande var i honom, och konungen var betänkt på att sätta honom över hela riket.
Då sökte de andra furstarna och satraperna att finna någon sak mot Daniel i det som angick riket.
Men de kunde icke finna någon sådan sak eller något som var orätt, eftersom han var trogen i sin tjänst; ingen försummelse och intet orätt var att finna hos honom.
Då sade männen: »Vi lära icke finna någon sak mot denne Daniel, om vi icke till äventyrs kunna finna en sådan i hans gudsdyrkan.»
Därefter skyndade furstarna och satraperna in till konungen och sade till honom så: »Må du leva evinnerligen, konung Darejaves!
Alla rikets furstar, landshövdingarna och satraperna, rådsherrarna och ståthållarna hava rådslagit om att en kunglig förordning borde utfärdas och ett förbud stadgas, av det innehåll att vilken som helst som under trettio dagar vänder sig med bön till någon annan, vare sig gud eller människa, än till dig, o konung, han skall kastas i lejongropen.
Så låt nu, o konung, härom utfärda ett förbud och sätta upp en skrivelse, som efter Mediens och Persiens oryggliga lag icke kan återkallas.»
I överensstämmelse härmed lät då konung Darejaves sätta upp en skrivelse och utfärda ett förbud.
Men så snart Daniel hade fått veta att skrivelsen var uppsatt, gick han in i sitt hus, varest han i sin övre sal hade fönster som voro öppna i riktning mot Jerusalem.
Där föll han tre gånger om dagen ned på sina knän och bad och tackade sin Gud, såsom han förut hade plägat göra.
När männen nu skyndade till, funno de Daniel bedjande och åkallande sin Gud.
Därefter gingo de till konungen och frågade honom angående det kungliga förbudet: »Har du icke låtit sätta upp ett förbud, av det innehåll att vilken som helst som under trettio dagar vänder sig med bön till någon annan, vare sig gud eller människa, än till dig, o konung, han skall kastas i lejongropen?»
Konungen svarade och sade: »Jo, och det påbudet står fast efter Mediens och Persiens oryggliga lag.»
Då svarade de och sade till konungen: »Daniel, en av de judiska fångarna, aktar varken på dig eller på det förbud som du har låtit sätta upp, utan förrättar sin bön tre gånger om dagen.»
När konungen hörde detta, blev han mycket bedrövad och gjorde sig bekymmer över huru han skulle kunna rädda Daniel; ända till solnedgången mödade han sig med att söka en utväg att hjälpa honom.
Då skyndade männen till konungen och sade till honom: »Vet, o konung, att det är en Mediens och Persiens lag att intet förbud och ingen förordning som konungen utfärdar kan återkallas.»
Då lät konungen hämta Daniel och kasta honom i lejongropen och konungen talade till Daniel och sade: »Din Gud, den som du så oavlåtligen dyrkar, han må rädda dig.»
Och man förde fram en sten och lade den över gropens öppning, och konungen förseglade den med sitt eget och med sina stormäns signet, för att ingen förändring skulle kunna göras i det som nu hade skett med Daniel.
Därefter gick konungen hem till sitt palats och tillbragte hela natten under fasta och lät inga kvinnor komma inför sig; och sömnen flydde honom.
Sedan om morgonen, när det dagades, stod konungen upp och gick med hast till lejongropen.
Och när han hade kommit nära intill gropen, ropade han på Daniel med ängslig röst; konungen talade till Daniel och sade: »Daniel, du den levande Gudens tjänare, har väl din Gud, den som du så oavlåtligen dyrkar, kunnat rädda dig från lejonen?»
Då svarade Daniel konungen: »Må du leva evinnerligen, o konung!
Min Gud har sänt sin ängel och tillslutit lejonens gap, så att de icke hava gjort mig någon skada.
Ty jag har inför honom befunnits oskyldig; ej heller har jag förbrutit mig mot dig, o konung.
Då blev konungen mycket glad, och befallde att man skulle taga Daniel upp ur gropen.
Och när Daniel hade blivit tagen upp ur gropen, kunde man icke upptäcka någon skada på honom; ty han hade trott på sin Gud.
Sedan lät konungen hämta de män som hade anklagat Daniel, och han lät kasta dem i lejongropen, med deras barn och hustrur; och innan de ännu hade hunnit till bottnen i gropen, föllo lejonen över dem och krossade alla deras ben.
Därefter lät konung Darejaves skriva till alla folk och stammar och tungomål som funnos på hela jorden: »Mycken frid vare med eder!
Härmed giver jag befallning att man inom mitt rikes hela område skall bäva och frukta för Daniels Gud.
Ty han är den levande Guden, som förbliver evinnerligen; och hans rike är sådant att det icke kan förstöras, och hans välde består intill änden.
Han är en räddare och hjälpare, och han gör tecken och under i himmelen och på jorden, han som har räddat Daniel ur lejonens våld.»
Och denne Daniel steg i ära och makt under Darejaves' och under persern Kores' regeringar.
I den babyloniske konungen Belsassars första regeringsår hade Daniel en dröm och såg en syn på sitt läger.
Sedan tecknade han upp drömmen och meddelade huvudsumman av dess innehåll.
Detta är Daniels berättelse: Jag hade en syn om natten, och såg i den huru himmelens fyra vindar stormade fram mot det stora havet.
Och fyra stora djur stego upp ur havet, det ena icke likt det andra.
Det första liknade ett lejon, men det hade vingar såsom en örn.
Medan jag ännu såg härpå, rycktes vingarna av djuret, och det restes upp från jorden, så att det blev ställt på två fötter såsom en människa, och ett mänskligt hjärta blev givet åt det.
Sedan fick jag se ännu ett djur, det andra i ordningen; det var likt en björn, och det reste upp sin ena sida, och det hade tre revben i sitt gap, mellan tänderna.
Och till det djuret blev så sagt: »Stå upp och sluka mycket kött.»
Därefter fick jag se ett annat djur, som liknade en panter, men på sina sidor hade det fyra fågelvingar; och djuret hade fyra huvuden, och välde blev givet åt det.
Därefter fick jag i min syn om natten se ett fjärde djur, övermåttan förskräckligt, fruktansvärt och starkt; det hade stora tänder av järn, det uppslukade och krossade, och vad som blev kvar trampade det under fötterna; det var olikt alla de förra djuren och hade tio horn.
Men under det att jag betraktade hornen, fick jag se huru mellan dem ett annat horn sköt upp, ett litet, för vilket tre av de förra hornen blevo bortstötta; och se, det hornet hade ögon lika människoögon, och en mun som talade stora ord.
Medan jag ännu såg härpå, blevo troner framsatta, och en som var gammal satte sig ned.
Hans klädnad var snövit, och håret på hans huvud var såsom ren ull; hans tron var av eldslågor, och hjulen därpå voro av flammande eld.
En flod av eld strömmade ut från honom, tusen gånger tusen voro hans tjänare, och tio tusen gånger tio tusen stodo där till hans tjänst.
Så satte man sig ned till doms, och böcker blevo upplåtna.
Medan jag nu såg härpå, skedde det att, för de stora ords skull som hornet talade -- medan jag ännu såg härpå -- djuret dödades och dess kropp förstördes och kastades i elden för att brännas upp.
Från de övriga djuren togs ock deras välde, ty deras livslängd var bestämd till tid och stund.
Sedan fick jag, i min syn om natten, se huru en som liknade en människoson kom med himmelens skyar; och han nalkades den gamle och fördes fram inför honom.
Åt denne gavs välde och ära och rike, och alla folk och stammar och tungomål måste tjäna honom.
Hans välde är ett evigt välde, som icke skall tagas ifrån honom, och hans rike skall icke förstöras.
Då kände jag, Daniel, min ande oroas i sin boning, och den syn som jag hade haft förskräckte mig.
Jag gick fram till en av dem som stodo där och bad honom om en tillförlitlig förklaring på allt detta Och han svarade mig och sade mig uttydningen därpå:
»De fyra stora djuren betyda att fyra konungar skola uppstå på jorden.
Men sedan skola den Högstes heliga undfå riket och taga det i besittning för evig tid, ja, för evigheters evighet.»
Därefter ville jag hava tillförlitlig förklaring angående det fjärde djuret, som var olikt alla de andra, det som var så övermåttan förskräckligt och hade tänder av järn och klor av koppar, det som uppslukade och krossade och sedan trampade under fötterna vad som blev kvar;
så ock angående de tio hornen på dess huvud, och angående det nya hornet, det som sedan sköt upp, och för vilket tre andra föllo av, det hornet som hade Ögon, och en mun som talade stora ord, det som var större att skåda än de övriga,
det hornet som jag ock hade sett; föra krig mot de heliga och bliva dem övermäktigt,
till dess att den gamle kom och rätt blev skipad åt den Högstes heliga och tiden var inne, då de heliga fingo taga riket i besittning.
Då svarade han så: »Det fjärde djuret betyder att ett fjärde rike skall uppstå på jorden, ett som är olikt alla de andra rikena.
Det skall uppsluka hela jorden och förtrampa och krossa den.
Och de tio hornen betyda att tio konungar skola uppstå i det riket; och efter dem skall uppstå en annan, som skall vara olik de förra, och som skall slå ned tre konungar.
Och denne skall upphäva sitt tal mot den Högste och föröda den Högstes heliga; han skall sätta sig i sinnet att förändra heliga tider och lagar; och de skola givas i hans hand under en tid, och tider, och en halv tid.
Men dom skall bliva hållen, och hans välde skall tagas ifrån honom och fördärvas och förgöras i grund.
Men rike och välde och storhet, utöver alla riken under himmelen, skall givas åt den Högstes heligas folk.
Dess rike skall vara ett evigt rike, och alla välden skola tjäna och lyda det.»
Här slutar berättelsen.
Men jag, Daniel, uppfylldes av många oroliga tankar, och färgen vek bort ifrån mitt ansikte; men jag bevarade i mitt hjärta vad som hade hänt.
I konung Belsassars tredje regeringsår såg jag, Daniel, en syn, en som kom efter den jag förut hade sett.
Då jag nu i denna syn såg till, tyckte jag mig vara i Susans borg i hövdingdömet Elam; och då jag vidare såg till i synen, fann jag mig vara vid floden Ulai.
Och när jag lyfte upp mina ögon, fick jag se en vädur stå framför floden, och han hade två horn; och båda hornen voro höga, men det ena var högre än det andra, och detta som var högre sköt sist upp.
Jag såg väduren stöta med hornen västerut och norrut och söderut, och intet djur kunde stå honom emot, och ingen kunde rädda ur hans våld; han for fram såsom han ville och företog sig stora ting.
Och när jag vidare gav akt, fick jag se en bock komma västerifrån och gå fram över hela jorden, dock utan att röra vid jorden; och bocken hade ett ansenligt horn i pannan.
Och han nalkades väduren med de båda hornen, den som jag hade sett stå framför floden, och sprang emot honom i väldig vrede.
Jag såg honom komma ända inpå väduren och störta över honom i förbittring, och han stötte till väduren och krossade hans båda horn, så att väduren icke hade någon kraft att stå emot honom.
Sedan slog han honom till jorden och trampade på honom; och ingen fanns, som kunde rädda väduren ur hans våld.
Och bocken företog sig mycket stora ting.
Men när han hade blivit som starkast, brast det stora hornet sönder, och fyra andra ansenliga horn sköto upp i dess ställe, åt himmelens fyra väderstreck.
Och från ett av dem gick ut ett nytt horn, i begynnelsen litet, och det växte övermåttan söderut och österut och åt »det härliga landet» till.
Och det växte ända upp till himmelens härskara och kastade några av denna härskara, av stjärnorna, ned till jorden och trampade på dem.
Ja, till och med mot härskarornas furste företog han sig stora ting: han tog bort ifrån honom det dagliga offret, och hans helgedoms boning slogs ned.
Jämte det dagliga offret bliver ock en härskara prisgiven, för överträdelses skull.
Och det slår sanningen ned till jorden och lyckas väl i vad det företager sig.
Sedan hörde jag en av de heliga tala, och en annan helig frågade denne som talade: »Huru lång tid avser synen om det dagliga offret, och om överträdelsen som kommer åstad förödelse, och om förtrampandet av både helgedom och härskara?»
Då svarade han mig: »Två tusen tre hundra aftnar och morgnar; därefter skall helgedomen komma till sin rätt igen.»
När nu jag, Daniel, hade sett denna syn och sökte att förstå den, fick jag se en som såg ut såsom en man stå framför mig.
Och mitt över Ulai hörde jag rösten av en människa som ropade och sade: »Gabriel, uttyd synen för denne.»
Då kom han intill platsen där jag stod, men jag blev förskräckt, när han kom, och föll ned på mitt ansikte.
Och han sade till mig: »Giv akt härpå, du människobarn; ty synen syftar på ändens tid.»
Medan han så talade med mig, låg jag i vanmakt, med mitt ansikte mot jorden; men han rörde vid mig och reste upp mig igen.
Därefter sade han: »Se, jag vill kungöra för dig vad som skall ske, när det lider mot slutet med vreden ty på ändens tid syftar detta.
Väduren som du såg, han med de två hornen, betyder Mediens och Persiens konungar.
Men bocken är Javans konung, och det stora hornet i hans panna är den förste konungen.
Men att det brast sönder, och att fyra andra uppstodo i dess ställe, det betyder att fyra riken skola uppstå av hans folk, dock icke jämlika med honom i kraft.
Och vid slutet av deras välde, när överträdarna hava fyllt sitt mått, skall en fräck och arglistig konung uppstå;
han skall bliva stor i kraft, dock icke jämlik med den förre i kraft och han skall komma åstad så stort fördärv att man måste förundra sig; och han skall lyckas väl och få fullborda sitt uppsåt.
Ja, han skall fördärva många, och jämväl de heligas folk.
Därigenom att han är så klok, skall han lyckas så väl med sitt svek, han skall föresätta sig stora ting, oförtänkt skall han fördärva många.
Ja, mot furstarnas furste skall han sätta sig upp; men utan människohand skall han då varda krossad.
Och synen angående aftnarna och morgnarna, varom nu är talat, är sanning.
Men göm du den synen, ty den syftar på en avlägsen framtid.»
Men jag, Daniel, blev maktlös och låg sjuk en tid.
Sedan stod jag upp och förrättade min tjänst hos konungen; och jag var häpen över synen, men ingen förstod den.
I Darejaves', Ahasveros' sons, första regeringsår -- hans som var av medisk släkt, men som hade blivit upphöjd till konung över kaldéernas rike --
i dennes första regeringsår kom jag, Daniel, att i skrifterna lägga märke till det antal år, som HERREN hade angivit för profeten Jeremia, när han sade att han ville låta sjuttio år gå till ända, medan Jerusalem låg öde.
Då vände jag mitt ansikte till Herren Gud med ivrig bön och åkallan, och fastade därvid i säck och aska.
Jag bad till HERREN, min Gud, och bekände och sade: »Ack Herre, du store och fruktansvärde Gud, du som håller förbund och bevarar nåd mot dem som älska dig och hålla dina bud!
Vi hava syndat och gjort illa och varit ogudaktiga och avfälliga; vi hava vikit av ifrån dina bud och rätter.
Vi hava icke hörsammat dina tjänare profeterna, som talade i ditt namn till våra konungar, furstar och fader och till allt folket i landet.
Du, Herre, är rättfärdig, men vi måste blygas, såsom vi ock nu göra, vi Juda man och Jerusalems invånare, ja, hela Israel, både de som bo nära och de som bo fjärran i alla andra länder dit du har fördrivit dem, därför att de voro otrogna mot dig.
Ja, Herre, vi med våra konungar, furstar och fäder måste blygas, därför att vi hava syndat mot dig.
Men hos Herren, vår Gud, är barmhärtighet och förlåtelse.
Ty vi voro avfälliga från
och hörde icke HERRENS, vår Guds, röst, så att vi vandrade efter hans lagar, dem som han förelade oss genom sina tjänare profeterna.
Nej, hela Israel överträdde din lag och vek av, utan att höra din röst.
Därför utgöt sig ock över oss den förbannelse som han hade svurit att sända, och som står skriven i Moses, Guds tjänares, lag; ty vi hade ju syndat mot honom.
Han höll sina ord, vad han hade talat mot oss, och mot domarna som dömde oss; och han lät en så stor olycka komma över oss, att ingenstädes under himmelen något sådant har skett, som det som nu har skett i Jerusalem.
I enlighet med vad som står skrivet i Moses lag kom all denna olycka över oss, men ändå sökte vi icke att blidka HERREN, vår Gud, genom att omvända oss från våra missgärningar och akta på din sanning.
Därför vakade ock HERREN över att olyckan drabbade oss; ty HERREN, vår Gud, är rättfärdig i alla de gärningar som han gör, men hörde icke hans röst.
Och nu, Herre, vår Gud, du som förde ditt folk ut ur Egyptens land med stark hand, och så gjorde dig ett namn, som är detsamma än i dag!
Vi hava syndat, vi hava varit ogudaktiga.
Men Herre, låt, för all din rättfärdighets skull, din vrede och förtörnelse vända sig ifrån din stad Jerusalem, ditt heliga berg; ty genom våra synder och genom våra faders missgärningar hava Jerusalem och ditt folk blivit till smälek för alla som bo omkring oss.
Och hör nu, du vår Gud, din tjänares bön och åkallan, och låt ditt ansikte lysa över din ödelagda helgedom, för Herrens skull.
Böj, min Gud, ditt öra härtill och hör; öppna dina ögon och se vilken förödelse som har övergått oss, och se till staden som är uppkallad efter ditt namn.
Ty icke i förlitande på vad rättfärdigt vi hava gjort bönfalla vi inför dig, utan i förlitande på din stora barmhärtighet.
O Herre, hör, o Herre, förlåt; o Herre, akta härpå, och utför ditt verk utan att dröja -- för din egen skull, min Gud, ty din stad och ditt folk äro uppkallade efter ditt namn.»
Medan jag ännu så talade och bad och bekände min egen och mitt folk Israels synd och inför HERREN, min Gud, frambar min förbön för min Guds heliga berg --
medan jag alltså ännu så talade i min bön, kom Gabriel till mig i flygande hast, den man som jag förut hade sett i min syn; och det var vid tiden för aftonoffret.
Han undervisade mig och talade till mig och sade: »Daniel, jag har nu begivit mig hit för att lära dig förstånd.
Redan när du begynte din bön, utgick befallning, och jag har kommit för att giva dig besked, ty du är högt benådad.
Så giv nu akt på ordet, och akta på synen.
Sjuttio veckor äro bestämda över ditt folk och över din heliga stad, innan en gräns sättes för överträdelsen och synderna få en ände och missgärningen varder försonad och en evig rättfärdighet framhavd, och innan syn och profetia beseglas och en höghelig helgedom bliver smord.
Så vet nu och förstå: Från den tid då ordet om att Jerusalem åter skulle byggas upp utgick, till dess en smord, en furste, kommer, skola sju veckor förgå; och under sextiotvå veckor skall det åter byggas upp med sina gator och sina vallgravar, om ock i tider av trångmål.
Men efter de sextiotvå veckorna skall en som är smord förgöras, utan att någon efterföljer honom.
Och staden och helgedomen skall en anryckande furstes folk förstöra; men själv skall denne få sin ände i störtfloden.
Och intill änden skall strid vara; förödelse är oryggligt besluten.
Och han skall med många sluta ett starkt förbund för en vecka, och för en halv vecka skola genom honom slaktoffer och spisoffer vara avskaffade; och på styggelsens vinge skall förödaren komma.
Detta skall fortgå, till dess att förstöring och oryggligt besluten straffdom utgjuter sig över förödaren.»
I den persiske konungen Kores' tredje regeringsår fick Daniel, som ock kallades Beltesassar, en uppenbarelse; den uppenbarelsen är sanning och bådar stor vedermöda.
Och han aktade på uppenbarelsen och lade märke till synen.
Jag, Daniel, hade då gått sörjande tre veckors tid.
Jag åt ingen smaklig mat, kött och vin kommo icke i min mun, ej heller smorde jag min kropp med olja, förrän de tre veckorna hade gått till ända.
På tjugufjärde dagen i första månaden, när jag var vid stranden av den stora floden, nämligen Hiddekel,
fick jag, då jag lyfte upp mina ögon, se en man stå där, klädd i linnekläder och omgjordad kring sina länder med ett bälte av guld från Ufas.
Hans kropp var såsom av krysolit hans ansikte liknade en ljungeld hans ögon voro såsom eldbloss, han armar och fötter såsom glänsande koppar; och ljudet av hans tal var såsom ett väldigt dån.
Och jag, Daniel, var den ende som såg synen; de män som voro med mig sågo den icke, men en stor förskräckelse föll över dem, så att de flydde bort och gömde sig.
Så blev jag allena kvar, och när jag såg den stora synen, förgick all min kraft; färgen vek bort ifrån mitt ansikte, så att det blev dödsblekt, och jag hade ingen kraft mer kvar.
Då hörde jag ljudet av hans tal; och på samma gång jag hörde ljudet av hans tal, där jag låg i vanmakt på mitt ansikte, med ansiktet mot jorden,
rörde en hand vid mig och hjälpte mig, så att jag skälvande kunde resa mig på mina knän och händer.
Sedan sade han till mig: »Daniel, du högt benådade man, giv akt på de ord som jag vill tala till dig, och res dig upp på dina fötter; ty jag har nu blivit sänd till dig.»
När han så talade till mig, reste jag mig bävande upp.
Och han sade till mig: »Frukta icke, Daniel, ty redan ifrån första dagen, då när du vände ditt hjärta till att söka förstånd och till att ödmjuka dig inför din Gud, hava dina ord varit hörda; och jag har nu kommit för dina ords skull.
Fursten för Persiens rike stod mig emot under tjuguen dagar; men då kom Mikael, en av de förnämsta furstarna, mig till hjälp, under det att jag förut hade stått där allena mot Persiens konungar.
Och nu har jag kommit för att undervisa dig om vad som skall hända ditt folk i kommande dagar; ty också detta är en syn som syftar på framtiden.»
Under det han så talade till mig, böjde jag mitt ansikte mot jorden och var stum.
Men se, han som var lik en människa rörde vid mina läppar.
Då upplät jag min mun och talade och sade till honom som stod framför mig: »Min herre, vid den syn jag såg har jag känt mig gripen av vånda, och jag har ingen kraft mer kvar.
Huru skulle också min herres tjänare, en sådan som jag, kunna tala med en sådan som min herre är?
Jag har nu ingen kraft mer i mig och förmår icke mer att andas.»
Då rörde han som såg ut såsom en människa åter vid mig och styrkte mig.
Han sade: »Frukta icke, du högt benådade man; frid vare med dig, var stark, ja, var stark.»
När han så talade med mig, kände jag mig styrkt och sade: »Tala, min herre, ty du har nu styrkt mig.»
Då sade han: »Kan du nu förstå varför jag har kommit till dig?
Men jag måste strax vända tillbaka för att strida mot fursten för Persien, och när jag är fri ifrån honom, kommer fursten för Javan.
Dock vill jag förkunna för dig vad som är upptecknat i sanningens bok.
Och ingen enda står mig bi mot dessa, förutom Mikael, eder furste.
Och jag stod vid hans sida såsom hans stöd och värn i medern Darejaves' första regeringsår.
Och nu skall jag förkunna för dig vad visst är.
Se, ännu tre konungar skola uppstå i Persien, och den fjärde skall förvärva sig större rikedomar än någon av de andra, och när han har blivit som starkast genom sina rikedomar, skall han uppbjuda all sin makt mot Javans rike.
Sedan skall en väldig konung uppstå, och han skall härska med stor makt och göra vad han vill.
Men knappt har han uppstått, så skall hans rike brista sönder och bliva delat efter himmelens förra väderstreck; och det skall icke tillfalla hans avkomlingar eller förbliva lika mäktigt som när han hade makten; ty hans rike skall omstörtas och tillfalla andra än dem.
Och konungen i Söderlandet skall bliva mäktig, så ock en av hans furstar; ja, denne skall bliva en ännu mäktigare härskare än han själv, och hans herradöme skall bliva stort.
Och efter några år skola de förbinda sig med varandra, och Söderlandskonungens dotter skall draga till konungen i Nordlandet för att komma åstad förlikning.
Men hon skall icke kunna behålla den makt hon vinner, ej heller skall han och hans makt bliva beståndande; utan hon skall bliva given till pris, hon jämte dem som läto henne draga dit, både hennes fader och den man som i sin tid tog henne till sig.
Men av telningarna från hennes rot skall en stiga upp på hans plats; denne skall draga mot Nordlandskonungens här och tränga in i hans fäste och göra med folket vad han vill och behålla övermakten.
Deras gudar och beläten och deras dyrbara håvor, både silver och guld, skall han ock föra såsom byte till Egypten.
Sedan skall han i några år lämna Nordlandskonungen i ro.
Däremot skall denne tränga in i Söderlandskonungens rike, men han skall få vända tillbaka till sitt land igen.
Och hans söner skola rusta sig till strid och samla en väldig krigs här; och den skall rycka fram och svämma över och utbreda sig; och den skall komma igen, och striden skall föras ända fram till hans fäste.
Då skall konungen i Söderlandet resa sig i förbittring och draga ut och strida mot konungen i Nordlandet; och denne skall ställa upp en stor härskara, men den härskaran skall varda given i den andres hand.
När då härskaran är sin kos, växer hans övermod; men om han än han slagit ned tiotusenden, får han dock icke makten.
Konungen i Nordlandet skall ställa upp en ny härskara, större än den förra; och efter en tid av några år skall han komma med en stor krigshär och stora förråd.
Vid samma tid skola många andra resa sig mot konungen i Söderlandet; våldsmän av ditt eget folk skola ock upphäva sig, för att synen skall fullbordas; men dessa skola falla.
Och konungen i Nordlandet skall rycka an och kasta upp vallar och intaga en välbefäst stad; och Söderlandets makt skall icke kunna hålla stånd, dess utvalda krigsfolk skall icke hava någon kraft till motstånd.
Och han som rycker emot honom skall göra vad han vill, och ingen skall kunna stå emot honom; han skall sätta sig fast i »det härliga landet», och förstöring skall komma genom hans hand.
Han skall rycka an med hela sitt rikes makt; dock är han hågad för förlikning, och en sådan skall han komma åstad.
En av sina döttrar skall han giva åt honom till hustru, henne till fördärv.
Men detta skall icke hava något bestånd och icke vara honom till gagn.
Därefter skall han vända sig mot öländerna och intaga många; men en härförare skall göra slut på hans smädelser, ja, låta hans smädelser vända tillbaka över honom själv.
Då skall han vända sig till sitt eget lands fästen; men han skall vackla och falla och sedan icke mer finnas till.
Och på hans plats skall uppstå en annan, en som låter en fogde draga igenom det land som är hans rikes prydnad; men efter några dagar skall han störtas, dock icke genom vrede, ej heller i krig.
Och på hans plats skall uppstå en föraktlig man, åt vilken konungavärdighet icke var ämnad; oförtänkt skall han komma och bemäktiga sig riket genom ränker.
Och översvämmande härar skola svämmas bort för honom och krossas, så ock förbundets furste.
Från den stund då man förbinder sig med honom skall han bedriva svek.
Han skall draga åstad och få övermakten, med allenast litet folk.
Oförtänkt skall han falla in i landets bördigaste trakter, och skall göra ting som hans fäder och hans fäders fäder icke hade gjort; byte och rov och gods skall han strö ut åt sitt folk; och mot fästena skall han förehava anslag, intill en viss tid.
Och han skall uppbjuda sin kraft; och sitt mod emot konungen i Söderlandet och komma med en stor här, men konungen i Söderlandet skall ock rusta sig till strid, med en mycket stor och talrik här; dock skall han icke kunna hålla stånd, för de anslags skull som göras mot honom.
De som äta hans bröd skola störta honom.
Och hans här skall svämma över, och många skola bliva slagna och falla.
Båda konungarna skola hava ont i sinnet, där de sitta tillhopa vid samma bord, skola de tala lögn, men det skall icke hava någon framgång; ty ännu dröjer änden, intill den bestämda tiden.
Han skall vända tillbaka till sitt land med stora förråd, och han skall lägga planer mot det heliga förbundet; och när han har fullbordat dem, skall han vända tillbaka till sitt land.
På bestämd tid skall han sedan åter draga åstad mot Söderlandet, men denna senare gång skall det ej gå såsom den förra.
Ty skepp från Kittim skola komma emot honom, och han skall förlora modet.
Då skall han vända om och rikta sin vrede mot det heliga förbundet och giva den fritt lopp.
Och när han har kommit hem, skall han lyssna till dem som hava övergivit det heliga förbundet.
Och härar, utsända av honom, skola komma och oskära helgedomens fäste och avskaffa det dagliga offret och ställa upp förödelsens styggelse.
Och dem som hava kränkt förbundet skall han med hala ord locka till helt avfall; men de av folket, som känna sin Gud, skola stå fasta och hålla ut.
Och de förståndiga bland folket skola lära många insikt; men de skola bliva hemsökta med svärd och eld, med fångenskap och plundring, till en tid;
dock skall under hemsökelsen en liten seger beskäras dem, och många skola då av skrymteri sluta sig till dem.
Hemsökelsen skall träffa somliga av de förståndiga, för att en luttring skall ske bland dem, så att de varda renade och tvagna till ändens tid; ty ännu dröjer denna, intill den bestämda tiden.
Och konungen skall göra vad han vill och skall förhäva sig och uppträda stormodigt mot allt vad gud heter; ja, mot gudars Gud skall han tala sådant att man måste förundra sig.
Och allt skall lyckas honom väl, till dess att vredens tid är ute, då när det har skett, som är oryggligt beslutet.
På sina fäders gudar skall han icke akta, ej heller skall han akta på den som är kvinnors lust eller på någon annan Gud, utan han skall uppträda stormodigt mot dem alla.
Men fästenas gud skall han i stället ära; en gud som hans fäder icke hava känt skall han ära med guld och silver och ädla stenar och andra dyrbara ting.
Och mot starka fästen skall han med en främmande guds hjälp göra vad honom lyster; dem som erkänna denne skall han bevisa stor ära, han skall sätta dem att råda över många, och han skall utskifta jord åt dem till belöning.
Men på ändens tid skall konungen i Söderlandet drabba samman med honom; och konungen i Nordlandet skall storma fram mot denne med vagnar och ryttare och många skepp, och skall falla in i främmande länder och svämma över och utbreda sig.
Han skall ock falla in i »det härliga landet», och många andra länder skola bliva hemsökta; men dessa skola komma undan hans hand: Edom och Moab och huvuddelen av Ammons barn.
Ja, han skall uträcka sin hand mot främmande länder, och Egyptens land skall icke slippa undan;
han skall bemäktiga sig skatter av guld och silver och allahanda dyrbara ting i Egypten; och libyer och etiopier skola följa honom åt.
Då skall han från öster och norr få höra rykten som förskräcka honom; och kan skall draga ut i stor vrede för att förgöra många och giva dem till spillo.
Och sina palatstält skall han slå upp mellan havet och helgedomens härliga berg.
Men han går till sin undergång, och ingen skall finnas, som hjälper honom.»
På den tiden skall Mikael träda upp, den store fursten som står såsom försvarare för dina landsmän; och då kommer en tid av nöd, vars like icke har funnits, allt ifrån den dag då människor blevo till och ända till den tiden.
Men på den tiden skola av ditt folk alla de varda frälsta, som finnas skrivna i boken.
Och många av dem som sova i mullen skola uppvakna, somliga till evigt liv, och somliga till smälek och evig blygd.
De förståndiga skola då lysa, såsom fästet lyser, och de som hava fört de många till rättfärdighet såsom stjärnor, alltid och evinnerligen.
Men du, Daniel, må gömma dessa ord och försegla denna skrift intill ändens tid; många komma att rannsaka den, och insikten skall så växa till.»
När nu jag, Daniel, såg till, fick jag se två andra stå där, en på flodens ena strand, och en på dess andra strand.
Och en av dem sade till mannen som var klädd i linnekläder, och som stod ovanför flodens vatten: »Huru länge dröjer det, innan änden kommer med dessa förunderliga ting?»
Och jag hörde på mannen som var klädd i linnekläder, och som stod ovanför flodens vatten, och han lyfte sin högra hand och sin vänstra hand upp mot himmelen och svor vid honom som lever evinnerligen att efter en tid, och tider, och en halv tid, och när det heliga folkets makt hade blivit krossad i grund, då skulle allt detta varda fullbordat.
Och jag hörde detta, men förstod det icke; och jag frågade: »Min herre, vad bliver slutet på allt detta?»
Då sade han: »Gå, Daniel, ty dessa ord skola förbliva gömda och förseglade intill ändens tid.
Många skola varda renade och tvagna och luttrade, men de ogudaktiga skola öva sin ogudaktighet, och ingen ogudaktig skall förstå detta; men de förståndiga skola förstå det.
Och från den tid då det dagliga offret bliver avskaffat och förödelsens styggelse uppställd skola ett tusen två hundra nittio dagar förgå.
Säll är den som förbidar och hinner fram till ett tusen tre hundra trettiofem dagar.
Men gå du åstad mot ändens tid; sedan du har vilat, skall du uppstå till din del, vid dagarnas ände.»
Detta är HERRENS ord som kom till Hosea, Beeris son, i Ussias, Jotams, Ahas' och Hiskias, Juda konungars, tid, och i Jerobeams, Joas' sons, Israels konungs, tid.
När HERREN först begynte tala genom Hosea, sade HERREN till honom: »Gå åstad och skaffa dig en trolös hustru och barn -- av en trolös moder; ty i trolös avfällighet löper landet bort ifrån HERREN.
Då gick han åstad och tog Gomer, Diblaims dotter; och hon blev havande och födde honom en son.
Och HERREN sade till honom: »Giv denne namnet Jisreel; ty när ännu en liten tid har förgått, skall jag hemsöka Jisreels blodskulder på Jehus hus och göra slut på konungadömet i Israels hus.
Och det skall ske på den dagen att jag skall bryta sönder Israels båge i Jisreels dal.»
Och hon blev åter havande och födde en dotter.
Då sade han till honom: »Giv denna namnet Lo-Ruhama; ty jag vill icke vidare förbarma mig över Israels hus, så att jag förlåter dem.
Men över Juda hus vill jag förbarma mig, och jag skall giva dem frälsning genom HERREN, deras Gud; icke genom båge och svärd och vad till kriget hör skall jag frälsa dem, icke genom hästar och ryttare.
Och när hon hade avvant Lo-Ruhama, blev hon åter havande och födde en son.
Då sade han: »Giv denne namnet Lo-Ammi; ty I ären icke mitt folk, ej heller vill jag höra eder till.»
Men antalet av Israels barn skall bliva såsom havets sand, som man icke kan mäta, ej heller räkna; och det skall ske, att i stället för att det sades till dem: »I ären icke mitt folk», skola de kallas »den levande Gudens barn».
Och Juda barn och Israels barn skola samla sig tillhopa, och skola sätta över sig ett gemensamt huvud, och skola draga upp ur landet; ty stor skall Jisreels dag vara.
Kallen då edra bröder Ammi och edra systrar Ruhama.
Gån till rätta med eder moder, gån till rätta; ty hon är icke min hustru, och jag är icke hennes man.
Må hon skaffa bort det lösaktiga väsendet från sitt ansikte och otuktsväsendet från sin barm.
Varom icke, skall jag kläda av henne, så att hon ligger naken, jag skall låta henne stå där sådan hon var den dag då hon föddes.
Jag skall göra henne lik en öken och låta henne bliva såsom ett torrt land och låta henne dö av törst.
Och mot hennes barn skall jag icke visa något förbarmande, eftersom de äro barn av en trolös moder;
ty deras moder var en trolös kvinna, ja, hon som födde dem bedrev skamliga ting.
Hon sade ju: »Jag vill följa efter mina älskare, som giva mig min mat och min dryck, min ull och mitt lin, min olja och mitt vin.»
Se, därför skall jag nu ock stänga din väg med törnen.
Ja, en mur skall jag resa framför henne, så att hon ej skall finna någon stig.
När hon då löper efter sina älskare, skall hon icke få dem fatt; när hon söker dem, skall hon ej finna dem.
Då skall hon säga: »Jag vill gå tillbaka till min förste man ty bättre var mig då än nu.»
Men hon har icke förstått att det var jag som skänkte åt henne både säden och vinet och oljan, och att det var jag som gav henne så mycket silver, så ock guld, varav de gjorde sin Baalsbild.
Därför skall jag taga tillbaka min säd, när tiden är inne, och mitt vin, när stunden kommer; jag skall taga bort min ull och mitt lin, det varmed hon skulle skyla sin blygd.
Ja, nu skall jag blotta hennes skam inför hennes älskares ögon, och ingen skall rädda henne ur min hand.
Och jag skall göra slut på all hennes fröjd, på hennes fester, nymånader och sabbater och på alla hennes högtider.
Jag skall föröda hennes vinträd och fikonträd, dem om vilka hon sade: »De äro en lön som mina älskare hava givit mig.» och jag skall göra därav en vildmark, och markens djur skola äta därav.
Så skall jag hemsöka henne för hennes Baalsdagar, då hon tände offereld åt Baalerna och prydde sig med ring och bröstspänne och följde efter sina älskare, men glömde mig, säger HERREN.
Se, fördenskull vill jag locka henne bort och föra henne ut i öknen och tala ljuvligt till henne.
Därefter skall jag giva henne tillbaka hennes vingårdar och göra Akors dal till en hoppets port.
Då skall hon sjunga såsom i sin ungdoms dagar, och såsom på den dag då hon drog upp ur Egyptens land.
Och det skall ske på den dagen, säger HERREN, att du skall ropa: »Min man!», och icke mer ropa till mig: »Min Baal!»
Ja, Baalernas namn skall jag skaffa bort ur hennes mun, så att de icke mer skola nämnas vid namn.
Och jag skall på den dagen för deras räkning sluta ett förbund med djuren på marken och med fåglarna under himmelen och med kräldjuren på jorden.
Och båge och svärd och vad till kriget hör skall jag bryta sönder och skaffa bort ur landet och låta dem bo där i trygghet.
Och jag skall trolova mig med dig för evig tid; jag skall trolova mig med dig rättfärdighet och rätt, i nåd och barmhärtighet.
Ja, i trofasthet skall jag trolova mig med dig, och du skall så lära känna HERREN.
Och det skall ske på den dagen att jag skall bönhöra, säger HERREN, jag skall bönhöra himmelen, och den skall bönhöra jorden,
och jorden skall bönhöra säden, så ock vinet och oljan, och de skola bönhöra Jisreel.
Och jag skall plantera henne åt mig i landet och förbarma mig över Lo-Ruhama och säga till Lo-Ammi: »Du är mitt folk.»
Och det skall svara: »Du är min Gud.»
Och HERREN sade till mig: »Gå ännu en gång åstad och giv din kärlek åt en kvinna som har en älskare och är en äktenskapsbryterska; likasom HERREN älskar Israels barn, fastän de vända sig till andra gudar och älska druvkakor.»
Och jag köpte henne åt mig och gav för henne femton siklar silver och en homer korn, och därutöver en letek korn.
Sedan sade jag till henne: »I lång tid skall du bliva sittande för min räkning, utan att få bedriva någon otukt, och utan att hava att skaffa med någon man; och jag skall bete mig sammalunda mot dig.
Ja, i lång tid skola Israels barn få sitta utan konung och furste, utan offer och stoder och utan efod och husgudar.
Sedan skola Israels barn omvända sig och söka HERREN, sin Gud, och David, sin konung; med fruktan skola de söka HERREN och hans goda, i kommande dagar.
Hören HERRENS ord, I Israels barn.
Ty HERREN har sak med landets inbyggare, eftersom ingen sanning och ingen kärlek och ingen Guds kunskap finnes i landet.
Man svär och ljuger, man mördar och stjäl och begår äktenskapsbrott; man far fram på våldsverkares vis, och blodsdåd följer på blodsdåd.
Därför ligger landet sörjande, och allt som lever där försmäktar både djuren på marken och fåglarna under himmelen; själva fiskarna i havet förgås.
Dock bör man icke så mycket gå till rätta med någon annan eller förebrå honom, eller förebrå ditt folk, som man bör gå till rätta med prästen.
Ja, du skall komma på fall om dagen, på fall skall ock profeten komma jämte dig om natten, jämväl din moder skall jag förgöra.
Det är förbi med mitt folk, därför att det ej får någon kunskap.
Men eftersom du har förkastat kunskap, därför skall ock jag förkasta dig, så att du upphör att vara min präst.
Och såsom du har förgätit din Guds lag, så skall ock jag förgäta dina barn.
Ju mer de hava fått växa till, dess mer hava de syndat mot mig; men deras ära skall jag förbyta i skam.
Av mitt folks synd föda de sig, och till dess missgärning står deras begår.
Men nu skall det gå prästen och folket lika: jag skall hemsöka dem för deras vägar, och för deras gärningar skall jag vedergälla dem.
När de äta, skola de icke bliva mätta, och genom sitt lösaktiga leverne skola de ej föröka sig; de hava ju upphört att hålla sig till HERREN.
Lösaktighet och vin och must taga bort förståndet.
Mitt folk frågar sin stock till råds och vill hämta besked av sin stav; ty en trolöshetens ande har fört dem vilse, så att de i trolös avfällighet hava lupit bort ifrån sin Gud.
På bergens toppar frambära de offer, och på höjderna tända de offereld, under ekar, popplar och terebinter, eftersom skuggan där är så god.
Så bliva edra döttrar skökor, och edra söners hustrur äktenskapsbryterskor.
Dock kan jag icke straffa edra döttrar för att de äro skökor, eller edra söners hustrur för att de äro äktenskapsbryterskor, ty männen själva gå ju avsides med skökor, och offra med tempeltärnor.
Så löper folket, som intet förstår, till sin undergång.
Om nu du Israel vill bedriva din otukt, så må dock Juda icke ådraga sig skuld.
Kommen då icke till Gilgal, dragen ej upp till Bet-Aven, och svärjen icke: »Så sant HERREN lever.»
Om Israel spjärnar emot såsom en obändig ko, månne HERREN ändå skall föra dem i bet såsom lamm i vida öknen
Nej, Efraim står i förbund med avgudar; må han då fara!
Deras dryckenskap är omåttlig. hejdlöst bedriva de sin otukt; de som skulle vara landets sköldar älska vad skamligt är.
Men en stormvind skall fatta dem med sina vingar, och de skola komma på skam med sina offer.
Hören detta, I präster, akten härpå, I av Israels hus, och I av konungens hus, lyssnen härtill; ty eder gäller domen.
Ty I haven varit en snara för Mispa och ett nät, utbrett på Tabor.
Mitt under sitt offrande har man sjunkit allt djupare, men jag skall bliva ett tuktoris för allasammans.
Jag känner Efraim, och Israel är icke fördold för mig.
Du Efraim, du har ju nu blivit en sköka, Israel har orenat sig.
De lägga sig icke vinn om att vända tillbaka till sin Gud, ty en trolöshetens ande bor i deras bröst, och HERREN känna de icke.
Men Israels stolthet vittnar emot honom, och Israel och Efraim komma på fall genom sin missgärning; Juda kommer ock på fall jämte dem.
Om de än med får och fäkreatur gå åstad för att söka HERREN, så finna de honom ändå icke; han har dragit sig undan från dem.
Mot HERREN hava de handlat trolöst, ja, de hava fött barn som icke äro hans.
Därför skall nu en nymånadsdag förtära dem, jämte det som de fingo på sin del.
Stöten i basun i Gibea, i trumpet i Rama, blåsen larmsignal i Bet-Aven.
Fienden är efter dig, Benjamin!
Efraim skall varda ödelagt på straffets dag; mot Israels stammar kungör jag vad visst är.
Juda furstar hava blivit råmärkflyttares likar; över dem skall jag utgjuta min vrede såsom vatten.
Efraim lider förtryck, och hans rätt våldföres, ty han har tagit sig till att vandra efter tomma stadgar.
Därför är jag nu för Efraim såsom mal och för Juda hus såsom röta i benen.
Och Efraim har märkt sin sjukdom och Juda sitt sår; därför har Efraim gått till Assur och sänt bud till Jarebs-konungen.
Men denne skall icke kunna hela eder; edert sår skall icke bliva läkt.
Ty jag skall vara såsom ett lejon mot Efraim och såsom ett ungt lejon mot Juda hus.
Själv griper jag mitt rov och går bort därmed; jag släpar det bort utan räddning.
Jag vill gå min väg, tillbaka till min boning, till dess att de hava fått lida vad de hava förskyllt och begynna söka mitt ansikte.
Ja, i sin nöd skola de söka mig: »Kommen, låtom oss vända om till HERREN.
Ty han har sargat oss, han skall ock hela oss.
Han har slagit oss, han skall ock förbinda oss.
Han skall om två dagar åter göra oss helbrägda; ja, på tredje dagen skall han låta oss stå upp, så att vi få leva inför honom.
Så låtom oss lära känna HERREN, ja, låtom oss fara efter att lära känna honom.
Hans uppgång är så viss som morgonrodnadens, och han skall komma över oss lik ett regn, lik ett vårregn, som vattnar jorden.»
Vad skall jag taga mig till med dig Efraim?
Vad skall jag taga mig till med dig, Juda?
Eder kärlek är ju lik morgonskyn, lik daggen, som tidigt försvinner.
Därför har jag utdelat mina hugg genom profeterna, därför har jag dräpt dem genom min muns tal; så skall domen över dig stå fram i ljuset.
Ty jag har behag till kärlek och icke till offer, och till Guds kunskap mer än till brännoffer.
Men dessa hava på människovis överträtt förbundet; däri hava de handlat trolöst mot mig.
Gilead är en stad av ogärningsmän, den är full med blodiga spår.
Och lik en rövarskara, som ligger i försåt för människor, är prästernas hop.
De mörda på vägen till Sikem, ja, vad skändligt är göra de.
I Israels hus har jag sett gruvliga ting; där bedriver Efraim sin otukt, där orenar sig Israel.
Också för dig, Juda, är en skördetid bestämd, när jag åter upprättar mitt folk.
När jag vill hela Israel, då uppenbarar sig Efraims missgärning och Samariens ondska.
Ty de öva falskhet, tjuvar göra inbrott, rövarskaror plundra på vägarna.
Och de betänka icke i sina hjärtan att jag lägger all deras ondska på minnet.
De äro nu kringrända av sina egna gärningar, ty dessa hava kommit inför mitt ansikte.
Med sin ondska bereda de konungen glädje och med sina lögner furstarna.
Allasammans äro de äktenskapsbrytare; de likna en ugn, upphettad av bagaren, som när han har knådat degen, underlåter att elda, till dess att degen är syrad.
På vår konungs dag drucko sig furstarna febersjuka av vin; själv räckte han bespottarna handen.
När de med sina anslag hava eldat upp sitt hjärta likasom en ugn, sover bagaren hela natten; men om morgonen brinner elden i ljus låga.
Allasammans äro de heta såsom en ugn och förbränna så sina domare; ja, alla deras konungar falla, ty bland dem finnes ingen som åkallar mig.
Efraim beblandar sig med andra folk; Efraim har blivit lik en ovänd kaka.
Främlingar hava förtärt hans kraft, men han förstår intet; fastän han har fått grå hår, förstår han ändå intet.
Men Israels stolthet vittnar emot honom; de vända icke om till HERREN, sin Gud, och de söka honom ej, allt detta oaktat.
Efraim har blivit lik en duva, enfaldig, utan förstånd.
Egypten påkalla de, till Assur gå de;
men bäst de gå där, breder jag ut mitt nät över dem och drager dem ned, såsom vore de fåglar under himmelen.
Ja, jag skall tukta dem, såsom det redan har sports i deras församling.
Ve över dem, ty de hava flytt bort ifrån mig!
Fördärv över dem, ty de hava avfallit från mig!
Och jag skulle förlossa dem, dem som föra mot mig så lögnaktigt tal!
De ropa icke till mig av hjärtat, allenast jämra sig på sina läger; de hava ångest för sin säd och sitt vin, men de äro gensträviga mot mig.
Det var jag som undervisade dem och stärkte deras armar, men de hava ont i sinnet mot mig.
De vända om, men icke till den som är därovan; de äro lika en båge som sviker.
Deras furstar skola falla genom svärd, därför att deras tungor äro så hätska.
Då skall man bespotta dem i Egyptens land.
Sätt basunen för din mun! »Såsom en örn kommer fienden över HERRENS hus, eftersom de hava överträtt mitt förbund och avfallit från min lag.
De ropa till mig: »Min Gud!
Vi känna dig, vi av Israel.»
Men eftersom Israel har förkastat vad gott är, skall fienden jaga honom.
Själva valde de sig konungar, som icke kommo från mig; de tillsatte furstar, utan att jag fick veta något därom av sitt silver och guld gjorde de sig avgudar, ty det skulle ju förstöras.
En styggelse är din kalv, Samarien!
Min vrede är upptänd mot dessa människor; huru länge skola de kunna undgå straff?
Från Israel har ju kalven kommit; en konstarbetare har gjort honom, och en gud är han icke.
Nej, Samariens kalv skall bliva krossad till smulor.
Ty vind så de, och storm skola de skörda.
Säd skola de icke få, deras gröda skall icke giva någon föda, och giver den någon, skola främlingar uppsluka den.
Uppslukad varder Israel!
Redan aktas de bland hedningarna såsom ett värdelöst ting.
Ty väl hava de dragit åstad upp till Assur, lika vildåsnor som gå sin egen väg, ja, väl vill Efraim köpslå om älskog;
men huru de än köpslå bland hedningarna, skall jag dock nu tränga dem tillhopa och låta dem begynna en tid av ringhet, under överkonungens förtryck.
Eftersom Efraim har gjort sig så många altaren till synd, skola ock hans altaren bliva honom till synd.
Om jag än skriver mina lagar för honom i tiotusental, så räknas de ju dock för en främlings lagar.
Såsom slaktoffergåvor åt mig offrar man kött som man sedan äter upp; HERREN har intet behag till sådana.
Nu kommer han ihåg deras missgärning och hemsöker deras synder; till Egypten skola de få vända tillbaka.
Och eftersom Israel har förgätit sin skapare och byggt sig palatser, och eftersom Juda har uppfört så många befästa städer, skall jag sända en eld mot hans städer, och den skall förtära palatsen i dem.
Gläd dig icke, Israel, så att du jublar såsom andra folk, du som i trolös avfällighet har lupit bort ifrån din Gud, du som har haft ditt behag i skökolön på alla sädeslogar.
Logen och vinpressen skola icke föda dem, och vinet skall slå fel för dem.
De skola icke få bo i HERRENS land; Efraim måste vända tillbaka till Egypten, och i Assyrien skola de nödgas äta vad orent är.
De skola ej få offra vin till drickoffer åt HERREN och skola icke vinna hans välbehag.
Deras slaktoffer skola vara för dem såsom sorgebröd; alla som äta därav skola bliva orena.
Ty det bröd de få stillar allenast deras hunger, det kommer icke in i HERRENS hus.
Vad skolen I då göra, när en högtidsdag kommer, en HERRENS festdag?
Ty se, om de undgå förödelsen, bliver det Egypten som får församla dem, Mof som får begrava dem.
Deras silver, som är dem så kärt, skola nässlor taga i besittning; törne skall växa i deras hyddor.
De komma, hemsökelsens dagar!
De komma, vedergällningens dagar!
Israel skall förnimma det.
Såsom en dåre står då profeten, såsom en vanvetting andans man, för din stora missgärnings skull; ty stor har din hätskhet varit.
Ja, en lurande fiende är Efraim mot min Gud; för profeten sättas fällor på alla hans vägar och utläggas snaror i hans Guds hus.
I djupt fördärv äro de nedsjunkna, nu såsom i Gibeas dagar.
Men han kommer ihåg deras missgärning, han hemsöker deras synder.
Såsom druvor i öknen fann jag Israel; jag såg edra fäder såsom förstlingsfrukter på ett fikonträd, då det begynner bära frukt.
Men när de kommo till Baal-Peor, invigde de sig åt skändlighetsguden och blevo en styggelse lika honom som de älskade.
Efraims härlighet skall flyga sin kos såsom en fågel; ingen skall där föda barn eller gå havande, ingen bliva fruktsam.
Och om de än få uppföda barn åt sig, skall jag taga dessa ifrån dem, så att ingen människa bliver kvar.
Ja, ve dem själva, när jag viker ifrån dem!
Väl är Efraim nu vad jag har sett Tyrus vara, en plantering på ängen; men Efraim skall en gång få föra ut sina söner till bödeln.
Giv dem, HERRE, vad du bör giva dem.
Giv dem ofruktsamma moderssköten och försinade bröst.
All deras ondska är samlad i Gilgal; ja, där fick jag hat till dem För deras onda väsendes skull vill jag driva dem ut ur mitt hus.
Jag skall icke längre bevisa dem kärlek; alla deras styresmän äro ju upprorsmän.
Efraim skall bliva nedbruten; deras rot skall förtorkas, de skola ej bära någon frukt.
Om de ock föda barn, skall jag döda deras livsfrukt, huru kär den än är dem.
Ja, min Gud skall förkasta dem, eftersom de icke ville höra honom; de skola bliva flyktingar bland hedningarna.
Israel var ett frodigt vinträd, som satte frukt.
Men ju mer frukt han fick, dess flera altaren gjorde han åt sig; ju bättre det gick hans land, dess präktigare stoder reste han.
Deras hjärtan voro hala; nu skola de lida vad de hava förskyllt.
Han skall själv bryta ned deras altaren, förstöra deras stoder.
Ja, nu skola de få säga: »Vi hava blivit utan konung, därför att vi icke fruktade HERREN.
Dock, en konung, vad skulle nu han kunna göra för oss?»
De tala tomma ord, de svärja falska eder, de sluta förbund; men såsom en bitter planta skjuter domen upp ur markens fåror.
För kalvarna i Bet-Aven skola Samariens inbyggare få bekymmer; ja, för en sådan skall hans folk hava sorg, och hans präster skola skria för hans skull, när hans skatter föras bort från honom.
Också han själv skall bliva släpad till Assyrien såsom en skänk åt Jarebs-konungen.
Skam skall Efraim uppbära, Israel skall komma på skam med sina rådslag.
Det är förbi med Samariens konung; såsom ett spån på vattnet far han hän.
Ödelagda bliva Avens offerhöjder, som Israel så har försyndat sig med; törne och tistel skall skjuta upp på deras altaren.
Då skall man säga till bergen: »Skylen oss», och till höjderna: »Fallen över oss.»
Israels synd når tillbaka ända till Gibeas dagar; där hava de förblivit stående.
Icke skulle hämndekriget mot de orättfärdiga kunna nå dem i deras Gibea?
Jo, när mig så lyster, tuktar jag dem; då skola folken församlas mot dem och oka dem ihop med deras båda missgärningsverk.
Efraim har varit en hemtam kalv, som fann behag i att gå på trösklogen; och jag har skonat hans frodiga hals.
Nu skall jag spänna Efraim i oket, Juda skall gå för plogen, Jakob för harven.
Sån ut åt eder i rättfärdighet, skörden efter kärlekens bud, bryten eder ny mark; ty det är tid att söka HERREN, för att han skall komma och låta rättfärdighet regna över eder.
I haven plöjt ogudaktighet, orättfärdighet haven I skördat, I haven ätit lögnaktighets frukt, i förlitande på eder väg, på edra många hjältar.
Men ett stridslarm skall uppstå bland edra stammar, och alla edra fästen skola ödeläggas, såsom Bet-Arbel ödelades av Salman på stridens dag, då man krossade både mödrar och barn.
Sådant skall Betel tillskynda eder, för eder stora ondskas skull.
När morgonrodnaden går upp, är det förbi, förbi med Israels konung!
När Israel var ung, fick jag honom kär, och ut ur Egypten kallade jag min son.
Men ju mer de hava blivit kallade, dess mer hava de dragit sig undan; de frambära offer åt Baalerna, och åt belätena tända de offereld.
Och likväl var det jag som lärde Efraim att gå, och som tog dem upp i mina armar.
Men de förstodo icke att jag ville hela dem.
Med lena band drog jag dem, med kärlekens tåg; jag lättade oket över deras halsar, jag sänkte mig ned till dem och gav dem föda.
Borde de då icke få vända tillbaka till Egyptens land eller få Assur till sin konung, eftersom de icke vilja omvända sig?
Ja, svärdet skall rasa i deras städer och förstöra deras bommar och frossa omkring sig, för deras anslags skull.
Ty mitt folks håg står till avfall från mig; och huru mycket man än kallar dem till den som är därovan, så höjer sig ändå ingen.
Men huru skall jag kunna giva dig till pris, Efraim, och låta dig fara, Israel?
Icke kan jag giva dig till pris såsom Adma och låta det gå dig såsom Seboim?
Mitt hjärta vänder sig i mig, all min barmhärtighet vaknar.
Jag vill icke låta dig känna min vredes glöd, jag skall icke vidare fördärva Efraim.
Ty jag är Gud och icke en människa; helig är jag bland eder, och med vrede vill jag ej komma.
Efter HERREN skola de så draga åstad, och han skall ryta såsom ett lejon; ja, han skall upphäva ett rytande, och hans barn skola då med bävan samlas västerifrån;
såsom fåglar skola de med bävan komma från Egypten och såsom duvor från Assurs land.
Och sedan skall jag låta dem bo kvar i sina hus, säger HERREN.
Efraim har omvärvt mig med lögn och Israels hus med svek Juda är alltjämt trolös mot Gud, mot den Helige, den Trofaste.
Efraim jagar efter vind och far efter östanväder; beständigt går han framåt i lögn och våld.
Med Assur sluter man förbund, och olja för man till Egypten.
Men HERREN skall gå till rätta med Juda och hemsöka Jakob, såsom hans vägar förtjäna; efter hans gärningar skall han vedergälla honom.
I moderlivet grep han sin broder i hälen, och i sin mandomskraft kämpade han med Gud.
Ja, han kämpade med ängeln och vann seger, han grät och bad honom om nåd.
I Betel mötte han honom, och där talade han med oss.
Och HERREN, härskarornas Gud, »HERREN» är hans namn.
Så vänd nu om till din Gud; håll fast vid kärlek och rätt, och förbida din Gud beständigt.
Kanaans folk går med falsk våg i sin hand, det älskar orättrådig vinning;
så säger ock Efraim: »Jag har ju blivit rik, jag har förvärvat mig gods; vad jag än gör, skall det ej draga över mig skuld som kan räknas för synd.»
Men jag som är HERREN, din Gud, alltsedan du var i Egyptens land, jag skall återigen låta dig bo i tält, likasom vid eder högtid.
Jag har talat till profeterna, jag har låtit dem skåda mångahanda syner, och genom profeterna har jag talat i liknelser.
Är nu Gilead ett ogärningsnäste, där allenast falskhet råder, och offrar man tjurar i Gilgal, så skola ock deras altaren bliva lika stenrösen vid markens fåror.
Och Jakob flydde till Arams mark Israel tjänade för en kvinna, för en kvinnas skull vaktade han hjorden.
Men genom en profet förde HERREN Israel upp ur Egypten, och genom en profet blev folket bevarat.
Efraim har uppväckt bitter förtörnelse; hans Herre skall låta hans blodskulder drabba honom och låta hans smädelser falla tillbaka på honom själv.
Så ofta Efraim tog till orda, uppstod skräck; högt tronade han i Israel.
Men han ådrog sig skuld genom Baal och måste så dö.
Och ännu fortgå de i sin synd; av sitt silver göra de sig gjutna beläten, avgudar efter sitt eget förstånd, alltsammans konstarbetares verk.
Till sådana ställa de sina böner; under det att de slakta människor, giva de sin hyllningskyss åt kalvar.
Därför skola de bliva lika morgonskyn, lika daggen som tidigt försvinner, lika agnar som blåsa bort ifrån tröskplatsen och lika rök som flyr hän ur ett rökfång.
Men jag är HERREN, din Gud, alltsedan du var i Egyptens land; utom mig vet du ej av någon Gud, och ingen annan frälsare finnes än jag.
Det var jag som lät mig vårda om dig i öknen, i den brännande torkans land.
Men ju bättre bete de fingo, dess mättare blevo de, och när de voro mätta till fyllest, blevo deras hjärtan högmodiga; och så glömde de mig.
Då blev jag mot dem såsom ett lejon; lik en panter lurar jag nu vid vägen.
Jag kommer över dem såsom en björninna från vilken man har tagit ungarna, jag river sönder deras hjärtans hölje; jag uppslukar dem på stället, lik en lejoninna, lik ett vilddjur som söndersliter dem.
Det har blivit ditt fördärv, o Israel, att du satte dig upp mot mig som var din hjälp.
Var är nu din konung, som skulle bereda dig frälsning i alla dina städer?
Och var har du dina domare, du som sade: »Låt mig få konung och furstar»?
Ja, en konung skall jag giva dig i min vrede, och i min förgrymmelse skall jag åter taga honom bort.
Efraims missgärning är samlad såsom i en pung, och hans synd är i förvar.
En barnaföderskas vånda skall komma över honom.
Han är ett oförnuftigt foster, som icke kommer fram i födseln. när tiden är inne.
Skulle jag förlossa sådana ur dödsrikets våld, köpa dem fria ifrån döden? -- Var har du dina hemsökelser, du död?
Var har du din pest, du dödsrike?
Ånger må vara fördold för mina ögon.
Bäst han står där frodig bland sina bröder skall en östanvind komma, ett HERRENS väder, som stiger upp från öknen; då skall hans brunn komma på skam och hans källa sina ut.
Den vinden rycker bort de skatter han har samlat av alla slags dyrbara håvor.
Samarien skall lida vad det har förskyllt genom sin gensträvighet mot sin Gud.
Inbyggarna skola falla för svärd, deras späda barn skola bliva krossade och deras havande kvinnor skall man upprista.
Vänd om, o Israel, till HERREN, din Gud; ty genom din missgärning har du kommit på fall.
Tagen med eder böneord, och vänden så åter till HERREN; sägen till honom: »Skaffa bort all missgärning, och tag fram goda håvor, så vilja vi hembära dig våra läppars offer, såsom man offrar tjurar.
Hos Assur skola vi ej mer söka vår frälsning, vi skola icke vidare stiga till häst. våra händers verk skola vi icke mer kalla för vår Gud.
Ty hos dig är det som den faderlöse undfår barmhärtighet.»
Ja, deras avfällighet vill jag hela, jag vill bevisa dem kärlek av hjärtat, ty min vrede har vänt sig ifrån dem.
Jag skall bliva för Israel såsom dagg, han skall blomstra såsom en lilja, och såsom Libanons skog skall han skjuta rötter.
Telningar skola utgå från honom, han skall bliva lik ett olivträd i fägring och doft skall han sprida såsom Libanon.
De som bo i hans skugga skola åter få odla säd och skola grönska såsom vinträd; hans namn skall vara såsom Libanons vin.
Men vad har jag då mer att skaffa med avgudarna, du Efraim!
Jag själv vill ju giva bönhörelse och se till honom.
Ja, lik en grönskande cypress vill jag bliva; hos mig skall finnas frukt att hämta för dig.
Den som är vis, han akte härpå; den som är förståndig, han besinne detta.
Ty HERRENS vägar äro rätta, och på dem vandra de rättfärdiga, men överträdarna komma där på fall.
Detta är HERRENS ord som kom till Joel, Petuels son.
Hören detta, I gamle, och lyssnen härtill, I landets alla inbyggare.
Har något sådant skett förut i edra dagar eller i edra fäders dagar?
Nej, om detta mån I förtälja för edra barn, och edra barn må förtälja därom för sina barn, och deras barn för ett kommande släkte.
Vad som blev kvar efter gräsgnagarna, det åto gräshopporna upp; och vad som blev kvar efter gräshopporna, det åto gräsbitarna upp; och vad som blev kvar efter gräsbitarna det åto gräsfrätarna upp.
Vaknen upp, I druckne, och gråten; ja, jämren eder, alla I som dricken vin, över att druvsaften är ryckt undan eder mun.
Ty ett folk har dragit upp över mitt land, ett mäktigt, ett som ingen kan räkna; det har tänder likasom lejon, och dess kindtänder likna lejoninnors.
Mina vinträd har det förött, och mina fikonträd har det brutit ned det har skalat dem nakna och kastat dem undan; vitnade äro deras rankor.
Klaga likasom en jungfru som bär sorgdräkt efter sin ungdoms brudgum
Spisoffer och drickoffer äro försvunna ifrån HERRENS hus; prästerna sörja, HERRENS tjänare.
Fälten äro förödda, marken ligger sörjande, ty säden är förödd, vinet borttorkat, oljan utsinad.
Åkermännen stå med skam, vingårdsmännen jämra sig, över vetet och över kornet; ty skörden på marken är förstörd.
Vinträden äro förtorkade och fikonträden försmäkta; granatträden och palmerna och äppelträden och alla andra träd på marken hava torkat bort.
Ja, all fröjd har vissnat och flytt ifrån människors barn.
Kläden eder i sorgdräkt och klagen, I präster; jämren eder, I som tjänen vid altaret; gån in och sitten i sorgdräkt natten igenom, I min Guds tjänare, eftersom eder Gud hus måste sakna spisoffer och drickoffer
Pålysen en helig fasta, lysen ut en högtidsförsamling; församlen de gamla, ja, alla landets inbyggare, till HERRENS, eder Guds, hus; och ropen så till HERREN.
Ve oss, vilken dag! ty HERRENS dag är nära, och såsom våld från den Allsvåldige kommer den.
Har icke vår bärgning blivit förstörd mitt för våra ögon? har icke glädje och fröjd försvunnit ifrån var Guds hus?
Utsädet ligger förtorkat under mullen, förrådshusen stå öde, ladorna få förfalla, ty säden är borttorkad.
Huru stönar icke boskapen!
Huru ängslas ej fäkreaturens hjordar!
De finna ju intet bete.
Ja, också fårhjordarna få lida under skulden.
Till dig, HERRE, ropar jag, nu då en eld har förtärt betesmarkerna i öknen och en eldslåga har förbränt alla träd på marken.
Ja, också markens djur ropa med trängtan till dig, eftersom vattenbäckarna äro uttorkade och betesmarkerna i öknen äro förtärda av eld.
Stöten i basun på Sion, och blåsen larmsignal på mitt heliga berg; må alla landets inbyggare darra!
Ty HERRENS dag kommer, ja, den är nära;
en dag av mörker och tjocka, en dag av moln och töcken, lik en gryning som breder ut sig över bergen.
Ett stort och mäktigt folk kommer, ett vars like aldrig någonsin har funnits och ej heller hädanefter skall uppstå, intill senaste släktens år.
Framför dem går en förtärande eld och bakom dem kommer en förbrännande låga.
Likt Edens lustgård var landet framför dem, men bakom dem är det en öde öken; ja, undan dem finnes ingen räddning.
De te sig likasom hästar, och såsom stridshästar hasta de åstad.
Med ett rassel likasom av vagnar spränga de fram över bergens toppar, med ett brus såsom av en eldslåga, när den förtär strå; de äro såsom ett mäktigt folk, ordnat till strid.
Vid deras åsyn gripas folken av ångest, alla ansikten skifta färg.
Såsom hjältar hasta de åstad, lika stridsmän bestiga de murarna; var och en går sin väg rakt fram, och ingen tager miste om sin stråt.
Den ene tränger icke den andre, var och en går sin givna bana; mitt igenom vapnen störta de fram utan hejd.
I staden rusa de in på murarna hasta de åstad, i husen tränga de upp, genom fönstren bryta de sig väg, såsom tjuvar göra.
Vid deras åsyn darrar jorden, och himmelen bävar; solen och månen förmörkas, och stjärnorna mista sitt sken.
Och HERREN låter höra sin röst framför sin här ty hans skara är mycket stor, mäktig är den skara som utför hans befallning.
Ja, HERRENS dag är stor och mycket fruktansvärd vem kan uthärda den?
Dock, nu mån I vända om till mig av allt edert hjärta, säger HERREN, med fasta och gråt och klagan.
Ja, riven sönder edra hjärtan, icke edra kläder, och vänden om till HERREN, eder Gud; ty nådig och barmhärtig är han, långmodig och stor i mildhet, och sådan att han ångrar det onda.
Måhända vänder han om och ångrar sig och lämnar kvar efter sig någon välsignelse, till spisoffer och drickoffer åt HERREN, eder Gud.
Stöten i basun på Sion, pålysen en helig fasta lysen ut en högtidsförsamling;
församlen folket, pålysen en helig sammankomst, kallen tillhopa de gamla församlen de små barnen, jämväl dem som ännu dia vid bröstet brudgummen må komma ur sin kammare och bruden ur sitt gemak.
Mellan förhuset och altaret må prästerna, HERRENS tjänare, hålla klagogråt och säga: »HERRE, skona ditt folk, och låt icke din arvedel bliva till smälek, till ett ordspråk bland hedningarna Varför skulle man få säga bland folken: 'Var är nu deras Gud?'»
Så upptändes då HERREN till nitälskan för sitt land, och han ömkade sig över sitt folk;
HERREN svarade och sade till sitt folk: Se, jag vill sända eder säd och vin och olja, så att I fån mätta eder därav, och jag skall icke mer låta eder bliva till smälek bland hedningarna.
Och nordlandsskaran skall jag förjaga långt bort ifrån eder, jag skall driva den undan till ett torrt och öde Land, dess förtrupp till Östra havet och dess eftertrupp till Västra havet.
Och stank skall stiga upp därav, ja, vämjelig lukt skall stiga upp därav, eftersom den har tagit sig för så stora ting.
Frukta icke, du land, utan fröjda dig och gläds, ty stora ting har HERREN tagit sig för
Frukten icke, I markens djur, ty betesmarkerna i öknen grönska, och träden bära sin frukt, fikonträden och vinträden giva sin kraft.
Och fröjden eder, I Sions barn, varen glada i HERREN, eder Gud; ty han giver eder höstregn, i rätt tid, han som ock förr sände ned över eder regn, både höst och vår.
Så skola logarna fyllas mod säd och pressarna flöda över av vin och olja.
Och jag skall giva eder gottgörelse för de årsgrödor som åtos upp av gräshopporna, gräsbitarna, gräsätarna och gräsgnagarna, den stora här som jag sände ut mot eder.
Och I skolen få äta till fyllest och bliva mätta; och då skolen I lova HERRENS, eder Guds, namn, hans som har handlat så underbart med eder; och mitt folk skall icke komma på skam evinnerligen.
Och I skolen förnimma att jag bor mitt i Israel, och att jag är HERREN, eder Gud, och eljest ingen.
Ja, mitt folk skall icke komma på skam evinnerligen.
Och det skall ske därefter att jag skall utgjuta min Ande över allt kött, och edra söner och edra döttrar skola profetera, edra gamla män skola hava drömmar edra ynglingar skola se syner;
också över dem som äro tjänare och tjänarinnor skall jag i de dagarna utgjuta min Ande.
Och jag skall låta tecken synas på himmelen och på jorden: blod och eld och rökstoder.
Solen skall vändas i mörker och månen i blod förrän HERRENS dag kommer, den stora och fruktansvärda.
Men det skall ske att var och en som åkallar HERRENS namn han skall varda frälst.
Ty på Sions berg och i Jerusalem skall finnas en räddad skara, såsom HERREN har sagt; och till de undsluppna skola höra de som HERREN kallar.
Ty se, i de dagarna och på den tiden, då jag åter upprättar Juda och Jerusalem,
då skall jag samla tillhopa alla hednafolk och föra dem ned till Josafats dal, och där skall jag hålla dom över dem, för mitt folks och min arvedels, Israels, skull, därför att de hava förskingrat dem bland hedningarna och utskiftat mitt land.
Ja, de hava kastat lott om mitt folk, gossarna hava de givit såsom betalning åt skökor, och flickorna hava de sålt för vin, som de hava druckit upp.
Och du, Tyrus, och du, Sidon, och I, Filisteens alla kretsar, vad förehaven också I mot mig?
Haven I något att vedergälla mig för, eller är det I som viljen begynna något mot mig?
Snart och med hast skall jag låta det I haven gjort komma tillbaka över edra egna huvuden,
eftersom I haven tagit mitt silver och mitt guld och fört mina skönaste klenoder in i edra palats,
och eftersom I haven sålt Judas och Jerusalems barn åt Javans barn, till att föras långt bort ifrån sitt land.
Se, jag skall kalla dem åter från den ort dit I haven sålt dem; och det som I haven gjort skall jag låta komma tillbaka över edra egna huvuden.
Jag skall sälja edra söner och döttrar i Juda barns hand, och de skola sälja dem till sabéerna, folket i fjärran land.
Ty så har HERREN talat.
Ropen ut detta bland hednafolken, båden upp dem till helig strid.
Manen på hjältarna, må alla stridsmännen komma och draga framåt.
Smiden edra plogbillar till svärd och edra vingårdsknivar till spjut; den svagaste må känna sig såsom en hjälte.
Skynden att komma, alla I folk har omkring, och samlen eder tillhopa.
Sänd, o HERRE, ditned dina hjältar.
Ja, må hednafolken resa sig och draga åstad till Josafats dal; ty där skall jag sitta till doms över alla folk häromkring.
Låten lien gå, ty skörden är mogen.
Kommen och trampen, ty pressen är full; presskaren flöda över, så stor är ondskan där.
Skaror hopa sig i Domens dal; ty HERRENS dag är nära i Domens dal.
Solen och månen förmörkas, och stjärnorna mista sitt sken.
Och HERREN upphäver ett rytande från Sion, och från Jerusalem låter han höra sin röst, så att himmelen och jorden bäva.
Men för sitt folk är HERREN en tillflykt och för Israels barn ett värn.
Och I skolen förnimma att jag är HERREN, eder Gud, som bor på Sion, mitt heliga berg.
Och Jerusalem skall vara en helgad plats och främlingar skola icke mer draga ditin.
På den tiden skall det ske att bergen drypa av druvsaft och höjderna flöda av mjölk; och alla bäckar i Juda skola flöda av vatten.
Och en källa skall rinna upp i HERRENS hus och vattna Akaciedalen.
Men Egypten skall bliva en ödemark, och Edom skall varda en öde öken därför att de hava övat våld mot Juda barn och utgjutit oskyldigt blod i sitt land.
Sedan skall Juda trona evinnerligen, och Jerusalem från släkte till släkte.
Och jag skall utplåna deras blodskulder, dem som jag icke allaredan har utplånat.
Och HERREN skall förbliva boende på Sion.
Detta är vad som talades av Amos, en bland herdarna från Tekoa, vad han skådade angående Israel i Ussias, Juda konungs, och Jerobeams, Joas' sons, Israels konungs, tid, två år före jordbävningen.
Han sade: HERREN upphäver ett rytande från Sion, och från Jerusalem låter han höra sin röst.
Då försänkas herdarnas betesmarker i sorg, och Karmels topp förtorkas.
Så säger HERREN: Eftersom Damaskus har trefalt förbrutit sig, ja, fyrfalt, skall jag icke rygga mitt beslut: eftersom de hava tröskat Gilead med sina tröskvagnar av järn.
Därför skall jag sända en eld mot Hasaels hus, och den skall förtära Ben-Hadads palatser.
Jag skall bryta sönder Damaskus' bommar och utrota invånarna i Bikeat-Aven och spirans bärare i Bet-Eden; och Arams folk skall bliva bortfört till Kir, säger HERREN.
Så säger HERREN: Eftersom Gasa har trefalt förbrutit sig, ja, fyrfalt, skall jag icke rygga mitt beslut: eftersom de hava fört bort allt folket såsom fångar och överlämnat dem åt Edom.
Därför skall jag sända en eld mot Gasas murar, och den skall förtära dess palatser.
Jag skall utrota invånarna i Asdod och spirans bärare i Askelon; och jag skall vända min hand mot Ekron, så att filistéernas sista kvarleva förgås, säger Herren, HERREN.
Så säger HERREN: Eftersom Tyrus har trefalt förbrutit sig, ja, fyrfalt, skall jag icke rygga mitt beslut: eftersom de hava överlämnat allt folket såsom fångar åt Edom, utan att tänka på sitt brödraförbund.
Därför skall jag sända en eld mot Tyrus' murar, och den skall förtära dess palatser.
Så säger HERREN: Eftersom Edom har trefalt förbrutit sig, ja, fyrfalt, skall jag icke rygga mitt beslut: eftersom han har förföljt sin broder med svärd och förkvävt all barmhärtighet, och eftersom han oupphörligt har låtit sin vrede rasa och ständigt behållit sin förgrymmelse.
Därför skall jag sända en eld mot Teman, och den skall förtära Bosras palatser.
Så säger HERREN: Eftersom Ammons barn hava trefalt förbrutit sig, ja, fyrfalt, skall jag icke rygga mitt beslut: eftersom de hava uppristat havande kvinnor i Gilead, när de ville utvidga sitt område.
Därför skall jag tända upp en eld mot Rabbas murar, och den skall förtära dess palatser, under härskri på stridens dag, under storm på ovädrets dag.
Och deras konung skall vandra bort i fångenskap, han själv och hans hövdingar med honom, säger HERREN.
Så säger HERREN: Eftersom Moab har trefalt förbrutit sig, ja, fyrfalt, skall jag icke rygga mitt beslut: eftersom han har förbränt Edoms konungs ben till aska.
Därför skall jag sända en eld mot Moab, och den skall förtära Keriots palatser; och Moab skall omkomma under stridslarm, under härskri vid basuners ljud,
Och jag skall utrota ur landet den som är domare där, och alla dess furstar skall jag dräpa jämte honom säger HERREN.
Så säger HERREN: Eftersom Juda har trefalt förbrutit sig, ja, fyrfalt, skall jag icke rygga mitt beslut: eftersom de hava förkastat HERRENS lag och icke hållit hans stadgar, utan låtit förleda sig av sina lögngudar, dem som ock deras fäder vandrade efter.
Därför skall jag sända en eld mot Juda, och den skall förtära Jerusalems palatser.
Så säger HERREN: Eftersom Israel har trefalt förbrutit sig, ja, fyrfalt, skall jag icke rygga mitt beslut: eftersom de sälja den oskyldige för penningar och den fattige för ett par skor.
Ty de längta efter att se stoft på de armas huvuden, och de vränga de ödmjukas sak.
Son och fader gå tillsammans till tärnan och ohelga så mitt heliga namn.
På pantade kläder sträcker man sig invid vart altare, och bötfälldas vin dricker man i sin Guds hus
Och dock var det jag som förgjorde för dem amoréerna, ett folk så högrest som cedrar och så väldigt som ekar; jag förgjorde deras frukt ovantill och deras rötter nedantill.
Det var jag som förde eder upp ur Egyptens land, och som ledde eder i öknen i fyrtio år, så att I intogen amoréernas land.
Och jag uppväckte somliga bland edra söner till profeter och somliga bland edra unga män till nasirer.
Är det icke så, I Israels barn? säger HERREN.
Men I gåven nasirerna vin att dricka, och profeterna bjöden I: »Profeteren icke.»
Se, därför skall jag låta ett gnissel uppstå i edert land, likt gnisslet av en vagn som är fullastad med kärvar.
Då skall ej ens den snabbaste finna någon undflykt, den starkaste har då intet gagn av sin kraft, och hjälten kan icke rädda sitt liv.
Bågskytten håller då icke stånd, den snabbfotade kan icke rädda sitt liv, ej heller kan ryttaren rädda sitt.
Ja, den som var modigast bland hjältarna skall på den dagen fly undan naken, säger HERREN.
Hören följande ord, som HERREN har talat mot eder, I Israels barn, ja, mot hela det släkte som jag har fört upp ur Egyptens land.
Så har han sagt:
Eder allena har jag utvalt bland alla släkter på jorden; därför skall jag ock hemsöka på eder alla edra missgärningar.
Färdas väl två tillsammans, utan att de hava blivit ense därom?
Ryter ett lejon i skogen, om det ej har funnit något rov?
Upphäver ett ungt lejon sin röst i kulan, utan att det har tagit ett byte?
Faller en fågel i snaran på marken, om intet garn har blivit utlagt för den?
Springer snaran upp från marken, utom när den gör någon fångst?
Eller stöter man i basun i en stad, utan att folket förskräckes?
Eller drabbas en stad av något ont, utan att HERREN har skickat det?
Sannerligen, Herren, HERREN gör alls intet utan att hava uppenbarat sitt råd för sina tjänare profeterna.
När lejonet ryter, vem skulle då icke frukta?
När Herren, HERREN talar, vem skulle då icke profetera?
Ropen ut över Asdods palatser och över palatsen i Egyptens land; sägen: Församlen eder till Samarias berg, och sen huru stor förvirring där råder, och huru man övar förtryck därinne.
Man förstår icke där att göra vad rätt är, säger HERREN; man hopar våld och fördärv i sina palats.
Därför säger Herren, HERREN så: Trångmål skall komma och omvärva landet, ditt starka fäste skall du mista, det skall störtas ned; och dina palats skola varda utplundrade.
Så säger HERREN: Likasom när en herde ur lejonets gap räddar allenast ett par benpipor eller snibben av ett öra, så skola Israels barn bliva räddade, desamma som nu i Samaria sitta i sina soffors hörn och på sina bäddars sidendamast.
Hören och betygen inför Jakobs hus, säger Herren, HERREN, härskarornas Gud:
Den dag då jag på Israel hemsöker dess överträdelser, då skall jag ock hemsöka Betels altaren, så att altarhornen bliva avhuggna och falla till jorden.
Och jag skall slå ned både vinterhus och sommarhus, och elfenbenshusen skola bliva förstörda, ja, en myckenhet av hus skall då få en ände, säger HERREN.
Hören detta ord, I Basans-kor på Samarias berg, I som förtrycken de arma och öven våld mot de fattiga, I som sägen till edra män: »Skaffen hit, så att vi få dricka.»
Herren, HERREN har svurit vid sin helighet: Se, dagar skola komma över eder, då man skall hämta upp eder med metkrokar och eder sista kvarleva med fiskkrokar.
Då skolen I söka eder ut, var och en genom närmaste rämna i muren, och eder Harmonsbild skolen I då kasta bort, säger HERREN.
Kommen till Betel och bedriven eder synd till Gilgal och bedriven än värre synd; frambären där på morgonen edra slaktoffer, på tredje dagen eder tionde.
Förbrännen syrat bröd till lovoffer, lysen ut och kungören frivilliga offer.
Ty sådant älsken I ju, I Israels barn, säger Herren, HERREN.
Jag lät eder gå med tomma munnar i alla edra städer, jag lät eder sakna bröd på alla edra orter.
Och likväl haven I icke omvänt eder till mig, säger HERREN.
Jag förhöll regnet för eder, när ännu tre månader återstodo till skördetiden; jag lät det regna över en stad, men icke över en annan; en åker fick regn, men en annan förtorkades, i det att regn icke kom därpå.
Ja, två, tre städer måste stappla bort till en och samma stad för att få vatten att dricka, utan att de ändå kunde släcka sin törst.
Och likväl haven I icke omvänt eder till mig, säger HERREN.
Jag slog eder säd med sot och rost; edra många trädgårdar och vingårdar, edra fikonträd och olivträd åto gräsgnagarna upp.
Och likväl haven I icke omvänt eder till mig, säger HERREN.
Jag sände ibland eder pest, likasom i Egypten; jag dräpte edra unga män med svärd och lät edra hästar bliva tagna såsom byte; och stanken av edra fallna skaror lät jag stiga upp och komma eder i näsan.
Och likväl haven I icke omvänt eder till mig, säger HERREN.
Jag lät omstörtning drabba eder, likasom när Gud omstörtade Sodom och Gomorra; och I voren såsom en brand, ryckt ur elden.
Och likväl haven I icke omvänt eder till mig, säger HERREN.
Därför skall jag göra så med dig, Israel; och eftersom jag nu skall göra så med dig, därför bered dig, Israel, att möta din Gud.
Ty se, han som har danat bergen och skapat vinden, han som kan yppa för människan hennes hemligaste tankar, han som kan göra morgonrodnaden till mörker, och som går fram över jordens höjder -- HERREN, härskarornas Gud, är hans namn.
Hören följande ord, som jag vill uppstämma såsom klagosång över eder, I av Israels hus:
»Fallen är hon och kan icke mer stå upp, jungfrun Israel!
Hon ligger slagen till marken i sitt land; ingen reser henne upp.»
Ty så säger Herren, HERREN: Den stad varifrån tusen plägade draga ut skall få behålla hundra kvar, och den stad varifrån hundra plägade draga ut skall få behålla tio kvar, i Israels hus.
Ty så säger HERREN till Israels hus: Söken mig, så fån I leva.
Men söken icke Betel, kommen icke till Gilgal, och dragen ej bort till Beer-Seba; ty Gilgal skall bliva bortfört i fångenskap, och Betel skall hemfalla åt fördärvet.
Söken HERREN så fån I leva; varom icke, så skall han komma över Josefs hus lik en eld; och elden skall bränna, och ingen skall släcka den, till att rädda Betel.
I som förvandlen rätten till malört och slån rättfärdigheten ned till jorden, veten:
han som har gjort Sjustjärnorna och Orion, han som kan förvandla svarta mörkret till morgon och göra dagen mörk såsom natten, han som kallar på havets vatten och gjuter det ut över jorden -- HERREN är hans namn.
Och han låter fördärv ljunga ned över starka fästen; ja, över fasta borgar kommer fördärv.
Dessa hata i porten den som försvarar vad rätt är och räkna såsom en styggelse den som talar sanning.
Därför, eftersom I trampen på den arme och tagen ifrån honom hans säd såsom skatt, därför hören; om I än byggen hus av huggen sten, skolen I icke få bo i dem, och om I än planteren sköna vingårdar, skolen I icke få dricka vin från dem.
Ty jag vet att edra överträdelser äro många och edra synder talrika, I den rättfärdiges förtryckare, som tagen mutor och vrängen rätten för de fattiga i porten.
Därför måste den förståndige tiga stilla i denna tid; ty det är en ond tid.
Söken vad gott är, och icke vad ont är, på det att I mån leva.
Då skall Herren, härskarornas Gud, vara med eder, såsom I menen honom vara.
Haten vad ont är, och älsken vad gott är, och hållen rätten vid makt i porten; kanhända skall då Herren, härskarornas Gud, vara nådig mot Josefs kvarleva.
Därför, så säger HERREN, härskarornas Gud, Herren: På alla torg skall dödsklagan ljuda, och på alla gator skall man ropa: »Ack ve!
Ack ve!»
Åkermännen skall man mana att brista ut i jämmer, och dödsklagan skall höjas av dem som äro förfarna i sorgesång;
ja, i alla vingårdar skall dödsklagan ljuda, ty jag skall gå fram mitt ibland eder, säger HERREN.
Ve eder som åstunden HERRENS dag!
Vad viljen I med HERRENS dag?
Den är mörker och icke ljus.
Då går det, såsom när någon flyr för ett lejon, men därvid mötes av en björn, och när han då söker tillflykt i sitt hus, bliver han stungen av en orm, vid det han sätter handen mot väggen.
Ja, HERRENS dag är mörker och icke ljus, den är töcken utan något solsken.
Jag hatar edra fester, jag är led vid dem, och jag finner intet behag i edra högtidsförsamlingar.
Ty om I än offren åt mig brännoffer, jämte edra spisoffer, så har jag dock ingen lust till dem, ej heller gitter jag se edra tackoffer av gödda kalvar.
Hav bort ifrån mig dina sångers buller; jag gitter icke höra ditt psaltarspel.
Men må rätten flöda fram såsom vatten, och rättfärdigheten lik en bäck som aldrig sinar.
Framburen I väl åt mig slaktoffer och spisoffer under de fyrtio åren i öknen, I av Israels hus?
Så skolen I nu nödgas taga med eder Sickut, eder konung, och Kiun, eder avgudabild, stjärnguden, som I haven gjort åt eder;
och jag skall låta eder föras åstad i fångenskap ända bortom Damaskus, säger han vilkens namn är HERREN, härskarornas Gud.
Ve eder, I säkre på Sion, I sorglöse på Samarias berg, I ädlingar bland förstlingsfolket, I som Israels hus plägar vända sig till!
Gån åstad till Kalne och sen efter, dragen därifrån till Stora Hamat, och faren så ned till filistéernas Gat: äro de bättre än rikena här, eller är deras område större än edert område?
Ve eder, I som menen att olycksdagen skall vara fjärran, men likväl inbjuden våldet att trona hos eder;
I som liggen på soffor av elfenben och haven det makligt på edra bäddar; I som äten lamm, utvalda ur hjorden, och kalvar, hämtade från gödstallet;
I som skrålen visor till harpans ljud och tänken ut åt eder musikinstrumenter såsom David;
I som dricken vin ur stora bålar och bruken salvor av yppersta olja, men icke bekymren eder om Josefs skada!
Fördenskull skola nu dessa främst föras bort i fångenskap; de som nu hava det så makligt få då sluta med sitt skrål.
Herren, HERREN har svurit vid sig själv, säger HERREN, härskarornas Gud: Jakobs stolthet är mig en styggelse, och hans palatser hatar jag; jag skall giva staden till pris med allt vad däri är.
Och det skall ske, att om än tio män finnas kvar i ett och samma hus, så skola de likväl alla dö.
När sedan en frände till någon av de döda med förbrännarens hjälp vill skaffa benen ut ur huset, och därvid ropar till en som är i det inre av huset: »Finnes här någon mer än du?», då måste denne svara: »Ingen»; och den förre skall då säga: »Rätt så, stillhet må råda; ty HERRENS namn får icke bliva nämnt.»
Ty se, på HERRENS bud skola de stora husen bliva slagna i spillror och de små husen i splittror.
Kunna väl hästar springa uppför en klippbrant, eller plöjer man där med oxar? -- eftersom I viljen förvandla rätten till en giftplanta och rättfärdighetens frukt till malört,
I som glädjen eder över det som är intet värt och sägen: »Genom vår egen styrka hava vi ju berett oss horn.»
Ty se, jag skall uppväcka ett folk mot eder, I av Israels hus, säger Herren, härskarornas Gud; och de skola förtrycka edert land, från det ställe där vägen går till Hamat ända till Hedmarksbäcken.
Följande syn lät Herren, HERREN mig se; Jag såg gräshoppor skapas, när sommargräset begynte växa upp; och det var sommargräset efter kungsslåttern.
När så dessa hade ätit upp alla markens örter, sade jag: »Herre, HERRE, förlåt.
Huru skall Jakob kunna bestå, han som är så ringa?»
Då ångrade HERREN detta. »Det skall icke ske», sade HERREN.
Följande syn lät Herren, HERREN mig se: Jag såg Herren, HERREN nalkas för att utföra sin sak genom eld; och elden förtärde det stora djupet och höll på att förtära arvedelslandet.
Då sade jag: »Herre, HERRE, håll upp.
Huru skall Jakob kunna bestå, han som är så ringa?»
Då ångrade HERREN detta. »Icke heller detta skall ske», sade Herren, HERREN.
Följande syn lät han mig se: Jag såg Herren stå på en mur, uppförd efter sänklod, och i sin hand höll han ett sänklod.
Och HERREN sade till mig: »Vad ser du, Amos?»
Jag svarade: »Ett sänklod.»
Då sade Herren: »Se, jag skall hänga upp ett sänklod mitt ibland mitt folk Israel; jag kan icke vidare tillgiva dem.
Isaks offerhöjder skola bliva ödelagda och Israels helgedomar förstörda, och mot Jerobeams hus skall jag uppresa mig med svärdet.»
Men Amasja, prästen i Betel, sände till Jerobeam, Israels konung, och lät säga: »Amos förehar en sammansvärjning mot dig, mitt i Israels hus.
Landet kan icke härda ut med allt hans ordande.
Ty så har Amos sagt: 'Jerobeam skall dö för svärd, och Israel skall föras bort i fångenskap ur sitt land.'»
Och Amasja sade till Amos: »Du siare, gå din väg och sök din tillflykt i Juda land; där må du äta ditt bröd, och där må du profetera.
Men i Betel får du icke vidare profetera, ty det är en konungslig helgedom och ett rikets tempel.»
Då svarade Amos och sade till Amasja: »Jag är varken en profet eller en profetlärljunge, jag är en boskapsherde, som lever av mullbärsfikon.
Men HERREN tog mig från hjorden; HERREN sade till mig: 'Gå åstad och profetera för mitt folk Israel.'
Så hör nu HERRENS ord.
Du säger: 'Profetera icke mot Israel och predika icke mot Isaks hus.'
Därför säger HERREN så: Din hustru skall bliva en sköka i staden, dina söner och döttrar skola falla för svärd, ditt land skall bliva utskiftat med mätsnöre, själv skall du dö i ett orent land, och Israel skall föras bort i fångenskap ur sitt land.»
Följande syn lät Herren, HERREN mig se; Jag såg en korg med mogen frukt.
Och han sade: »Vad ser du, Amos?»
Jag svarade: »En korg med mogen frukt.»
Då sade HERREN till mig: »Mitt folk Israel är moget till undergång; jag kan icke vidare tillgiva dem.
Och sångerna i palatset skola på den dagen förbytas i jämmer, säger Herren, HERREN; man skall få se lik i mängd, överallt skola de ligga kastade; ja, stillhet må råda!»
Hören detta, I som stån den fattige efter livet och viljen göra slut på de ödmjuka i landet,
I som sägen: »När är då nymånadsdagen förbi, så att vi få sälja säd, och sabbaten, så att vi få öppna vårt sädesförråd?
Då vilja vi göra efa-måttet mindre och priset högre och förfalska vågen, så att den visar orätt vikt.
Då vilja vi köpa de arma för penningar och den fattige för ett par skor; och avfall av säden vilja vi då sälja såsom säd.»
HERREN har svurit vid Jakobs stolthet: Aldrig skall jag förgäta detta allt som de hava gjort.
Skulle jorden icke darra, när sådant sker, och skulle icke alla dess inbyggare sörja?
Skulle icke hela jorden höja sig såsom Nilen och röras upp och åter sjunka såsom Egyptens flod?
Och det skall ske på den dagen, säger Herren, HERREN, att jag skall låta solen gå ned i dess middagsglans och låta jorden sjunka i mörker mitt på ljusa dagen.
Jag skall förvandla edra högtider till sorgetider och alla edra sånger till klagovisor.
Jag skall hölja säcktyg kring allas länder och göra alla huvuden skalliga.
Jag skall låta det bliva, såsom när man sörjer ende sonen, och låta det sluta med en bedrövelsens dag.
Se dagar skola komma, säger Herren, HERREN, då jag skall sända hunger i landet: icke en hunger efter bröd, icke en törst efter vatten, utan efter att höra HERRENS ord.
Då skall man driva omkring från hav till hav, och från norr till öster, och färdas hit och dit för att söka efter HERRENS ord, men man skall icke finna det.
På den dagen skola de försmäkta av törst, edra sköna jungfrur och edra unga män,
desamma som nu svärja vid Samariens syndaskuld och säga: »Så sant din gud lever, o Dan», och: »Så sant den lever, som man dyrkar i Beer-Seba.»
De skola falla och icke mer stå upp.
Jag såg HERREN stå invid altaret, och han sade: Slå till pelarhuvudena, så att trösklarna bäva, och låt spillrorna falla över huvudet på alla där.
Deras sista kvarleva skall jag sedan dräpa med svärd.
Ingen av dem skall kunna undfly, ingen av dem kunna rädda sig.
Om de än bröte sig in i dödsriket, så skulle min hand hämta dem fram därifrån; och fore de än upp till himmelen, så skulle jag störta dem ned därifrån.
Gömde de sig än på toppen av Karmel, så skulle jag där leta fram dem och hämta dem ned; och dolde de sig än undan min åsyn på havets botten, så skulle jag där mana ormen fram att stinga dem.
Om de läte föra sig bort i fångenskap av sina fiender, skulle jag bjuda svärdet att där komma och dräpa dem.
Ja, jag skall låta mitt öga vila på dem, till deras olycka och icke till deras lycka.
Ty Herren, HERREN Sebaot, han som rör vid jorden, då försmälter den av ångest och alla dess inbyggare sörja, ja, hela jorden höjer sig såsom Nilen och sjunker åter såsom Egyptens flod;
han som bygger sin sal i himmelen och befäster sitt valv över jorden, han som kallar på havets vatten och gjuter det ut över jorden -- HERREN är hans namn.
Ären I icke för mig lika med etiopiernas barn, I Israels barn? säger HERREN.
Förde jag icke Israel upp ur Egyptens land och filistéerna ifrån Kaftor och araméerna ifrån Kir?
Se, Herrens, HERRENS ögon äro vända mot detta syndiga rike, och jag skall förgöra det från jordens yta.
Dock vill jag icke alldeles förgöra Jakobs hus, säger HERREN.
Ty se, jag skall låta ett bud utgå, att Israels hus må bliva siktat bland alla hednafolken, såsom siktades det i ett såll; icke det minsta korn skall falla på jorden.
Alla syndare i mitt folk skola dö för svärdet, de som nu säga: »Oss skall olyckan ej nalkas, över oss skall den icke komma.»
På den dagen skall jag upprätta Davids förfallna hydda; jag skall mura igen dess revor och upprätta dess ruiner och bygga upp den, sådan den var i forna dagar;
så att de få taga i besittning vad som är kvar av Edom och av alla hedningar som hava uppkallats efter mitt namn, säger HERREN, han som skall göra detta.
Se, dagar skola komma, säger HERREN, då plöjaren skall följa skördemannen i spåren, och druvtramparen såningsmannen, då bergen skola drypa av druvsaft och alla höjder skola försmälta.
Då skall jag åter upprätta mitt folk Israel; när de bygga upp sina ödelagda städer, skola de ock få bo i dem; när de plantera vingårdar, skola de ock få dricka vin från dem; när de anlägga trädgårdar, skola de ock få äta deras frukt.
Jag skall då plantera dem i deras eget land, och de skola icke mer ryckas upp ur det land som jag har givit dem, säger HERREN, din Gud.
Detta är Obadjas syn.
Så säger Herren, HERREN om Edom: Ett budskap hava vi hört från HERREN, och en budbärare är utsänd bland folken: »Upp, ja, låt oss stå upp och strida mot det!»
Se, jag skall göra dig ringa bland folken, djupt föraktad skall du bliva.
Ditt hjärtas övermod har bedragit dig, där du sitter ibland bergsklyftorna i den höga boning och säger i ditt hjärta: »Vem kan störta mig ned till jorden?»
Om du än byggde ditt näste så högt uppe som örnen, ja, om det än bleve förlagt mitt ibland stjärnorna, så skulle jag dock störta dig ned därifrån, säger HERREN.
När tjuvar komma över dig, och rövare om natten, ja då är det förbi med dig.
Sannerligen, de skola stjäla så mycket dem lyster.
När vinbärgare komma över dig, sannerligen, en ringa efterskörd skola de lämna kvar.
Huru genomsökt skall icke Esau bliva, huru skola ej hans dolda skatter letas fram!
Ut till gränsen skola de driva dig, alla dina bundsförvanter; dina vänner skola svika dig och skola taga väldet över dig.
I stället för att giva dig bröd skola de lägga en snara på din väg, där du icke kan märka den.
Sannerligen, på den dagen, säger HERREN skall jag förgöra de vise i Edom och allt förstånd på Esaus berg.
Dina hjältar, o Teman, skola då bliva slagna av förfäran; och så skall var man på Esaus berg bliva utrotad och dräpt.
Ja, för det våld du övade mot din broder Jakob skall du höljas med skam och bliva utrotad till evig tid.
På den dag då du lämnade honom i sticket, på den dag då främlingar förde bort hans gods och utlänningar drogo in genom hans port och kastade lott om Jerusalem, då var ju ock du såsom en av dem.
Men se icke så med lust på din broders dag, på hans motgångs dag; gläd dig icke så över Juda barn på deras undergångs dag; spärra icke upp munnen så stort på nödens dag.
Drag icke in genom mitt folks port på deras ofärds dag; se ej så hans olycka med lust, också du, på hans ofärds dag; och räck icke ut din hand efter hans gods på hans ofärds dag.
Ställ dig icke vid vägskälet för att nedgöra hans flyktingar, och giv icke hans undsluppna till pris på nödens dag.
Ty HERRENS dag är nära för alla hednafolk.
Såsom du har gjort, så skall man ock göra mot dig; dina gärningar skola komma tillbaka över ditt eget huvud.
Ja, såsom I haven druckit på mitt heliga berg, så skola ock alla hednafolk få dricka beständigt, de skola få dricka kalken i botten och bliva såsom hade de ej varit till.
Men på Sions berg skall finnas en räddad skara, och det skall vara en helig plats; och Jakobs hus skall åter få råda över sina besittningar.
Då skall Jakobs hus bliva en eld och Josefs hus en låga, och Esaus hus skall varda såsom strå, och de skola antända det och förtära det, och ingen skall slippa undan av Esaus hus; ty så har HERREN talat.
Och Sydlandets folk skall taga Esaus berg i besittning, och Låglandets folk skall taga filistéernas land; ja, också Efraims mark skall man taga i besittning, så ock Samariens mark.
Och Benjamin skall taga Gilead.
Och de bortförda av denna Israels barns här, de som bo i Kanaan allt intill Sarefat, så ock de bortförda från Jerusalem, de som leva i Sefarad, dessa skola taga Sydlandets städer i besittning.
Och frälsare skola draga upp på Sions berg till att döma Esaus berg.
Och så skall riket vara HERRENS.
Och HERRENS ord kom till Jona, Amittais son; han sade:
»Stå upp och begiv dig till Nineve, den stora staden, och predika för den; ty deras ondska har kommit upp inför mitt ansikte.»
Men Jona stod upp och ville fly till Tarsis, undan HERRENS ansikte.
Och han for ned till Jafo och fann där ett skepp som skulle gå till Tarsis.
Och sedan han hade erlagt betalning för resan, steg han ombord därpå för att fara med till Tarsis, undan HERRENS ansikte.
Men HERREN sände en stark vind ut över havet, så att en stark storm uppstod på havet; och skeppet var nära att krossas.
Då betogos sjömännen av fruktan och ropade var och en till sin gud; och vad löst som fanns i skeppet kastade de i havet för att bereda sig lättnad.
Men Jona hade gått ned i det inre av fartyget och låg där i djup sömn.
Då gick skepparen till honom och sade till honom: »Huru kan du sova så?
Stå upp och åkalla din Gud.
Kanhända skall den Guden tänka på oss, så att vi icke förgås.»
Och folket sade till varandra: »Välan, låt oss kasta lott, så att vi få veta för vems skull denna olycka har kommit över oss.»
När de så kastade lott, föll lotten på Jona.
Då sade de till honom: »Säg oss för vems skull denna olycka har kommit över oss.
Vad är ditt ärende, och varifrån kommer du?
Från vilket land och av vad folk är du?»
Han svarade den; »Jag är en hebré, och jag dyrkar HERREN, himmelens Gud, som har gjort havet och det torra.»
Då betogos männen av stor fruktan och sade till honom: »Vad är det du har gjort!»
Ty männen fingo genom det han berättade dem veta att han flydde undan HERRENS ansikte.
Och de sade till honom: »Vad skola vi göra med dig, så att havet stillar sig för oss?»
Ty havet stormade mer och mer.
Då svarade han dem: »Tagen mig och kasten mig i havet, så skall havet stillas för eder; ty jag vet att det är för min skull som denna starka storm har kommit över eder.»
Och männen strävade med all makt att komma tillbaka till land, men de kunde icke; ty havet stormade mer och mer emot dem.
Då ropade de till HERREN och sade: »Ack HERRE, låt oss icke förgås för denne mans själs skull, och låt icke oskyldigt blod komma över oss.
Ty du, HERRE, har gjort såsom dig täckes.»
Därefter togo de Jona och kastade honom i havet.
Då lade sig havets raseri.
Och männen betogos av stor fruktan för HERREN, och de offrade slaktoffer åt HERREN och gjorde löften.
Men HERREN sände en stor fisk, som slukade upp Jona.
Och Jona var i fiskens buk tre dagar och tre nätter.
Och Jona bad till HERREN, sin Gud, i fiskens buk.
Han sade: »Jag åkallade HERREN i min nöd, och han svarade mig; från dödsrikets buk ropade jag, och du hörde min röst.
Du kastade mig i djupet, mitt i havet, och strömmen omslöt mig, alla dina svallande böljor gingo över mig.
Jag tänkte då: 'Jag är bortdriven ifrån dina ögon.'
Men jag skall åter få skåda upp mot ditt heliga tempel.
Vatten omvärvde mig in på livet, djupet omslöt mig; sjögräs omsnärjde mitt huvud.
Till bergens grund sjönk jag ned, jordens bommar slöto sig bakom mig för evigt.
Men du förde min själ upp ur graven, HERRE, min Gud.
När min själ försmäktade i mig, då tänkte jag på HERREN, och min bön kom till dig, i ditt heliga tempel.
De som hålla sig till fåfängliga avgudar, de låta sin nåds Gud fara.
Men jag vill offra åt dig, med högljudd tacksägelse; vad jag har lovat vill jag infria; frälsningen är hos HERREN!»
Och på HERRENS befallning kastade fisken upp Jona på land.
Och HERRENS ord kom för andra gången till Jona; han sade:
»Stå upp och begiv dig till Nineve, den stora staden, och predika för den vad jag skall tala till dig.»
Då stod Jona upp och begav sig till Nineve, såsom HERREN hade befallt.
Men Nineve var en stor stad inför Gud, tre dagsresor lång.
Och Jona begav sig på väg in i staden, en dagsresa, och predikade och sade: »Det dröjer ännu fyrtio dagar, så skall Nineve bliva omstörtat.»
Då trodde folket i Nineve på Gud, och lyste ut en fasta och klädde sig i sorgdräkt, både stora och små.
Och när saken kom för konungen i Nineve, stod han upp från sin tron och lade av sin mantel och höljde sig i sorgdräkt och satte sig i aska.
Sedan utropade och förkunnade man i Nineve, enligt konungens och hans stores påbud, och sade: »Ingen människa må smaka något, icke heller något djur, vare sig av fäkreaturen eller småboskapen; de må icke föras i bet, ej heller vattnas.
Och både människor och djur skola hölja sig i sorgdräkt och ropa till Gud med all makt.
Och var och en må vända om från sin onda väg och från den orätt som han har haft för händer.
Vem vet, kanhända vänder Gud då om och ångrar sig och vänder sig ifrån sin vredes glöd, så att vi icke förgås.»
Då nu Gud såg vad de gjorde, att de vände om från sin onda väg, ångrade han det onda som han hade hotat att göra mot dem, och han gjorde icke så.
Men detta förtröt Jona högeligen, och hans vrede upptändes.
Och han bad till HERREN och sade: »Ack Herre, var det icke detta jag tänkte, när jag ännu var i mitt land!
Därför ville jag ock i förväg fly undan till Tarsis.
Jag visste ju att du är en nådig och barmhärtig Gud, långmodig och stor i mildhet, och sådan att du ångrar det onda.
Så tag nu, Herre, mitt liv ifrån mig; ty jag vill hellre vara död än leva.»
Men HERREN sade: »Menar du att du har skäl till att vredgas?»
Och Jona gick ut ur staden och stannade öster om staden; där gjorde han sig en hydda och satt i skuggan därunder, för att se huru det skulle gå med staden.
Och HERREN Gud lät en ricinbuske skjuta upp över Jona, för att den skulle giva skugga åt hans huvud och hjälpa honom ur hans förtrytelse; och Jona gladde sig högeligen över ricinbusken.
Men dagen därefter, när morgonrodnaden gick upp, sände Gud maskar som frätte ricinbusken, så att den vissnade.
När sedan solen hade gått upp, sände Gud en brännande östanvind, och solen stack Jona på huvudet, så att han försmäktade.
Då önskade han sig döden och sade: »Jag vill hellre vara död än leva.»
Men Gud sade till Jona: »Menar du att du har skäl till att vredgas för ricinbuskens skull?»
Han svarade: »Jag må väl hava skäl att vredgas till döds.»
Då sade HERREN: »Du ömkar dig över ricinbusken, som du icke har haft någon möda med och icke har dragit upp, som kom till på en natt och förgicks efter en natt.
Och jag skulle icke ömka mig över Nineve, den stora staden, där mer än ett hundra tjugu tusen människor finnas, som icke förstå att skilja mellan höger och vänster, och därtill djur i myckenhet!»
Detta är HERRENS ord som kom till morastiten Mika i Jotams, Ahas' och Hiskias, Juda konungars, tid, vad han skådade angående Samaria och Jerusalem.
Hören, I folk, allasammans; akta härpå, du jord med allt vad på dig är.
Och vare Herren, HERREN ett vittne mot eder, Herren i sitt heliga tempel.
Ty se, HERREN träder ut ur sin boning, han far ned och går fram över jordens höjder.
Bergen smälta under hans fötter, och dalar bryta sig fram -- såsom vaxet gör för elden, såsom vattnet, när det störtar utför branten.
Genom Jakobs överträdelse sker allt detta och genom Israels hus' synder.
Vem är då upphovet till Jakobs överträdelse?
Är det icke Samaria?
Och vem till Juda offerhöjder?
Är det icke Jerusalem?
Så skall jag då göra Samaria till en stenhop på marken, till en plats för vingårdsplanteringar; jag skall vräka hennes stenar ned i dalen, och hennes grundvalar skall jag blotta.
Alla hennes beläten skola bliva krossade, alla hennes skökoskänker uppbrända i eld, alla hennes avgudar skall jag förstöra; ty av skökolön har hon hopsamlat dem, och skökolön skola de åter bliva.
Fördenskull måste jag klaga och jämra mig, jag måste gå barfota och naken; jag måste upphäva klagoskri såsom en schakal och sorgelåt såsom en struts.
Ty ohelbara äro hennes sår; slaget har nått ända till Juda, det har drabbat ända till mitt folks port, ända till Jerusalem.
Förkunnen det icke i Gat; gråten icke så bittert.
I Bet-Leafra vältrar jag mig i stoftet.
Dragen åstad, I Safirs invånare, i nakenhet och skam.
Saanans invånare våga sig icke ut.
Klagolåten i Bet-Haesel tillstädjer eder ej att dröja där.
Ty Marots invånare våndas efter tröst; ned ifrån HERREN har ju en olycka kommit, intill Jerusalems port.
Spännen travare för vagnen, I Lakis' invånare, I som voren upphovet till dottern Sions synd; ty hos eder var det som Israels överträdelser först funnos.
Därför måste du giva skiljebrev åt Moreset-Gat.
Husen i Aksib hava för Israels konungar blivit såsom en försinande bäck.
Ännu en gång skall jag låta erövraren komma över eder, I Maresas invånare.
Ända till Adullam skall Israels härlighet komma.
Raka dig skallig och skär av ditt hår, i sorg över barnen, som voro din lust; gör ditt huvud så kalt som gamens, ty de skola föras bort ifrån dig.
Ve dessa som tänka ut vad fördärvligt är och bereda vad ont är på sina läger, och som sätta det i verket, så snart morgonen gryr, allenast det står i deras makt;
dessa som hava begärelse till sin nästas åkrar och röva dem, eller till hans hus och tillägna sig dem; dessa som öva våld mot både människor och hus, mot både ägare och egendom!
Därför säger HERREN så: Se, jag tänker ut mot detta släkte vad ont är; och I skolen icke kunna draga eder hals därur, ej heller skolen I sedan gå så stolta, ty det bliver en ond tid.
På den dagen skall man stämma upp en visa över eder och sjunga en sorgesång; man skall säga: »Det är ute med oss, vi äro förstörda i grund!
Mitt folks arvslott bliver nu given åt en annan.
Ja i sanning, den ryckes ifrån mig, och åt avfällingar utskiftas våra åkrar.»
Så sker det att hos dig icke mer finnes någon som får spänna mätsnöre över en lott i HERRENS församling.
»Hören då upp att predika», så är deras predikan; »om sådant får man icke predika; det är ju ingen ände på smädelser!»
Är detta ett tillbörligt tal, du Jakobs hus?
Har då HERREN varit snar till vrede?
Hava hans gärningar visat något sådant?
Äro icke fastmer mina ord milda mot den som vandrar redligt?
Men nu sedan en tid uppreser sig mitt folk såsom en fiende.
I sliten manteln bort ifrån kläderna på människor som trygga gå sin väg fram och ej vilja veta av strid.
Mitt folks kvinnor driven I ut från de hem där de hade sin lust; deras barn beröven I för alltid den berömmelse de hade av mig.
Stån upp och gån eder väg!
Här skolen I icke hava någon vilostad, för eder orenhets skull, som drager i fördärv, ja, i gruvligt fördärv.
Om någon som fore med munväder och falskhet sade i sin lögnaktighet: »Jag vill predika för dig om vin och starka drycker» -- det vore en predikare för detta folk!
Jag vill församla dig, Jakob, ja, hela ditt folk.
Jag vill hämta tillhopa Israels kvarlevor, jag vill föra dem tillsammans såsom fåren till fållan, såsom en hjord till dess betesmark, så att där uppstår ett gny av människor.
En vägbrytare drager ut framför dem; de bryta sig igenom och tåga fram, genom porten vandra de ut.
Deras konung tågar framför dem, HERREN går i spetsen för dem.
Och jag sade: Hören, I Jakobs hövdingar och I furstar av Israels hus.
Tillkommer det ej eder att veta vad rätt är,
I som haten det goda och älsken det onda, I som sliten huden av kroppen på människorna och köttet från deras ben?
Men eftersom dessa äta mitt folks kött och riva huden av deras kropp och bryta sönder deras ben, för att stycka dem likasom det man kastar i grytan, ja, likasom kött som lägges i kitteln,
därför skall HERREN icke svara dem, när de ropa till honom; han skall dölja sitt ansikte för dem på den tiden, för deras onda väsendes skull.
Så talar HERREN mot de profeter som föra mitt folk vilse, mot dem som ropa: »Allt står väl till!», så länge de hava något att tugga med sina tänder, men båda upp folket till helig strid mot den som ej giver dem något i gapet.
Därför skall natt komma över eder, så att det bliver slut på edra syner, och mörker, så att det bliver slut på edra spådomar.
Ja, solen skall gå ned över profeterna och dagen varda mörk över dem.
Siarna skola stå där med skam, och spåmännen skola få blygas; de skola alla nödgas skyla sitt skägg, då nu intet svar mer kommer från Gud.
Men jag, jag är uppfylld med kraft, ja, med HERRENS Ande, med rättsinne och frimodighet, så att jag kan förkunna för Jakob hans överträdelse och för Israel hans synd.
Hören då detta, I hövdingar av Jakobs hus och I furstar av Israels hus, I som hållen för styggelse vad rätt är och gören krokigt allt vad rakt är,
I som byggen upp Sion med blodsdåd och Jerusalem med orättfärdighet --
den stad vars hövdingar döma för mutor, vars präster undervisa för betalning, och vars profeter spå för penningar, allt under det de stödja sig på HERREN och säga: »Är icke HERREN mitt ibland oss?
Olycka skall ej komma över oss.»
Därför skall för eder skull Sion varda upplöjt till en åker och Jerusalem bliva en stenhop och tempelberget en skogbevuxen höjd.
Men det skall ske i kommande dagar att det berg där HERRENS hus är skall stå där fast grundat, ypperst ibland bergen, och vara upphöjt över andra höjder; och folk skall strömma ditupp,
ja, många hednafolk skola gå åstad och skola säga: »Upp, låt oss draga åstad till HERRENS berg, upp till Jakobs Guds hus, för att han må undervisa oss om sina vägar, så att vi kunna vandra på hans stigar.»
Ty från Sion skall lag utgå, och HERRENS ord från Jerusalem.
Och han skall döma mellan många folk och skipa rätt åt mäktiga hednafolk, ända bort i fjärran land.
Då skola de smida sina svärd till plogbillar och sina spjut till vingårdsknivar.
Folken skola ej mer lyfta svärd mot varandra och icke mer lära sig att strida.
Och var och en skall sitta under sitt vinträd och sitt fikonträd, och ingen skall förskräcka honom; ty så har HERREN Sebaots mun talat.
Ja, alla andra folk vandra vart och ett i sin guds namn, men vi vilja vandra i HERRENS, vår Guds, namn, alltid och evinnerligen.
På den dagen, säger HERREN, skall jag församla de haltande och hämta tillhopa de fördrivna och dem som jag har hemsökt med olyckor.
Och jag skall låta de haltande bliva en kvarleva och de långt bort förjagade ett mäktigt folk; och HERREN skall vara konung över dem på Sions berg från nu och till evig tid.
Och du Herdetorn, du dotter Sions kulle, till dig skall det komma, ja, till dig skall det återvända, det forna herradömet, dottern Jerusalems konungavälde.
Men varför skriar du nu så högt?
Finnes då ingen konung i dig, har du icke mer någon rådklok man, eftersom ångest, lik en barnaföderskas, har gripit dig?
Ja, väl må du vrida dig i födslosmärtor såsom en barnaföderska, du dotter Sion; ty nu måste du ut ur staden, du måste bo på öppna fältet; ja, du skall komma ända till Babel -- där skall du finna räddning, där skall HERREN förlossa dig ur dina fienders hand.
Nu hava många hednafolk församlat sig mot dig, och de säga: »Må hon varda skändad, så att våra ögon få skåda med lust på Sion.»
Men dessa känna icke HERRENS tankar, de förstå icke hans rådslut, att han har samlat dem såsom kärvar till tröskplatsen.
Upp då och tröska, du dotter Sion!
Ty jag skall giva dig horn av järn och giva dig klövar av koppar, för att du må sönderkrossa många folk.
Och deras byte skall du giva till spillo åt HERREN och deras skatter åt hela jordens HERRE.
Nu må du samla dina skaror, du skarornas stad.
Bålverk har man rest upp mot oss; Israels domare slår man med ris på kinden.
Men du Bet-Lehem Efrata, som är så ringa för att vara bland Juda släkter, av dig skall åt mig utgå en som skall bliva en furste i Israel, en vilkens härkomst tillhör förgångna åldrar, forntidens dagar.
Därför skola de prisgivas intill den tid då hon som skall föda har fött; då skall återstoden av hans bröder få vända tillbaka till Israels barn.
Och han skall träda fram och vakta sin hjord i HERRENS kraft, i HERRENS, sin Guds, namns höghet; och den skall hava ro, ty han skall då vara stor intill jordens ändar.
Och tryggheten skall vara sådan, att om Assur vill falla in i vårt land och tränga in i våra palats, så kunna vi ställa upp mot honom sju herdar, ja, åtta furstliga herrar;
och dessa skola avbeta Assurs land med svärd och Nimrods land ända in i dess portar.
Så skall han rädda oss från Assur, om denne vill falla in i vårt land och tränga fram över våra gränser.
Då skall Jakobs kvarleva vara bland många folk såsom dagg från HERREN, såsom en regnskur på gräs, vilken icke dröjer för någon mans skull eller väntar för människobarns skull.
Och Jakobs kvarleva skall då vara bland hedningarna, mitt ibland många folk, såsom ett lejon bland boskap i skogen, såsom ett ungt lejon bland fårhjordar, vilket förtrampar, var det går fram, och griper sitt rov utan räddning.
Ja, må din hand vara upplyft över dina ovänner, och må alla dina fiender bliva utrotade!
Och det skall ske på den dagen, säger HERREN, att jag skall utrota dina hästar ur ditt land och förstöra dina vagnar;
jag skall utrota städerna i ditt land och riva ned alla dina fästen;
jag skall utrota all trolldom hos dig, och inga teckentydare skola mer träffas hos dig;
jag skall utrota dina beläten och dina stoder ur ditt land, så att du icke mer skall tillbedja dina händers verk;
jag skall omstörta dina Aseror och skaffa dem bort ur ditt land; och dina städer skall jag ödelägga.
Och i vrede och förtörnelse skall jag utkräva hämnd av hednafolken, dem som icke hava varit hörsamma.
Hören vad HERREN säger: Stå upp och utför din sak inför bergen, och låt höjderna höra din röst.
Ja, hören HERRENS sak, I berg och I fasta klippor, jordens grundvalar!
Ty HERREN har sak mot sitt folk, och med Israel vill han gå till rätta.
Mitt folk, vad har jag gjort mot dig, och varmed har jag betungat dig?
Svara mig!
Jag förde dig ju upp ur Egyptens land, och ur träldomshuset förlossade jag dig; och Mose, Aron och Mirjam lät jag gå framför dig.
Mitt folk, kom ihåg vad Balak, konungen i Moab, hade i sinnet, och vad Bileam, Beors son, svarade honom; kom ihåg huru det var mellan Sittim och Gilgal, och lär dig så förstå HERRENS rättfärdighets gärningar.
Varmed skall jag träda fram inför HERREN, och varmed böja mig ned inför Gud i höjden?
Skall jag träda fram inför honom med brännoffer, med årsgamla kalvar?
Har HERREN behag till vädurar i tusental, till oljeströmmar i tiotusental?
Skall jag giva min förstfödde till offer för min överträdelse, min livsfrukt till syndoffer för min själ?
Nej, vad gott är har han kungjort för dig, o människa.
Ty vad annat begär HERREN av dig, än att du gör vad rätt är och vinnlägger dig om kärlek och vandrar i ödmjukhet inför din Gud?
Hör huru HERREN ropar till staden!
Ja, säll är den som aktar på ditt namn.
Hören om straffet, och vem han är, som har bestämt det.
Kunna ogudaktighetens skatter framgent få stanna i den ogudaktiges hus?
Kan där få finnas ett undermåligt efa-mått, värt att förbannas?
Vore jag rättfärdig, om jag fördroge orätt våg och falska vikter i pungen,
om de rika i staden finge vara fulla av orättrådighet, om dess invånare finge tala lögn och hava falsk tunga i sin mun?
Nej, och därför måste jag slå dig med oläkliga sår, hemsöka dig med förödelse för dina synders skull.
När du äter något, skall du icke bliva mätt, och tomhet skall råda i din buk.
Vad du skaffar undan skall du ändå icke kunna rädda, och vad du räddar skall jag giva åt svärdet.
Du skall så, men icke få skörda; du skall pressa oliver, men icke få smörja din kropp med oljan, du skall pressa ut druvmust, men icke få dricka vinet.
Vid Omris stadgar håller man fast, man efterföljer alla Ahabs hus' gärningar; ty efter dessas rådslag är det I vandren.
Därför skall jag göra dig till ett föremål för häpnad, och invånarna i staden till ett mål för begabberi; ja, mitt folks smälek skolen I få bära.
Ve mig!
Det är mig, såsom när frukten är insamlad om sommaren, eller såsom när efterskörden efter vinbärgningen är slut och ingen druvklase mer finnes att äta, intet förstlingsfikon av dem jag hade haft lust till.
De fromma äro försvunna ur landet, och ingen redlig man finnes bland människorna.
Alla ligga de på lur efter blod; envar vill fånga den andre i sitt nät.
Till att främja det onda äro deras händer redo: fursten begär gåvor, och domaren står efter vinning; den mäktige kräver öppet vad honom lyster; så bedriva de vrånghet.
Den bäste ibland dem är såsom ett törnsnår, den redligaste värre än en taggig häck.
Men när dina siares dag är inne, ja, när hemsökelsen når dig, då skall bestörtning komma ibland dem.
Man får icke tro på någon vän, icke lita på någon förtrogen; för henne som vilar i din famn måste du vakta din muns dörrar.
Ty sonen föraktar sin fader, dottern sätter sig upp mot sin moder, sonhustrun mot sin svärmoder, och envar har sitt eget husfolk till fiender.
Men jag vill skåda efter HERREN, jag vill hoppas på min frälsnings Gud; min Gud skall höra mig.
Glädjens icke över mig, I mina fiender.
Om jag än har fallit, skall jag dock stå upp igen; om jag än sitter i mörkret, är dock HERREN mitt ljus.
Eftersom jag har syndat mot HERREN, vill jag bära hans vrede, till dess att han utför min sak och skaffar mig rätt, till dess att han för mig ut i ljuset, så att jag med lust får se på hans rättfärdighet.
När mina fiender se det, skola de höljas med skam, desamma som säga till mig: »Var är nu HERREN, din Gud?»
Mina ögon skola se med lust på dem; ty då skola de bliva nedtrampade såsom orenlighet på gatan.
En dag skall komma, då dina murar skola byggas upp; på den dagen skola dina gränser sträcka sig vida.
På den dagen skall man komma till dig både från Assur och från Egyptens städer, ja från Egypten och ända ifrån floden, och från hav till hav, och från berg till berg.
Men eljest skall jorden bliva en ödemark för sina inbyggares skull; det skall vara deras gärningars frukt.
Vakta med din stav ditt folk, din arvedels hjord, så att den får hava sin avskilda boning i skogen på Karmel; låt den gå i bet i Basan och i Gilead, likasom under forna dagar.
Ja, likasom i de dagar då du drog ut ur Egyptens land skall jag låta dem se underbara ting.
Hedningarna skola se det och komma på skam med all sin makt.
De skola nödgas lägga handen på munnen, deras öron skola vara bedövade.
De skola slicka stoftet såsom ormar; lika maskar som kräla på jorden skola de med bävan övergiva sina borgar.
Med förskräckelse skola de söka HERREN, vår Gud; Ja, för dig skola de frukta.
Vem är en sådan Gud som du? -- du som förlåter kvarlevan av din arvedel dess missgärning och tillgiver den dess överträdelse, du som icke behåller vrede evinnerligen, ty du har lust till nåd,
och du skall åter förbarma dig över oss och trampa våra missgärningar under fötterna.
Ja, du skall kasta alla deras synder i havets djup.
Du skall bevisa trofasthet mot Jakob och nåd mot Abraham, såsom du med ed har lovat våra fäder i forntidens dagar.
Detta är en utsaga om Nineve, den bok som innehåller elkositen Nahums syn.
HERREN är en nitälskande Gud och en hämnare, ja, en hämnare är HERREN, en som kan vredgas.
En hämnare är HERREN mot sina ovänner, vrede behåller han mot sina fiender.
HERREN är långmodig, men han är stor i kraft, och ingalunda låter han någon bliva ostraffad.
HERREN har sin väg i storm och oväder och molnen äro dammet efter hans fötter.
Han näpser havet och låter det uttorka och alla strömmar låter han sina bort.
Då försmäkta Basan och Karmel, Libanons grönska försmäktar.
Bergen bäva för honom, och höjderna försmälta av ångest.
Jorden röres upp för hans ansikte, jordens krets med alla som bo därpå.
Vem kan bestå för hans ogunst, och vem kan uthärda hans vrede glöd?
Hans förtörnelse utgjuter sig såsom eld, och klipporna rämna inför honom.
HERREN är god, ett värn i nödens tid, och han låter sig vårda om dem som förtrösta på honom.
Men genom en störtflod gör han ände på platsen där den staden står, och hans fiender förföljas av mörker.
Ja, på edert anslag mot HERREN gör han ände, icke två gånger behöver hemsökelsen drabba.
Ty om de ock äro hopslingrade såsom törnsnår och så fulla av livssaft, som deras dryck är av must, skola de likväl alla förbrännas såsom torrt strå.
Ty från dig drog ut en man som hade onda anslag mot HERREN, en vilkens rådslag voro fördärv.
Så säger HERREN: »Huru starka och huru många de ock må vara, skola de ändå mejas av och försvinna; och om jag förr har plågat dig, så skall jag nu ej göra det mer.
Ty nu skall jag bryta sönder de ok han har lagt på dig, och hans band skall jag slita av.»
Men om dig bjuder HERREN så »Ingen avkomma av ditt namn skall mer få finnas.
Ur dina gudars hus skall jag utrota alla beläten, både skurna och gjutna.
En grav bereder jag åt dig, ty på skam har du kommit.»
Se, över bergen nalkas glädjebudbärarens fötter hans som förkunnar frid: »Fira dina högtider, Juda, infria dina löften.
Ty ej mer skall fördärvaren draga fram mot dig; han varder förgjord i grund.»
En folkförskingrare drager upp mot dig; bevaka dina fästen.
Speja utåt vägen, omgjorda dina länder bruka din kraft, så mycket du förmår.
Ty HERREN vill återställa Jakobs höghet såsom Israels höghet, då nu plundrare så hava ödelagt dem och så fördärvat deras vinträd.
Hans hjältars sköldar äro färgade röda, stridsmännen gå klädda i scharlakan; vagnarna gnistra av eld, när han gör dem redo till strid; och man skakar lansar av cypressträ.
På vägarna storma vagnarna fram, de köra om varandra på fälten; såsom bloss äro de att skåda lika ljungeldar fara de åstad.
Han vet nogsamt vilka väldiga kämpar han äger; de störta överända, där de rusa framåt.
De hasta mot stadens murar, och stormtaken göras redo.
Strömportarna måste öppna sig, och palatset försmälter av ångest.
Ja, domen står fast: hon bliver blottad, bortsläpad; hennes tärnor måste sucka likasom duvor och slå sig för sitt bröst.
I all sin tid var Nineve lik en vattenrik damm, men nu flyr vattnet bort. »Stannen!
Stannen!» -- Nej, ingen vänder sig om.
Röven nu silver, röven guld.
Här finnas skatter utan ände, överflöd på alla dyrbara håvor.
Ödeläggelse och förödelse och förstörelse!
Förfärade hjärtan och skälvande knän!
Darrande länder allestädes!
Allas ansikten hava skiftat färg.
Var är nu lejonens kula, den plats där de unga lejonen förtärde sitt rov, där lejonet och lejoninnan hade sin gång, där lejonungen gick omkring, utan att någon skrämde bort den?
Var är lejonet som tog rov, så mycket dess ungar ville hava, och dödade åt sina lejoninnor, ja, uppfyllde sina hålor med rov och sina kulor med rövat gods?
Se, jag skall vända mig mot dig, säger HERREN Sebaot; dina vagnar skall jag låta gå upp i rök, och dina unga lejon skall svärdet förtära.
Jag skall utrota ditt rövade gods från jorden och man skall ej mer höra dina sändebuds röst
Ve dig, du blodstad, alltigenom så full av lögn och våld, du som aldrig upphör att röva!
Hör, piskor smälla!
Hör, vagnshjul dåna!
Hästar jaga fram, och vagnar rulla åstad.
Ryttare komma i fyrsprång; svärden ljunga, och spjuten blixtra.
Slagna ser man i mängd och lik i stora hopar; igen ände är på döda, man stupar över döda.
Allt detta för den myckna otukt hon bedrev, hon, den fagra och trollkunniga skökan, som prisgav folkslag genom sin otukt och folkstammar genom sina trolldomskonster.
Se, jag skall vända mig mot dig, säger HERREN Sebaot; jag skall lyfta upp ditt mantelsläp över ditt ansikte och låta folkslag se din blygd och konungariken din skam.
Och jag skall kasta på dig vad styggeligt är, jag skall låta dig bliva föraktad, ja, göra dig till ett skådespel.
Var och en som ser dig skall sky dig och skall säga: »Nineve är ödelagt, men vem kan ömka det?»
Ja, var finner man någon som vill trösta dig?
Är du då bättre än No-Amon, hon som tronade vid Nilens strömmar, omsluten av vatten -- ett havets fäste, som hade ett hav till mur?
Etiopier i mängd och egyptier utan ände, putéer och libyer voro dig till hjälp.
Också hon måste ju gå i landsflykt och fångenskap, också hennes barn blevo krossade i alla gathörn; om hennes ädlingar kastade man lott, och alla hennes stormän blevo fängslade med kedjor
Så skall ock du bliva drucken och sjunka i vanmakt; också du skall få leta efter något värn mot fienden.
Alla dina fästen likna fikonträd med brådmogen frukt: vid minsta skakning falla de i munnen på den som vill äta dem.
Se, ditt manskap är hos dig såsom kvinnor; ditt lands portar stå vidöppna för dina fiender; eld förtär dina bommar.
Hämta dig vatten till förråd under belägringen, förstärk dina fästen.
Stig ned i leran och trampa i murbruket; grip till tegelformen.
Bäst du står där, skall elden förtära dig och svärdet utrota dig.
Ja, såsom av gräsmaskar skall du bliva uppfrätt, om du ock själv samlar skaror så talrika som gräsmaskar, skaror så talrika som gräshoppor.
Om du ock har krämare flera än himmelens stjärnor, så vet: gräsmaskarna fälla sina vingars höljen och flyga bort.
Ja, dina furstar äro såsom gräshoppor och dina hövdingar såsom gräshoppssvärmar: de stanna inom murarna, så länge det är svalt, men när solen kommer fram, då fly de bort, och sedan vet ingen var de finnas.
Dina herdar hava slumrat in, du Assurs konung; dina väldige ligga i ro.
Ditt folk är förstrött uppe på bergen, och ingen församlar det.
Det finnes ingen bot för din skada oläkligt är ditt sår.
Alla som höra vad som har hänt dig klappa i händerna över dig.
Ty över vem gick ej din ondska beständigt?
Detta är den utsaga som uppenbarades för profeten Habackuk.
Huru länge, HERRE, skall jag ropa, utan att du hör klaga inför dig över våld, utan att du frälsar?
Varför låter du mig se sådan ondska?
Huru kan du själv skåda på sådan orättrådighet, på det fördärv och det våld jag har inför mina ögon?
Så uppstår ju kiv, och så upphäva sig trätor.
Därigenom bliver lagen vanmäktig, och rätten kommer aldrig fram.
Ty den ogudaktige snärjer den rättfärdige; så framstår rätten förvrängd.
Sen efter bland hedningarna och skåden; häpnen, ja, stån där med häpnad Ty en gärning utför han i edra dagar, som I icke skolen tro, när den förtäljes.
Ty se, jag skall uppväcka kaldéerna det bistra och oförvägna folket, som drager ut så vitt som jorden når och inkräktar boningar som icke äro deras.
Det folket är förskräckligt och fruktansvärt; rätt och myndighet tager det sig självt.
Dess hästar äro snabbare än pantrar och vildare än vargar om aftonen; dess ryttare jaga fram i fyrsprång.
Ja, fjärran ifrån komma dess ryttare, de flyga åstad såsom örnen, när han störtar sig över sitt rov
Alla hasta de till våld, av sin stridslust drivas de framåt; och fångar hopa de såsom sand.
Konungar äro dem ett åtlöje, och furstar räkna de för lekverk; åt alla slags fästen le de, de kasta upp jordvallar och intaga dem.
Så fara de åstad såsom vinden, alltjämt framåt till att åsamka sig skuld; ty deras egen kraft är deras gud.
Är du då icke till av ålder?
Jo, HERRE, min Gud, min Helige, vi skola ej dö!
HERRE, till en dom är det du har satt dem, och till en tuktan har du berett dem, du vår klippa.
Du vilkens ögon äro för rena för att se på det onda, du som icke lider att skåda på orättrådighet, huru kan du ändå skåda på dessa trolösa människor och tiga stilla, när den ogudaktige fördärvar den som har rätt mot honom?
Så vållar du att människorna bliva lika fiskar i havet, lika kräldjur, som icke hava någon herre.
Ja, denne drager dem allasammans upp med sin krok, han fångar dem i sitt nät och församlar dem i sitt garn; däröver är han glad och fröjdar sig.
Fördenskull frambär han offer åt sitt nät och tänder offereld åt sitt garn; genom dem bliver ju hans andel så fet och hans mat så kräslig.
Men skall han därför framgent få tömma sitt nät och beständigt dräpa folken utan någon förskoning
Jag vill stiga upp på min vaktpost och ställa mig på muren; jag vill speja för att se vad han skall tala genom mig, och vilket svar på mitt klagomål jag skall få att frambära.
Och HERREN svarade mig och sade: Skriv upp din syn, och uppteckna den på skrivtavlor, med tydlig skrift, så att den lätt kan läsas.
Ty ännu måste synen vänta på sin men den längtar efter fullbordan och skall icke slå fel.
Om den dröjer, så förbida den, ty den kommer förvisso, den skall ej utebliva.
Se, uppblåst och orättrådig är dennes själ i honom; men den rättfärdige skall leva genom sin tro.
Ty såsom vinet icke är att lita på, så skall denne övermodige ej bestå, om han ock spärrar upp sitt gap såsom dödsriket och är omättlig såsom döden, om han ock har församlat till sig alla folk och hämtat tillhopa till sig alla folkslag.
Sannerligen, de skola allasammans stämma upp en visa över honom, ja, en smädesång om honom med välbetänkta ord; man skall säga: Ve dig som hopar vad som icke är ditt och belastar dig med utpantat gods -- men för huru länge!
Sannerligen, oförtänkt skola borgenärer resa sig mot dig och anfäktare vakna upp mot dig, och du skall bliva ett byte för dem.
Såsom du själv har plundrat många folk, så skola ock alla andra folk få plundra dig, för dina blodsdåd mot människor och ditt våld mot länder, mot städer och alla som bo i dem.
Ve dig som söker orätt vinning åt ditt hus, för att kunna bygga ditt näste högt uppe och så skydda dig undan olyckans våld!
Med dina rådslag drager du skam över ditt hus, i det att du gör ände på många folk och så syndar mot dig själv.
Ty stenarna i muren skola ropa, och bjälkarna i trävirket skola svara dem.
Ve dig som bygger upp städer med blodsdåd och befäster orter med orättfärdighet!
Se, av HERREN Sebaot är det ju sagt: »Så möda sig folken för det som skall förbrännas av elden- och folkslagen arbeta sig trötta för det som skall bliva till intet.»
Ty jorden skall varda full av HERRENS härlighets kunskap, likasom havsdjupet är fyllt av vattnet.
Ve dig som iskänker vin åt din nästa och blandar ditt gift däri och berusar honom, för att få skåda hans blygd!
Med skam skall du få mätta dig i stället för med ära.
Ja, du skall också själv få dricka, till dess du ligger där med blottad förhud.
Kalken skall i sin ordning räckas dig av HERRENS hand, och smälek skall hölja din ära.
Ty över dig skall komma en hemsökelse, lik Libanons, och en förhärjelse, lik den som skrämmer bort dess djur, för dina blodsdåd mot människor och ditt våld mot länder, mot städer och alla som bo i dem.
Vad kan ett skuret beläte hjälpa, eftersom en snidare vill slöjda sådant?
Och vad ett gjutet beläte, en falsk vägvisare, eftersom dess formare så förtröstar därpå, att han gör sig stumma avgudar?
Ve dig som säger till stocken: »Vakna!», och till döda stenen: »Vakna upp!»
Kan en sådan giva någon vägvisning?
Visst är den överdragen med guld och silver, men alls ingen ande är däri.
Men HERREN är i sitt heliga tempel.
Hela jorden vare stilla inför honom.
En bön av profeten Habackuk; till Sigjonót.
HERRE, jag har hört om dig och häpnat.
HERRE, förnya i dessa år dina gärningar, låt oss förnimma dem i dessa år.
Mitt i din vrede må du tänka på förbarmande.
Gud kommer från Teman, den helige från berget Paran.
Sela.
Hans majestät övertäcker himmelen, och av hans lov är jorden full.
Då uppstår en glans såsom av solljus, strålar gå ut ifrån honom, och han höljer i dem sin makt.
Framför honom går pest, och feberglöd följer i hans spår.
Han träder fram -- därmed kommer han jorden att darra; en blick -- och han kommer folken att bäva.
De uråldriga bergen splittras, de eviga höjderna sjunka ned.
Han vandrar de vägar han fordom gick.
Jag ser Kusans hyddor hemsökta av fördärv; tälten darra i Midjans land.
Harmas då HERREN på strömmar?
Ja, är din vrede upptänd mot strömmarna eller din förgrymmelse mot havet, eftersom du så färdas fram med dina hästar, med dina segerrika vagnar?
Framtagen och blottad är din båge, ditt besvurna ords pilar.
Sela.
Till strömfåror klyver du jorden.
Bergen se dig och bäva; såsom en störtskur far vattnet ned.
Djupet låter höra sin röst, mot höjden lyfter det sina händer.
Sol och måne stanna i sin boning för skenet av dina farande pilar, för glansen av ditt blixtrande spjut.
I förgrymmelse går du fram över jorden, i vrede tröskar du sönder folken.
Du drager ut för att frälsa ditt folk, för att bereda frälsning åt din smorde.
Du krossar taket på de ogudaktigas hus, du bryter ned huset, från grunden till tinnarna.
Sela.
Du genomborrar deras styresmans huvud med hans egna pilar, när de storma fram till att förskingra oss, under fröjd, såsom gällde det att i lönndom äta upp en betryckt.
Du far med dina hästar fram över havet, över de stora vattnens svall.
Jag hör det och darrar i mitt innersta, vid dånet skälva mina läppar; maktlöshet griper benen i min kropp, jag darrar på platsen där jag står.
Ty jag måste ju stilla uthärda nödens tid, medan det kommer, som skall tränga folket.
Ja, fikonträdet blomstrar icke mer, och vinträden giva ingen skörd, olivträdets frukt slår fel och fälten alstra ingen äring, fåren ryckas bort ur fållorna, och inga oxar finnas mer i stallen.
Likväl vill jag glädja mig i HERREN och fröjda mig i min frälsnings Gud.
HERREN, Herren är min starkhet; han gör mina fötter såsom hindens och låter mig gå fram över mina höjder.
För sångmästaren, med mitt strängaspel.
Detta är HERRENS ord som kom till Sefanja, son till Kusi, son till Gedalja, son till Amarja, son till Hiskia, i Josias, Amons sons, Juda konungs, tid.
Jag skall rycka bort och förgöra allt vad på jorden är, säger HERREN;
jag skall förgöra människor och djur, jag skall förgöra fåglarna under himmelen och fiskarna i havet, det vacklande riket jämte de ogudaktiga människorna; ja, människorna skall jag utrota från jorden, säger HERREN.
Jag skall uträcka min hand mot Juda och mot Jerusalems alla invånare och utrota från denna plats Baals sista kvarleva, avgudaprofeternas namn jämte prästerna;
dem som på taken tillbedja himmelens härskara, och dem som tillbedja HERREN och svärja vid honom och svärja vid Malkam;
dem som hava vikit bort ifrån HERREN, och dem som aldrig hava sökt HERREN eller frågat efter honom.
Varen stilla inför Herren, HERREN!
Ty HERRENS dag är nära; HERREN har tillrett ett slaktoffer, han har invigt sina gäster.
Och det skall ske på HERRENS slaktoffers dag att jag skall hemsöka furstarna och konungasönerna och alla som kläda sig i utländska kläder;
Jag skall på den dagen hemsöka alla som hoppa över tröskeln, dem som fylla sin herres hus med våld och svek.
På den dagen, säger HERREN, skall klagorop höras ifrån Fiskporten och jämmer från Nya staden och stort brak från höjderna.
Jämren eder, I som bon i Mortelkvarteret, ty det är förbi med hela krämarskaran; utrotade äro alla de penninglastade.
Och det skall ske på den tiden att jag skall genomleta Jerusalem med lyktor och hemsöka de människor som nu ligga där i ro på sin drägg, dem som säga i sina hjärtan: »HERREN gör intet, varken gott eller ont.»
Deras ägodelar skola då lämnas till plundring och deras hus till ödeläggelse.
Om de bygga sig hus, skola de ej få bo i dem, och om de plantera vingårdar, skola de ej få dricka vin från dem.
HERRENS stora dag är nära, ja, den är nära, den kommer med stor hast.
Hör, det är HERRENS dag!
I ångest ropa nu hjältarna.
En vredens dag är den dagen, en dag av ångest och trångmål, en dag av ödeläggelse och förödelse en dag av mörker och tjocka, en dag av moln och töcken,
en dag då basunljud och härskri höjes mot de fastaste städer och mot de högsta murtorn.
Då skall jag bereda människorna sådan ångest att de gå där såsom blinda, därför att de hava syndat mot HERREN.
Deras blod skall spridas omkring såsom stoft, och deras kroppar skola kastas ut såsom orenlighet.
Varken deras silver eller deras guld skall kunna rädda dem på HERRENS vredes dag.
Av hans nitälskans eld skall hela jorden förtäras.
Ty en ände, ja, en ände med förskräckelse skall han göra på alla jordens inbyggare.
Besinna dig och kom till sans, du folk utan blygsel,
innan ännu rådslutet är fullgånget -- den dagen hastar fram, såsom agnar fara! -- och innan HERRENS vredes glöd kommer över eder, ja, innan HERRENS vredes dag kommer över eder.
Söken HERREN, alla I ödmjuke i landet, som hållen hans lag.
Söken rättfärdighet, söken ödmjukhet; kanhända bliven I så beskärmade på HERRENS vredes dag.
Ty Gasa skall bliva övergivet och Askelon varda en ödemark; mitt på ljusa dagen skall Asdods folk drivas ut, och Ekron skall ryckas upp med roten.
Ve eder som bebon landsträckan utmed havet, I av keretéernas folk!
Ett HERRENS ord skall nå dig, Kanaan, du filistéernas land; ja, jag skall fördärva dig, så att ingen mer bor i dig.
Och landsträckan utmed havet skall ligga såsom betesmarker, där herdarna hava sina brunnar och fåren sina fållor.
Och den skall tillfalla de kvarblivna av Juda hus såsom deras lott; där skola de föra sin boskap i bet.
I Askelons hus skola de få lägra sig, när aftonen kommer.
Ty HERREN, deras Gud, skall se till dem och skall åter upprätta dem.
Jag har hört Moabs smädelser och Ammons barns hån, huru de hava smädat mitt folk och förhävt sig mot dess land.
Därför, så sant jag lever, säger HERREN Sebaot, Israels Gud: det skall gå Moab såsom Sodom, och Ammons barn såsom Gomorra.
Ett tillhåll för nässlor och en saltgrop skola de bliva, och en ödemark till evig tid.
Kvarlevan av mitt folk skall plundra dem. och återstoden av min menighet skall få dem till sin arvedel.
Så skall det gå dem, till lön för deras högmod därför att de hava smädat och förhävt sig mot HERREN Sebaots folk.
Fruktansvärd skall HERREN bevisa sig mot dem; ty han skall göra alla jordens gudar maktlösa, och alla hedningarnas havsländer skola tillbedja honom, vart folk på sin ort --
också I etiopier, I som av mig bliven slagna med svärd.
Och han skall uträcka sin hand mot norr och fördärva Assur, han skall göra Nineve till en ödemark, förtorkat såsom en öken.
Och därinne skola hjordar lägra sig, allahanda vilda djur i skaror; pelikaner och rördrommar skola taga natthärbärge på pelarhuvudena därinne; fåglalåt skall ljuda i fönstren och förödelse bo på trösklarna, nu då cederpanelningen är bortriven.
Så skall det gå den glada staden, som satt så trygg, och som sade i sitt hjärta: »Jag och ingen annan!»
Huru har den icke blivit en ödemark, en lägerstad för vilda djur!
Alla som gå där fram skola vissla åt den och slå ihop händerna.
Ve henne, den gensträviga och befläckade staden, förtryckets stad!
Hon hör icke på någons röst, hon tager ej emot tuktan; på HERREN förtröstar hon icke, till sin Gud vill hon ej komma.
Furstarna därinne äro rytande lejon; hennes domare äro såsom vargar om aftonen, de spara intet till morgondagen.
Hennes profeter äro stortaliga trolösa män; hennes präster ohelga vad heligt är, de våldföra lagen.
HERREN är rättfärdig därinne, han gör intet orätt. var morgon låter han sin rätt gå fram i ljuset, den utebliver aldrig; men de orättfärdiga veta icke av någon skam.
Jag utrotade folkslag, deras murtorn blevo förstörda, deras gator gjorde jag öde, så att ingen mer gick där fram; deras städer blevo förhärjade, så att de lågo tomma på människor, blottade på invånare.
Jag tillsade henne att allenast frukta mig och taga emot tuktan; då skulle hennes boning undgå förstörelse, med allt vad jag hade givit i hennes vård.
Men i stället ävlades de att göra allt vad fördärvligt var.
Därför man I vänta på mig, säger HERREN, och på den dag jag står upp för att taga byte.
Ty mitt domslut är: jag skall församla folk och hämta tillhopa konungariken, för att utgjuta över dem min ogunst, all min vredes glöd; ty av min nitälskans eld skall hela jorden förtäras.
Se, då skall jag giva åt folken nya, renade läppar, så att de allasammans åkalla HERRENS namn och endräktigt tjäna honom.
Ända ifrån länderna bortom Etiopiens strömmar skola mina tillbedjare, mitt förskingrade folk, frambära offer åt mig.
På den tiden skall du slippa att längre blygas för alla de överträdelser som du har begått mot mig.
Ty då skall jag avskilja från dig dem som nu jubla så segerstolt i dig; och du skall då icke vidare förhäva dig på mitt heliga berg.
Men jag skall lämna kvar i dig ett folk, betryckt och armt; och de skola förtrösta på HERRENS namn.
Kvarlevan av Israel skall då icke mer göra något orätt, ej heller tala lögn, och i deras mun skall icke finnas en falsk tunga.
Ja, de skola få beta och ligga i ro, utan att någon förskräcker dem.
Jubla, du dotter Sion, höj glädjerop, du Israel; var glad och fröjda dig av allt hjärta, du dotter Jerusalem.
HERREN har avvänt straffdomarna ifrån dig, han har röjt din fiende ur vägen.
HERREN, som bor i dig, är Israels konung; du behöver ej mer frukta något ont.
På den tiden skall det sägas till Jerusalem; »Frukta icke, Sion låt ej modet falla.
HERREN, din Gud, bor i dig en hjälte som kan frälsa.
Han gläder sig över dig med lust, han tiger stilla i sin kärlek, han fröjdas över dig med jubel.»
Dem som med bedrövelse måste sakna högtiderna, dem skall jag då församla, dem som levde skilda från dig, du som själv bar smälekens börda.
Ty se, jag skall på den tiden utföra mitt verk på alla dina förtryckare. jag skall frälsa de haltande och hämta tillhopa de fördrivna, jag skall låta dem bliva ett ämne till lovsång och till berömmelse på hela jorden, där de voro så smädade.
På den tiden skall jag låta eder komma tillbaka ja, på den tiden skall jag hämta eder tillhopa.
Ty jag vill låta eder bliva ett ämne till berömmelse och till lovsång bland alla jordens folk, i det att jag åter upprättar eder, så att I sen det med egna ögon, säger HERREN.
I konung Darejaves' andra regeringsår, i sjätte månaden, på första dagen i månaden, kom HERRENS ord genom profeten Haggai Serubbabel, Sealtiels son, Juda ståthållare, och till översteprästen Josua, Josadaks son; han sade:
Så säger HERREN Sebaot: Detta folk säger: »Ännu är icke tiden kommen att gå till verket, tiden att HERRENS hus bygges upp.»
Men HERRENS ord kom genom profeten Haggai; han sade:
Är då tiden kommen för eder att själva bo i panelade hus, medan detta hus ligger öde?
Därför säger nu HERREN Sebaot så: Given akt på huru det går eder.
I sån mycket, men inbärgen litet; I äten, men fån icke nog för att bliva mätta; I dricken, men fån icke nog för att bliva glada; I tagen på eder kläder, men haven icke nog för att bliva varma.
Och den som får någon inkomst, han far den allenast för att lägga den i en söndrig pung.
Ja, så säger HERREN Sebaot: Given akt på huru det går eder.
Men dragen nu upp till bergen, hämten trävirke och byggen upp mitt hus, så vill jag hava behag därtill och bevisa mig härlig, säger HERREN.
I väntaden på mycket, men se, det blev litet, och när I förden det hem, då blåste jag på det.
Varför gick det så? säger HERREN Sebaot.
Jo, därför att mitt hus får ligga öde, under det att envar av eder hastar med sitt eget hus.
Fördenskull har himmelen ovan eder förhållit eder sin dagg och jorden förhållit sin gröda.
Och jag har bjudit torka komma över land och berg, och över säd, vin och olja och alla andra jordens alster, och över människor och djur, och över all frukt av edra händers arbete.
Och Serubbabel, Sealtiels son, och översteprästen Josua, Josadaks son med hela kvarlevan av folket lyssnade till HERRENS, sin Guds, röst och till profeten Haggais ord, eftersom HERREN, deras Gud, hade sänt honom; och folket fruktade för HERREN.
Då sade Haggai, HERRENS sändebud, efter HERRENS uppdrag, till folket så: »Jag är med eder, säger HERREN.»
Och HERREN uppväckte Serubbabels, Sealtiels sons, Juda ståthållares, ande och översteprästen Josuas, Josadaks sons, ande och allt det kvarblivna folkets ande, så att de gingo till verket och arbetade på HERREN Sebaots; sin Guds, hus.
Detta skedde på tjugufjärde dagen i sjätte månaden av konung Darejaves' andra regeringsår.
I sjunde månaden, på tjuguförsta dagen i månaden, kom HERRENS ord genom profeten Haggai han sade:
Säg till Serubbabel, Sealtiels son Juda ståthållare, och till översteprästen Josua, Josadaks son, och till kvarlevan av folket:
Leva icke ännu bland eder män kvar, som hava sett detta hus i dess forna härlighet?
Och hurudant sen I det nu vara?
Är det icke såsom intet i edra ögon?
Men var likväl nu frimodig, du Serubbabel, säger HERREN; och var frimodig, du överstepräst Josua, Josadaks son; och varen frimodiga och arbeten, alla I som hören till folket i landet, säger HERREN; ty jag är med eder, säger HERREN Sebaot.
Det förbund som jag slöt med eder, när I drogen ut ur Egypten, vill jag låta stå fast, och min Ande skall förbliva ibland eder; frukten icke.
Ty så säger HERREN Sebaot: Ännu en gång, inom en liten tid, skall jag komma himmelen och jorden, havet och det torra att bäva;
och alla hednafolk skall jag komma att bäva, och så skola dyrbara håvor från alla hednafolk föras hit; och jag skall fylla detta hus med härlighet, säger HERREN Sebaot.
Ty mitt är silvret, och mitt är guldet, säger HERREN Sebaot.
Den tillkommande härligheten hos detta hus skall bliva större än dess forna var, säger HERREN Sebaot; och på denna plats skall jag låta friden råda, säger HERREN Sebaot.
På tjugufjärde dagen i nionde månaden av Darejaves' andra regeringsår kom HERRENS ord till profeten Haggai; han sade:
Så säger HERREN Sebaot: Fråga prästerna om lag och säg:
»Om någon bär heligt kött i fliken av sin mantel och så med fliken kommer vid något bakat eller kokt, eller vid vin eller olja, eller vid något annat som man förtär, månne detta därigenom bliver heligt?»
Prästerna svarade och sade: »Nej.»
Åter frågade Haggai: »Om den som har blivit orenad genom en död kommer vid något av allt detta, månne det då bliver orenat?»
Prästerna svarade och sade: »Ja.»
Då tog Haggai till orda och sade: »Så är det med detta folk och så är det med detta släkte inför mig, säger HERREN, och så är det med allt deras händers verk: vad de där offra, det är orent.
Och given nu akt på huru det hittills har varit, före denna dag, och under tiden innan man ännu hade begynt lägga sten på sten till HERRENS tempel
huru härförinnan, om någon kom till en sädesskyl som skulle giva tjugu mått, den gav allenast tio, och huru, om någon kom till vinpressen för att ösa upp femtio kärl, den gav allenast tjugu.
Vid allt edra händers arbete slog jag eder säd med sot och rost och hagel, och likväl vänden I eder icke till mig, säger HERREN.
Given alltså akt på huru det hittills har varit, före denna dag; ja, given akt på huru det har varit före tjugufjärde dagen i nionde månaden, denna dag då grunden har blivit lagd till HERRENS tempel.
Finnes någon säd ännu i kornboden?
Nej; och varken vinträdet eller fikonträdet eller granatträdet eller olivträdet har ännu burit någon frukt.
Men från denna dag skall jag giva välsignelse.»
Och HERRENS ord kom för andra gången till Haggai, på tjugufjärde dagen i samma månad; han sade:
Säg till Serubbabel, Juda ståthållare: Jag skall komma himmelen och jorden att bäva;
jag skall omstörta konungatroner och göra hednarikenas makt till intet; jag skall omstörta vagnarna med sina kämpar, och hästarna skola stupa med sina ryttare.
Den ene skall falla för den andres svärd.
På den tiden, säger HERREN Sebaot, skall jag taga dig, min tjänare Serubbabel, Sealtiels son, säger HERREN, och skall akta dig såsom min signetring; ty dig har jag utvalt, säger HERREN Sebaot.
I åttonde månaden av Darejaves' andra regeringsår kom HERRENS ord till Sakarja, son till Berekja, son till Iddo, profeten, han sade:
Svårt förtörnad var HERREN på edra fäder.
Säg därför nu till folket så säger HERREN Sebaot: Vänden om till mig, säger HERREN Sebaot, så vill jag vända om till eder, säger HERREN Sebaot.
Varen icke såsom edra fäder, för vilka forna tiders profeter predikade och sade: »Så säger HERREN Sebaot: Vänden om från edra onda vägar och edra onda gärningar»; men de ville icke höra och aktade icke på mig säger HERREN.
Edra fäder, var äro de?
Och profeterna, leva de kvar evinnerligen?
Nej, men mina ord och mina rådslut, de som jag betrodde åt mina tjänare profeterna, de träffade ju edra fäder, så att de måste vända om och säga: »Såsom HERREN Sebaot hade beslutit att göra med oss, och såsom våra vägar och våra gärningar förtjänade, så har han ock gjort med oss.»
På tjugufjärde dagen i elfte månaden, det är månaden Sebat, i Darejeves' andra regeringsår, kom HERRENS ord till Sakarja, son till Berekja, son till Iddo, profeten; han sade:
Jag hade en syn om natten: Jag fick se en man som red på en röd häst; och han höll stilla bland myrtenträden i dalsänkningen.
Och bakom honom stodo andra hästar, röda, bruna och vita.
Då frågade jag: »Vad betyda dessa, min herre?»
Ängeln som talade med mig svarade mig: »Jag vill låta dig förstå vad dessa betyda.»
Och mannen som stod bland myrtenträden tog till orda och sade: »Det är dessa som HERREN har sänt ut till att fara omkring på jorden.»
Och själva togo de till orda och sade till HERRENS ängel, som stod bland myrtenträden: »Vi hava farit omkring på jorden och hava funnit hela jorden lugn och stilla.»
Då tog HERRENS ängel åter till orda och sade: »HERRE Sebaot, huru länge skall det dröja, innan du förbarmar dig över Jerusalem och Juda städer?
Du har ju nu varit vred på dem i sjuttio år.»
Och HERREN svarade ängeln som talade med mig goda och tröstliga ord;
och ängeln som talade med mig sade sedan till mig: »Predika och säg: Så säger HERREN Sebaot: Jag har stor nitälskan för Jerusalem och Sion;
och jag är storligen förtörnad på hednafolken, som sitta så säkra; ty när jag var allenast litet förtörnad, hjälpte de ytterligare till att fördärva.
Därför säger HERREN så: Jag vill åter vända mig till Jerusalem i barmhärtighet; mitt hus skall där bliva uppbyggt, säger HERREN Sebaot, och mätsnöret skall spännas över Jerusalem.
Ytterligare må du predika och säga: Så säger HERREN Sebaot: Ännu en gång skola mina städer få njuta överflöd av goda håvor; ja, HERREN skall ännu en gång trösta Sion, och ännu en gång skall han utvälja Jerusalem.»
Sedan lyfte jag upp mina ögon och fick då se fyra horn.
Då frågade jag ängeln som talade med mig: »Vad betyda dessa?»
Han svarade mig: »Detta är de horn som hava förstrött Juda, Israel och Jerusalem.»
Sedan lät HERREN mig se fyra smeder.
Då frågade jag: »I vad ärende hava dessa kommit?»
Han svarade: »De förra voro de horn som förströdde Juda, så att ingen kunde upplyfta sitt huvud; men nu hava dessa kommit för att injaga skräck hos dem, och för att slå av hornen på de hednafolk som hava lyft sitt horn mot Juda land, till att förströ dess inbyggare.»
Sedan lyfte jag upp mina ögon och fick då se en man som hade ett mätsnöre i sin hand.
Då frågade jag: »Vart går du?»
Han svarade mig: »Till att mäta Jerusalem, för att se huru brett och huru långt det skall bliva.»
Då fick jag se ängeln som talade ned mig komma fram, och en annan ängel kom emot honom.
Och han sade till denne: »Skynda åstad och tala till den unge mannen där och säg: 'Jerusalem skall ligga såsom en obefäst plats; så stor myckenhet av människor och djur skall finnas därinne.
Men jag själv, säger HERREN, skall vara en eldsmur däromkring, och jag skall bevisa mig härlig därinne.'»
Upp, upp!
Flyn bort ur nordlandet, säger HERREN, I som av mig haven blivit förströdda åt himmelens fyra väderstreck, säger HERREN.
Upp, Sion!
Rädda dig, du som nu bor hos dottern Babel!
Ty så säger HERREN Sebaot, han som har sänt mig åstad för att förhärliga sig, så säger han om hednafolken, vilka plundrade eder (ty den som rör vid eder, han rör vid hans ögonsten):
»Se, jag lyfter min hand mot dem, och de skola bliva ett byte för sina forna trälar; och I skolen så förnimma att HERREN Sebaot har sänt mig.»
Jubla och gläd dig, du dotter Sion; ty se, jag kommer för att aga min boning i dig, säger HERREN.
Och då skola många hednafolk sluta sig till HERREN och bliva mitt folk.
Ja, jag skall taga min boning i dig; och du skall förnimma att HERREN Sebaot har sänt mig till dig.
Och HERREN skall hava Juda till I sin arvedel i det heliga landet, och ännu en gång skall han utvälja Jerusalem.
Allt kött vare stilla inför HERREN; ty han har stått upp och trätt fram ur sin heliga boning.
Sedan lät han mig se översteprästen Josua stående inför HERRENS ängel; och Åklagaren stod vid hans högra sida för att anklaga honom.
Men HERREN sade till Åklagaren: »HERREN skall näpsa dig, du Åklagare; ja, HERREN skall näpsa dig, han som har utvalt Jerusalem.
Är då icke denne en brand, ryckt ur elden?»
Och Josua var klädd i orena kläder, där han stod inför ängeln
Och denne tog till orda och sade till dem som stodo där såsom hans tjänare: »Tagen av honom de orena kläderna.»
Och till honom själv sade han: »Se, jag har tagit bort ifrån dig din missgärning, och man skall nu kläda dig i högtidskläder.»
Då sade jag: »Må man ock sätta en ren bindel på hans huvud.»
Och de satte en ren bindel på hans huvud och klädde på honom andra kläder, medan HERRENS ängel stod därbredvid.
Och HERRENS ängel betygade för Josua och sade:
»Så säger HERREN Sebaot: Om du vandrar på mina vägar och håller vad jag har bjudit dig hålla, så skall du ock få styra mitt hus och vakta mina gårdar; och jag skall låta dig hava din gång bland dessa som här göra tjänst.
Hör härpå, Josua, du överstepräst, med dina medbröder, som sitta här inför dig (ty dessa män skola vara ett tecken): Se, jag vill låta min tjänare Telningen komma;
ty se, i den sten som jag har lagt inför Josua -- över vilken ena sten sju ögon vaka -- i den skall jag inrista den inskrift som hör därtill, säger HERREN Sebaot; och jag skall utplåna detta lands missgärning på en enda dag.
På den tiden, säger HERREN Sebaot, skall var och en av eder kunna inbjuda den andre till gäst under sitt vinträd och fikonträd.»
Sedan blev jag av ängeln som talade med mig åter uppväckt, likasom när någon väckes ur sömnen.
Och han sade till mig: »Vad ser du?»
Jag svarade: »Jag ser en ljusstake, alltigenom av guld, med sin oljeskål ovantill och med sina sju lampor; och sju rör gå till de särskilda lamporna därovantill.
Och två olivträd sträcka sig över den, ett på högra sidan om skålen och ett på vänstra.»
Sedan frågade jag och sade till ängeln som talade med mig: »Vad betyda dessa ting, min herre?»
Men ängeln som talade med mig svarade och sade till mig: »Förstår du då icke vad de betyda?»
Jag svarade: »Nej, min herre.»
Då talade han och sade till mig: »Detta är HERRENS ord till Serubbabel: Icke genom någon människas styrka eller kraft skall det ske, utan genom min Ande, säger HERREN Sebaot.
Vilket du än må vara, du stora berg som reser dig mot Serubbabel, så skall du ändå förvandlas till jämn mark.
Ty han skall få föra fram slutstenen under jubelrop: 'Nåd, nåd må vila över den!'»
Vidare kom HERRENS ord till mig; han sade:
»Serubbabels händer hava lagt grunden till detta hus; hans händer skola ock få fullborda det.
Och du skall förnimma att HERREN Sebaot har sänt mig till eder.
Ty vem är den som vill förakta: den ringa begynnelsens dag, när dessa sju glädjas över att se murlodet i Serubbabels hand, dessa HERRENS ögon, som överfara hela jorden?»
Och jag frågade och sade till honom: »Vad betyda dessa två olivträd, det på högra och det på vänstra sidan om ljusstaken?»
Och ytterligare frågade jag och sade till honom: »Vad betyda de två olivkvistar som sträcka sig intill de två gyllene rännor genom vilka den gyllene oljan ledes ditned?»
Då sade han till mig: »Förstår du då icke vad de betyda?»
Jag svarade: »Nej, min herre.»
Då sade han: »Dessa äro de två oljesmorda som stå såsom tjänare inför hela jordens Herre.»
När jag sedan åter lyfte upp mina ögon, fick jag se en bokrulle flyga fram.
Och han sade till mig: »Vad ser du?»
Jag svarade: »Jag ser en bokrulle flyga fram; den är tjugu alnar lång och tio alnar bred.»
Då sade han till mig: »Detta är Förbannelsen, som går ut över hela landet; ty i kraft av den skall var och en som stjäl varda bortrensad härifrån, och i kraft av den skall var och en som svär varda bortrensad härifrån.
Jag har låtit den gå ut, säger HERREN Sebaot, för att den skall komma in i tjuvens hus och in i dens hus, som svär falskt vid mitt namn; och den skall stanna där i huset och fräta upp det med både trävirke och stenar.»
Sedan kom ängeln som talade med mig fram och sade till mig: »Lyft upp dina ögon och se vad det är som där kommer fram.
Och jag frågade: »Vad är det?»
Han svarade: »Det är en sädesskäppa som kommer fram.»
Ytterligare sade han: »Så är det beställt med dem i hela landet.»
Jag fick då se huru en rund skiva av bly lyfte sig; och nu syntes där en kvinna som satt i skäppan.
Därefter sade han: »Detta är Ogudaktigheten.»
Och så stötte han henne åter ned i skäppan och slog igen blylocket över dess öppning.
När jag sedan lyfte upp mina ögon, fick jag se två kvinnor komma fram; och vinden fyllde deras vingar, ty de hade vingar lika hägerns.
Och de lyfte upp skäppan mellan jord och himmel.
Då frågade jag ängeln som talade med mig: »Vart föra de skäppan?»
Han svarade mig: »De hava i sinnet att bygga ett hus åt henne i Sinears land; och när det är färdigt, skall hon där bliva nedsatt på sin plats.»
När jag sedan åter lyfte upp mina ögon, fick jag se fyra vagnar komma fram mellan två berg, och bergen voro av koppar.
För den första vagnen voro röda hästar, för den andra vagnen svarta hästar,
för den tredje vagnen vita hästar, och för den fjärde vagnen fläckiga hästar, starkare än de andra.
Då tog jag till orda och frågade ängeln som talade med mig: »Vad betyda dessa, min herre?»
Ängeln svarade och sade till mig: »Det är himmelens fyra vindar, vilka nu draga ut, sedan de hava fått träda inför hela jordens Herre.
Vagnen med de svarta hästarna drager mot nordlandet, de vita följa efter dem, och de fläckiga draga mot sydlandet.»
Men när de som voro starkast skulle draga ut, voro de ivriga att få fara omkring på jorden.
Då sade han: »Ja, I mån fara omkring på jorden.»
Och de foro åstad omkring på jorden.
Därefter ropade han på mig och talade till mig och sade: »Se, genom dem som draga ut mot nordlandet skall jag släcka min vrede på nordlandet.»
Och HERRENS ord kom till mig; han sade:
Tag emot av Heldai gåvorna från de landsflyktiga, från Tobia och Jedaja; du själv må redan samma dag gå åstad bort till Josias, Sefanjas sons, hus, dit dessa hava kommit från Babel.
När du så har fått silver och guld, skall du därav låta göra kronor; och du skall sätta en på översteprästen Josuas, Josadaks sons, huvud.
Och du skall säga till honom: »Så säger HERREN Sebaot: Se, där är en man som skall kallas Telningen.
Under honom skall det gro, och han skall bygga upp HERRENS tempel.
Ja, han skall bygga upp HERRENS tempel och förvärva majestät och sitta på sin tron och regera; och en präst skall han vara på sin tron; och fridens rådslag skola vara mellan båda.
Men kronorna skola förvaras i HERRENS tempel, till en åminnelse av Helem, Tobia och Jedaja och Hen, Sefanjas son.
Och fjärran ifrån skall man komma och bygga på HERRENS tempel; och I skolen så förnimma att HERREN Sebaot har sänt mig till eder.
Och så skall ske, om I troget hören HERRENS, eder Guds, röst.»
Och i konung Darejaves' fjärde regeringsår hände sig att HERRENS ord kom till Sakarja, på fjärde dagen i nionde månaden, det är Kisleu.
Ty från Betel hade då Sareser och Regem-Melek med sina män blivit sända för att bönfalla inför HERREN;
de skulle nämligen fråga prästerna i HERREN Sebaots hus och profeterna sålunda: »Skola vi framgent hålla gråtodag och späka oss i femte månaden, såsom vi hava gjort nu i så många år?»
Så kom då HERREN Sebaots ord till mig; han sade:
Säg till allt folket i landet och till prästerna: När I nu under sjuttio år haven hållit faste- och klagodagar i femte och i sjunde månaden, har det då varit åt mig som I haven hållit fasta?
Och när I äten och dricken, är det icke då för eder egen räkning som I äten och dricken?
Haven I icke förnummit de ord som HERREN lät predika genom forna tiders profeter, medan Jerusalem ännu tronade i god ro med sina städer omkring sig, och medan Sydlandet och Låglandet ännu voro bebodda?
Vidare kom HERRENS ord till Sakarja; han sade:
Så sade ju HERREN Sebaot: »Dömen rätta domar, och bevisen varandra kärlek och barmhärtighet.
Förtrycken icke änkan och den faderlöse, främlingen och den fattige, och tänken icke i edra hjärtan ut ont mot varandra.»
Men de ville icke akta därpå, utan spjärnade emot i gensträvighet och tillslöto sina öron för att slippa att höra.
ja, de gjorde sina hjärtan hårda såsom diamant, för att slippa att höra den lag och de ord som HERREN Sebaot genom sin Ande hade sänt, förmedelst forna tiders profeter.
Därför utgick stor vrede från HERREN Sebaot.
Och det skedde, att likasom de icke hade velat höra, när han ropade, så sade nu HERREN Sebaot: »Jag vill icke höra, när de ropa;
utan jag skall förströ dem såsom genom en stormvind bland allahanda hednafolk som de icke känna.»
Så har nu landet blivit öde efter dem, så att ingen färdas där, vare sig fram eller tillbaka; ty de hava så gjort det ljuvliga landet till en ödemark.
Vidare kom HERREN Sebaots ord; han sade:
Så säger HERREN Sebaot: Jag har stor nitälskan för Sion, ja, med stor vrede nitälskar jag för henne.
Så säger HERREN: Jag vill vända: åter till Sion och taga min boning i Jerusalem; och Jerusalem skall kallas »den trogna staden», och HERREN Sebaots berg »det heliga berget».
Så säger HERREN Sebaot: Ännu en gång skola gamla män och gamla kvinnor vara att finna på gatorna i Jerusalem, var och en med sin stav i handen, för hög ålders skull.
Och stadens gator skola vara fulla av gossar och flickor, som leka där på gatorna,
Så säger HERREN Sebaot.
Om än sådant på den tiden kan komma att synas alltför underbart för kvarlevan av detta folk, icke måste det väl därför synas alltför underbart också för mig? säger HERREN Sebaot.
Så säger HERREN Sebaot: Se, jag skall frälsa mitt folk ut ur både österland och västerland
och låta dem komma och bosätta sig i Jerusalem; och de skola vara mitt folk, och jag skall vara deras Gud, i sanning och rättfärdighet.
Så säger HERREN Sebaot: Fatten mod, I som i denna tid hören dessa ord av samma profeters mun, som talade på den tid då grunden lades till HERREN Sebaots hus, templet som skulle byggas upp.
Ty före den tiden var människornas arbete lönlöst och djurens arbete fåfängt; ingen hade någon ro för sina ovänner, vare sig han gick ut eller in, ty jag eggade alla människor mot varandra.
Men nu är jag icke mer så sinnad mot kvarlevan av detta folk som jag var i forna dagar, säger HERREN Sebaot.
Ty nu skall friden skaffa utsäde, vinträdet skall giva sin frukt, jorden skall giva sin gröda, och himmelen skall giva sin dagg; och jag skall låta kvarlevan av detta folk få allt detta till sin arvedel.
Och det skall ske, att likasom I, både Juda hus och Israels hus, haven varit ett exempel som man har nämnt, när man förbannade bland hedningarna, så skolen I nu, då jag har frälsat eder, tvärtom bliva nämnda, när man välsignar.
Frukten icke, utan fatten mod.
Ty så säger HERREN Sebaot: Likasom jag, när edra fäder förtörnade mig, beslöt att göra eder ont, säger HERREN Sebaot, och icke sedan ångrade det,
så har jag tvärtom i denna tid beslutit att göra gott mot Jerusalem och Juda hus; frukten icke.
Men detta är vad I skolen göra: Talen sanning med varandra; domen rätta och fridsamma domar i edra portar.
Tänken icke i edra hjärtan ut ont mot varandra, och älsken icke falska eder; ty allt sådant hatar jag, säger HERREN.
Och HERREN Sebaots ord kom till mig; han sade:
Så säger HERREN Sebaot: Fastedagarna i fjärde, femte, sjunde och tionde månaden skola för Juda hus bliva till fröjd och glädje och till sköna högtider.
Men älsken sanning och frid.
Så säger HERREN Sebaot: Ännu en gång skall det ske att folk skola komma hit och många städers invånare;
och invånarna i den ena staden skola gå till den andra och säga: »Upp, låtom oss gå åstad och bönfalla inför HERREN och söka HERREN Sebaot; jag själv vill ock gå åstad.»
Ja, många folk och mäktiga hednafolk skola komma och söka HERREN Sebaot i Jerusalem och bönfalla inför HERREN,
Så säger HERREN Sebaot: På den tiden skall det ske att tio män av allahanda tungomål som talas bland hednafolken skola fatta en judisk man i mantelfliken och säga: »Låt oss gå med eder, ty vi hava hört att Gud är med eder.»
Detta är en utsaga som innehåller HERRENS ord över Hadraks land; också i Damaskus skall den slå ned -- ty HERREN har sitt öga på andra människor såväl som på Israels alla stammar.
Den drabbar ock Hamat, som gränsar därintill, så ock Tyrus och Sion, där man är så vis.
Tyrus byggde sig ett fäste; hon hopade silver såsom stoft och guld såsom orenlighet på gatan.
Men se, Herren skall åter göra henne fattig, han skall bryta hennes murar ned i havet, och hon själv skall förtäras av eld.
Askelon må se det med fruktan, och Gasa med stor bävan, så ock Ekron, ty dess hopp skall komma på skam.
Gasa mister sin konung, Askelon bliver en obebodd plats
Asdod skall bebos av en vanbördig hop; så skall jag utrota filistéernas stolthet.
Men när jag har ryckt blodmaten ur deras mun och styggelserna undan deras tänder då skall också av dem bliva en kvarleva åt vår Gud, de skola bliva såsom stamfurstar i Juda, och Ekrons folk skall bliva såsom jebuséerna.
Och jag skall slå upp mitt läger till ett värn för mitt hus, mot härar som komma eller gå, och ej mer skall någon plågare komma över dem; ty jag vaktar nu med öppna ögon.
Fröjda dig storligen, du dotter Sion; höj jubelrop, du dotter Jerusalem.
Se, din konung kommer till dig; rättfärdig och segerrik är han.
Han kommer fattig, ridande på en åsna, på en åsninnas fåle.
Så skall jag utrota vagnar Efraim och hästar ur Jerusalem; ja, stridens bågar skola utrotas, och han skall tala frid till folken.
Och hans herradöme skall nå från hav till hav, och ifrån floden intill jordens ändar.
För ditt förbundsblods skull vill jag ock släppa dina fångar fria ur gropen där intet vatten finnes.
Så vänden då åter till edert fäste, I fångar som nu haven ett hopp.
Ja, det vare eder förkunnat i dag att jag vill giva eder dubbelt igen.
Ty jag skall spänna Juda såsom min båge och lägga Efraim såsom pil på den, och dina söner, du Sion, skall jag svänga såsom spjut mot dina söner, du Javan, och göra dig lik en hjältes svärd.
Ja, HERREN skall uppenbara sig i höjden, och såsom en ljungeld skall hans pil fara ut; Herren, HERREN skall stöta i basunen, och med sunnanstormar skall han draga fram.
HERREN Sebaot, han skall beskärma dem; de skola uppsluka sina fiender och trampa deras slungstenar under fötterna; under stridslarm skola de svälja sina fiender såsom vin, till dess de själva äro så fulla av blod som offerskålar och altarhörn.
Och HERREN, deras Gud, skall på den tiden giva dem seger, ty de äro ju det folk som han har till sin hjord.
Ja, ädelstenar äro de i en krona, strålande över hans land.
Huru stor bliver icke deras lycka, huru stor deras härlighet!
Av deras säd skola ynglingar blomstra upp, och jungfrur av deras vin.
HERREN mån I bedja om regn, när vårregnets tid är inne; HERREN är det som sänder ljungeldarna.
Regn skall han då giva människorna i ymnigt mått, gröda på marken åt var och en.
Men husgudarnas tal är fåfänglighet, spåmännens syner äro lögn, tomma drömmar är vad de tala, och den tröst de giva är ett intet.
Därför måste folket draga hädan såsom en fårhjord och fara illa, där det går utan herde.
Mot herdarna är min vrede upptänd och bockarna skall jag hemsöka.
Ja, HERREN Sebaot skall vårda sig om sin hjord, Juda hus, och skall så göra den till en stolt stridshäst åt sig.
Från den hjorden skall en hörnsten komma, från den en stödjepelare, från den en båge till striden, från den allt vad styresman heter.
Och de skola vara lika hjältar, som gå fram i striden, likasom trampade de i orenlighet på gatan.
Ja, strida skola de, ty HERREN är med dem, och ryttarna på sina hästar skola då komma på skam.
Jag skall giva styrka åt Juda hus, och åt Josefs hus skall jag giva seger.
Jag skall i min barmhärtighet låta dem komma tillbaka, och det skall bliva såsom hade jag aldrig förkastat dem.
Ty jag är HERREN, deras Gud, och skall bönhöra dem.
Och Efraims män skola bliva lika hjältar, och deras hjärtan skola glädja sig såsom av vin.
Deras barn skola ock se det och bliva glada; deras hjärtan skola fröjda sig i HERREN.
Jag skall locka på dem och samla dem tillhopa, ty jag förlossar dem; och de skola bliva lika talrika som de fordom voro.
Och när jag planterar ut dem bland folken, skola de tänka på mig i fjärran land; och med sina barn skola de få leva och komma tillbaka.
Ja, från Egyptens land skall jag låta dem komma tillbaka och från Assur skall jag församla dem.
Sedan skall jag föra dem till Gileads land och till Libanon; och där skall icke finnas rum nog för dem.
Han skall draga fram genom havet på en trång väg, böljorna i havet skall han slå ned, och alla Nilflodens djup skola torka ut.
Så skall Assurs stolthet bliva nedbruten och spiran tagen ifrån Egypten.
Men dem skall jag göra starka i HERREN, och i hans namn skola de gå fram, säger HERREN.
Öppna dina dörrar, Libanon, ty eld skall nu förtära dina cedrar.
Jämra dig, du cypress, ty cedern måste falla, de härliga träden skola förödas.
Jämren eder, I Basans ekar, ty skogen, den ogenomträngliga, varder fälld.
Hör huru herdarna jämra sig, när deras härlighet bliver förödd!
Hör huru de unga lejonen ryta, när Jordanbygdens snår varda förödda!
Så sade HERREN, min Gud: »Bliv en herde för slaktfåren,
ty deras köpare slakta dem utan all försyn, och deras säljare säga: 'Lovad vare HERREN att jag bliver allt rikare.'
Ej heller skonas de av sina egna herdar.»
»Se, jag vill nu icke mer skona landets inbyggare», säger HERREN, »utan låta människorna falla i varandras hand och i sina konungars hand, och dessa skola fördärva landet, och jag skall icke rädda någon ur deras hand.»
Så blev jag en herde för slaktfåren, de arma fåren.
Och jag tog mig två stavar, den ena kallade jag Ljuvlig ro, den andra kallade jag Endräkt; och jag vaktade så fåren
Men sedan jag inom en månad hade förgjort de tre herdarna, blev jag led vid fåren, likasom ock deras sinne var avogt mot mig.
Då sade jag: »Jag vill icke mer vara eder herde.
Vad som vill dö, det må dö, och vad som vill förgås, det må förgås; och de som sedan bliva kvar må äta varandras kött.»
Så tog jag min stav Ljuvlig ro och bröt sönder den, till att upplösa det förbund som jag hade slutit med alla folk.
Och när detta nu på den dagen blev upplöst, förnummo de arma fåren, som aktade på mig, att det var HERRENS ord.
Därefter sade jag till dem: »Om I så finnen för gott, så given mig min lön; varom icke, må det så vara.»
Och de vägde upp trettio siklar silver såsom lön åt mig.
Då sade HERREN till mig: »Kasta det åt krukmakaren» -- det härliga pris vartill jag hade blivit värderad av dem!
Och jag tog de trettio silversiklarna och kastade dem i HERRENS hus åt krukmakaren.
Därefter bröt jag sönder min andra stav, Endräkt, till att upplösa broderskapet mellan Juda och Israel.
Och HERREN sade till mig: »Tag dig nu redskap såsom en oförnuftig herde;
ty se, jag vill låta en herde uppstå i landet, som icke vårdar sig om de får som hålla på att förgås, icke uppsöker det förskingrade, icke helar det sargade, icke sörjer för det som är helbrägda, utan allenast äter köttet av de feta och river sönder klövarna på dem.»
Ve över denne ovärdige herde, som övergiver sin hjord!
Må ett svärd träffa hans arm och hans högra öga!
Må hans arm alldeles förtvina och hans högra öga förmörkas i grund!
Detta är en utsaga som innehåller HERRENS ord över Israel.
Så säger HERREN, han som har utspänt himmelen och grundat jorden och danat människans ande i henne:
Se, jag skall göra Jerusalem till an berusningens kalk för alla folk runt omkring; jämväl över Juda skall det komma, när Jerusalem bliver belägrat.
Och det skall ske på den tiden att jag skall göra Jerusalem till en lyftesten för alla folk; var och en som försöker lyfta den skall illa sarga sig därpå.
Och alla jordens folk skola församla sig mot det.
På den tiden, säger HERREN, skall jag slå alla hästar med förvirring och deras ryttare med vanvett.
Men över Juda hus skall jag upplåta mina ögon, när jag bland hednafolken slår alla hästar med blindhet.
Då skola Juda stamfurstar säga i sina hjärtan: »Jerusalems invånare äro vår styrka, genom HERREN Sebaot, sin Gud.»
På den tiden skall jag låta Juda stamfurstar bliva såsom brinnande fyrfat bland ved, och såsom eldbloss bland halmkärvar, så att de förbränna alla folk runt omkring, både åt höger och åt vänster; men Jerusalem skall framgent trona på sin plats, där Jerusalem nu är.
Och först skall HERREN giva seger åt Juda hyddor, för att icke Davids hus och Jerusalems invånare skola tillräkna sig större ära än Juda.
På den tiden skall HERREN beskärma Jerusalems invånare; den skröpligaste bland dem skall på den tiden vara såsom David, och Davids hus skall vara såsom ett gudaväsen, såsom HERRENS ängel framför dem.
Och jag skall på den tiden sätta mig i sinnet att förgöra alla folk som komma mot Jerusalem.
Men över Davids hus och över Jerusalems invånare skall jag utgjuta en nådens och bönens ande, så att de se upp till mig, och se vem de hava stungit.
Och de skola hålla dödsklagan efter honom, såsom man håller dödsklagan efter ende sonen, och skola bittert sörja honom, såsom man sörjer sin förstfödde.
Ja, på den tiden skall i Jerusalem hållas stor dödsklagan, sådan den var, som hölls i Hadadrimmon på Megiddons slätt.
Och släkterna i landet skola hålla dödsklagan var för sig: Davids hus släkt för sig, och dess kvinnor för sig, Natans hus' släkt för sig, och dess kvinnor för sig,
Levi hus' släkt för sig, och dess kvinnor för sig, Simeis släkt för sig, och dess kvinnor för sig;
så ock alla övriga släkter var för sig, och deras kvinnor för sig.
På den tiden skola Davids hus och Jerusalems invånare få en öppen brunn, till att avtvå sin synd och orenhet.
Och det skall ske på den tiden, säger HERREN Sebaot, att jag skall utrota avgudarnas namn ur landet, så att de icke mer skola nämnas; profeterna och orenhetens ande skall jag ock skaffa bort ur landet.
Och det skall ske, att om någon därefter uppträder såsom profet, så skola hans egna föräldrar, hans fader och moder, säga till honom: »Du kan icke få leva, du som talar lögn i HERRENS namn.»
Och hans egna föräldrar, hans fader och moder, skola stinga ihjäl honom, när han vill profetera.
Och det skall ske på den tiden att alla profeter skola blygas för sina syner, när de vilja profetera; och för att icke bliva röjda skola de icke mer kläda sig i mantel av hår.
Och var och en av dem skall säga: »Jag är ingen profet, en åkerman är jag; redan i min ungdom blev jag köpt till träl.»
Och om man då frågar honom: »Vad är det för sår du har på din kropp?» så skall han svara: »Dem har jag fått därhemma, hos mina närmaste.»
Svärd, upp mot min herde, mot den man som fick stå mig nära! säger HERREN Sebaot.
Må herden bliva slagen, så att fåren förskingras; ty jag vill nu vända min hand mot de svaga.
Och det skall ske i hela landet, säger HERREN, att två tredjedelar där skola utrotas och förgås; allenast en tredjedel skall där lämnas kvar.
Och den tredjedelen skall jag låta gå genom eld; jag skall luttra dem, såsom man luttrar silver, och pröva dem, såsom man prövar guld.
Så skola de åkalla mitt namn, och jag skall bönhöra dem.
Jag skall säga: »Detta är mitt folk.»
Och det skall svara: »HERREN är min Gud.»
Se, en dag skall komma, en HERRENS dag, då man i dig skall utskifta byte.
Ty jag skall församla alla folk till strid mot Jerusalem; och staden skall intagas, och husen skola plundras och kvinnorna skändas.
Och hälften av folket i staden skall föras bort i fångenskap.
Men återstoden därav skall icke bliva utrotad ur staden;
ty HERREN skall draga ut och strida mot de folken, såsom han stridde förr på drabbningens dag.
Och han skall den dagen stå med sina fötter på Oljeberget, gent emot Jerusalem, österut; och Oljeberget skall rämna mitt itu, mot öster och väster, till en mycket stor dal, i det att ena hälften av berget viker undan mot norr, och andra hälften därav mot söder.
Och I skolen fly ned i dalen mellan mina berg, ty dalen mellan bergen skall räcka ända till Asel; I skolen fly, såsom I flydden för jordbävningen i Ussias, Juda konungs, tid.
Då skall HERREN, min Gud, komma, ja, du själv och alla heliga med dig.
Och det skall ske på den dagen att ljuset skall bliva borta, ty himlaljusen skola förmörkas.
Och det bliver en dag som är ensam i sitt slag, och som är känd av HERREN, en dag då det varken är dag eller natt, en dag då det bliver ljust, när aftonen kommer.
Och det skall ske på den tiden att rinnande vatten skola utgå från Jerusalem, ena hälften mot Östra havet och andra hälften mot Västra havet; både sommar och vinter skall det vara så.
Och HERREN skall då vara konung över hela jorden; ja, på den tiden skall HERREN vara en, och hans namn ett.
Hela landet från Geba till Rimmon, söder om Jerusalem, skall då förvandlas till en slättmark; men själva staden skall trona på sin höjd, och sträcka sig från Benjaminsporten ända till den plats där den förra porten stod, till Hörnporten och Hananeltornet och till de kungliga vinpressarna;
och folket skall bo där i ro och icke mer givas till spillo, ty Jerusalem skall trona i trygghet.
Men denna hemsökelse skall HERREN låta drabba alla de folk som drogo ut för att strida mot Jerusalem: han skall låta deras kött ruttna, medan de ännu stå på sina fötter; deras ögon skola ruttna i sina hålor och deras tunga skall ruttna i deras mun.
Och det skall ske på den tiden att HERREN skall sända en stor förvirring bland dem; de skola bära hand på varandra, och den enes hand skall lyftas mot den andres.
Också Juda skall strida mot Jerusalem.
Och skatter skola samlas tillhopa från alla folk runt omkring: guld, silver och kläder i stor myckenhet.
En likadan hemsökelse skall ock drabba hästar, mulåsnor, kameler, åsnor och alla andra djur som finnas där i lägren.
Och det skall ske att alla överblivna ur alla de folk som kommo mot Jerusalem skola år efter år draga ditupp, för att tillbedja konungen HERREN Sebaot, och för att fira lövhyddohögtiden.
Men om någon av jordens folkstammar icke drager upp till Jerusalem, för att tillbedja konungen HERREN Sebaot, då skall över den icke komma något regn.
Om Egyptens folkstam icke drager åstad och kommer ditupp, så skall ej heller över den komma regn.
Detta bliver den hemsökelse som HERREN skall låta drabba de folk som icke draga upp för att fira lövhyddohögtiden.
Ja, så skall Egypten drabbas av sin synd, så skola ock alla andra folk drabbas av sin synd, om de icke draga upp för att fira lövhyddohögtiden.
På den tiden skall på hästarnas bjällror stå att läsa: »Helgad åt HERREN», och grytorna i HERRENS hus skola vara såsom offerskålarna framför altaret.
Och var gryta i Jerusalem och Juda skall vara helgad åt HERREN Sebaot, så att var och en som vill offra kan komma och taga en sådan och koka i den.
Och ingen kanané skall mer finnas i HERREN Sebaots hus, på den tiden.
Detta är en utsaga, som innehåller HERRENS ord till Israel genom Malaki.
Jag har bevisat eder kärlek, säger HERREN.
Nu frågen I: »Varmed har du då bevisat oss kärlek?»
Esau var ju en broder till Jakob, säger HERREN, och jag älskade Jakob,
men Esau hatade jag; därför gjorde jag hans berg till en ödemark och hans arvedel till ett hemvist för öknens schakaler.
Om nu Edom säger: »Ja, vi äro förstörda, men vi skola åter bygga upp det ödelagda», så svarar HERREN Sebaot: Väl må de bygga upp, men jag skall åter riva det ned, och så skall man få kalla det 'ogudaktighetens land' och 'det folk, på vilket HERREN evinnerligen vredgas'.
I skolen få se det med egna ögon, och då skolen I säga: 'HERREN är stor utöver Israels gränser.'
En son skall hedra sin fader och en tjänare sin herre.
Om nu jag är fader, var är då den heder, som skulle visas mig?
Och om jag är en herre, var är då den fruktan, som man skulle hava för mig? -- så säger HERREN Sebaot till eder, I präster, som förakten mitt namn.
Nu frågen I: »Varmed hava vi då visat förakt för ditt namn?»
Jo, därmed att I bären fram ovärdig spis på mitt altare.
Åter frågen I: »På vad sätt hava vi betett oss ovärdigt mot dig?»
Jo, i det att I tänken: »HERRENS bord behöver man icke mycket akta.»
När i fören fram ett offerdjur, som är blint, då räknen I sådant icke för ont; när I fören fram ett som är lytt eller svagt, då räknen I ej heller sådant för ont.
Kom med något sådant till din ståthållare, så får du se, om han tager gunstigt emot dig och bliver dig bevågen, säger HERREN Sebaot.
Bönfallen alltså nu inför Gud, att han må bliva oss nådig.
Kan han väl vara eder bevågen, då I haven begått sådant? säger HERREN Sebaot.
Ack att bland eder funnes någon som ville stänga tempeldörrarna, så att I icke längre förgäves upptänden eder eld på mitt altare!
Jag har icke behag till eder, säger HERREN Sebaot, och till offergåvor av eder hand har jag icke lust.
Från solens uppgång ända till dess nedgång är ju mitt namn stort bland folken, och överallt frambäras rökoffer och rena offergåvor åt mitt namn; ja, mitt namn är stort bland folken, säger HERREN Sebaot.
Men I ohelgen det, i det att I sägen: »Herrens bord kan man gärna försumma, och den spis, som gives därtill, behöver man icke mycket akta.»
Ja, I sägen: »Icke är det mödan värt!», och så handhaven I det vanvördigt, säger HERREN Sebaot.
När I alltså frambären eder offergåva, då fören I fram, vad som är rövat och vad som är lytt och svagt.
Skulle jag hava behag till sådana gåvor av eder hand? säger HERREN.
Nej, förbannad vare den bedragare, som i sin hjord har ett djur av hankön, men ändå, när han har gjort ett löfte, offrar åt Herren ett djur, som icke duger.
Ty jag är en stor konung, säger HERREN Sebaot, och mitt namn är fruktansvärt bland folken.
Därför kommer nu följande bud till eder, I präster.
Om I icke hörsammen det och akten därpå, så att I given mitt namn ära, säger HERREN Sebaot, så skall jag sända förbannelse över eder och förbanna edra välsignelser; ja, jag har redan förbannat dem, eftersom I icke akten därpå.
Se, jag skall låta min näpst drabba eder avkomma, och jag skall kasta orenlighet i ansiktet på eder, orenligheten efter edra högtidsoffer; ja, I skolen själva bliva kastade i denna.
Då skolen I förstå, att jag har sänt till eder detta bud, för att mitt förbund med Levi skall bestå, säger HERREN Sebaot.
Jag hade ett förbund med honom, och däri var liv och frid.
Sådant gav jag åt honom, för att han skulle frukta mig; och han fruktade mig och bävade för mitt namn.
Rätt undervisning var i hans mun, och ingen orätt fanns på hans läppar; fridsamt och redligt vandrade han i min umgängelse och omvände många från missgärning.
Ty prästens läppar skola förvara kunskap, och undervisning skall man hämta ur hans mun; han är ju HERREN Sebaots sändebud.
Men I haven vikit av ifrån vägen; genom eder undervisning haven I kommit många på fall.
I haven fördärvat förbundet med Levi, säger HERREN Sebaot.
Därför har ock jag gjort eder föraktade och låga i allt folkets ögon, eftersom I icke hållen mina vägar, utan haven anseende till personen, när I handhaven undervisningen.
Hava vi icke alla en och samma fader?
Har icke en och samma Gud skapat oss?
Varför handla vi då trolöst mot varandra och bryta våra fäders förbund?
Juda har handlat trolöst, och styggelse är bedriven i Israel och i Jerusalem; ty Juda har oskärat HERRENS helgedom, den som han älskar, och de hava tagit till äkta kvinnor, som dyrka främmande gudar.
Hos den man som så gör må HERREN utrota var levande själ ur Jakobs hyddor, jämväl den som frambär offergåvor till HERREN Sebaot.
Och ännu något annat gören I: I vållen, att HERRENS altare höljes med tårar, med gråt och klagan, så att han icke mer vill se till offergåvorna, ej heller med välbehag kan taga emot något ur eder hand.
Nu frågen I: »Huru så?»
Jo, HERREN var ju vittne mellan dig och din ungdoms hustru, henne som du nu har varit trolös emot, fastän hon är din maka, din äkta hustru.
Hava vi då icke en och samma skapare, den, i vilkens hand det står, att vår ande bevaras?
Och vad vill nu denne ene?
Han vill ju hava ett gudaktigt släkte.
Tagen eder därför väl till vara, så att ingen bliver trolös mot sin ungdoms hustru.
Ty jag hatar äktenskapsskillnad, säger HERREN, Israels Gud, och att man höljer sig i våld såsom i en överklädnad, säger HERREN Sebaot.
Tagen eder därför väl till vara, så att I icke bliven trolösa.
I trötten ut HERREN med edert tal.
Nu frågen I: »Varmed trötta vi då ut honom?»
Jo, därmed att I sägen: »Den som gör ont är ändå god i HERRENS ögon, och till sådana har han behag.
Ty varför kommer icke eljest domens Gud?»
Se, jag skall sända ut min ängel, och han skall bereda väg för mig.
Och med hast skall han komma till sitt tempel, den Herre, som I åstunden, ja, förbundets ängel, som I begären, se, han kommer, säger HERREN Sebaot.
Men vem kan uthärda hans tillkommelses dag, och vem kan bestå, när han uppenbarar sig?
Ty han skall vara såsom en guldsmeds eld och såsom valkares såpa.
Och han skall sätta sig ned och smälta silvret och rena det; han skall rena Levi söner och luttra dem såsom guld och silver; och sedan skola de frambära åt HERREN offergåvor i rättfärdighet.
Och Juda offergåvor och Jerusalems skola då behaga HERREN väl likasom i forna dagar och i förgångna år.
Ja, jag skall komma till eder för att hålla dom, och jag skall vara ett snarfärdigt vittne mot trollkarlar, äktenskapsbrytare och menedare, så ock mot dem som förhålla dagakarlen hans lön eller förtrycka änkan och den faderlöse eller vränga rätten för främlingen, men icke frukta mig, säger HERREN Sebaot.
Ty jag, HERREN, har icke förändrats, och I, Jakobs barn, haven icke heller hört upp:
allt ifrån edra fäders dagar haven I vikit av ifrån mina stadgar och icke hållit dem Vänden om till mig, så vill jag vända om till eder, säger HERREN Sebaot.
Nu frågen I: »Varutinnan skola vi vända om?»
Menen I då, att en människa får röva från Gud?
Ty I röven ju från mig.
Åter frågen I: »På vad sätt hava vi rövat från dig?»
Jo, i fråga om tionden och offergärden.
Förbannelse har drabbat eder, men ändå röven I från mig, så många I ären.
Fören full tionde till förrådshuset, så att i mitt hus finnes mat, och pröven så, hurudan jag sedan bliver, säger HERREN Sebaot.
Förvisso skall jag då öppna himmelens fönster över eder och utgjuta över eder riklig välsignelse.
Och jag skall näpsa gräshopporna för eder, så att de icke mer fördärva eder frukt på marken; ej heller skola edra vinträd mer slå fel på fältet, säger HERREN Sebaot.
Och alla folk skola prisa eder sälla, ty edert land skall då vara ljuvligt, säger HERREN Sebaot.
I haven talat hårda ord mot mig, säger HERREN.
Nu frågen I: »Vad hava vi då med varandra talat mot dig?»
I haven sagt: »Det är fåfängt att tjäna Gud.
Eller vad vinning hava vi därav att vi hålla, vad han har bjudit oss hålla, och därav att vi gå i sorgdräkt inför HERREN Sebaot?
Nej, de fräcka vilja vi nu prisa sälla; ty de som göra, vad ogudaktigt är, bliva upprättade, de gå fria, huru de än fresta Gud.»
Men därunder hava också de som frukta HERREN talat med varandra; och HERREN har aktat på dem och hört dem, och en minnesbok har blivit skriven inför hans ansikte till åminnelse av dessa som frukta HERREN och tänka på hans namn.
Och dessa, säger HERREN Sebaot, skall jag hava såsom min egendom på den dag, då jag utför mitt verk; och jag skall skona dem, såsom en fader skonar sin son, som tjänar honom.
Och I skolen då åter få se, vilken skillnad det är mellan den rättfärdige och den ogudaktige, mellan den som tjänar Gud och den som icke tjänar honom.
Ty se, dagen kommer, och den skall brinna såsom en ugn.
Då skola alla fräcka människor och alla som göra, vad ogudaktigt är, bliva lika strå, och dagen, den som kommer, skall förbränna dem, säger HERREN Sebaot, så att varken rot eller krona lämnas kvar av dem.
Men för eder, I som frukten mitt namn, skall rättfärdighetens sol gå upp med läkedom under sina vingar.
Då skolen I slippa ut och hoppa såsom kalvar, som hava varit instängda i stallet.
Och de ogudaktiga skolen I trampa ned, ty de skola bliva såsom aska under edra fötter på den dag, då jag utför mitt verk, säger HERREN Sebaot.
Tänken på Moses lag, min tjänares, åt vilken jag på Horeb gav stadgar och rätter för hela Israel.
Se, jag skall sända till eder profeten Elia, förrän HERRENS stora och fruktansvärda dag kommer.
Och han skall vända fädernas hjärtan till barnen och barnens hjärtan till deras fäder, för att jag icke, när jag kommer, skall slå landet med tillspillogivning.
Detta är Jesu Kristi, Davids sons, Abrahams sons, släkttavla.
Abraham födde Isak, Isak födde Jakob, Jakob födde Judas och hans bröder;
Judas födde Fares och Sara med Tamar, Fares födde Esrom, Esrom födde Aram;
Aram födde Aminadab, Aminadab födde Naasson, Naasson födde Salmon;
Salmon födde Boes med Rakab, Boes födde Jobed med Rut, Jobed födde Jessai;
Jessai födde David, konungen, David födde Salomo med Urias' hustru;
Salomo födde Roboam, Roboam födde Abia.
Abia födde Asaf;
Asaf födde Josafat, Josafat födde Joram, Joram födde Osias;
Osias födde Joatam, Joatam födde Akas, Akas födde Esekias;
Esekias födde Manasses, Manasses födde Amos, Amos födde Josias;
Josias födde Jekonias och hans bröder, vid den tid då folket blev bortfört i fångenskap till Babylonien.
Sedan folket hade blivit bortfört i fångenskap till Babylonien, födde Jekonias Salatiel, Salatiel födde Sorobabel;
Sorobabel födde Abiud, Abiud födde Eljakim, Eljakim födde Asor;
Asor födde Sadok, Sadok födde Akim, Akim födde Eliud;
Eliud födde Eleasar, Eleasar födde Mattan, Mattan födde Jakob;
Jakob födde Josef, Marias man, och av henne föddes Jesus, som kallas Kristus.
Så utgöra släktlederna från Abraham intill David tillsammans fjorton leder, och från David intill dess att folket blev bortfört i fångenskap till Babylonien fjorton leder, och från det att folket blev bortfört i fångenskap till Babylonien intill Kristus fjorton leder.
Med Jesu Kristi födelse gick det så till.
Sedan Maria, hans moder, hade blivit trolovad med Josef, befanns hon, förrän de kommo tillsammans, vara havande av helig ande.
Nu var Josef, hennes man, en rättsinnig man och ville icke utsätta henne for vanära; därför beslöt han att hemligen skilja sig från henne.
Men när han hade fått detta i sinnet, se, då visade sig i drömmen en Herrens ängel för honom och sade: »Josef, Davids son, frukta icke att taga till dig Maria, din hustru; ty det som är avlat i henne är av helig ande.
Och hon skall föda en son, och honom skall du giva namnet Jesus, ty han skall frälsa sitt folk ifrån deras synder.»
Allt detta har skett, för att det skulle fullbordas, som var sagt av Herren genom profeten som sade:
»Se, jungfrun skall bliva havande och föda en son, och man skall giva honom namnet Emmanuel» (det betyder Gud med oss).
När Josef hade vaknat upp ur sömnen, gjorde han som Herrens ängel hade befallt honom och tog sin hustru till sig.
Och han kände henne icke, förrän hon hade fött en son; och honom gav han namnet Jesus.
När nu Jesus var född i Betlehem i Judeen, på konung Herodes' tid, då kommo vise män från österns länder till Jerusalem
och sade: »Var är den nyfödde judakonungen?
Vi hava nämligen sett hans stjärna i östern och hava kommit för att giva honom vår hyllning.»
När konung Herodes hörde detta, blev han förskräckt, och hela Jerusalem med honom.
Och han församlade alla överstepräster och skriftlärde bland folket och frågade dem var Messias skulle födas.
De svarade honom: »I Betlehem i Judeen; ty så är skrivet genom profeten:
'Och du Betlehem, du judiska bygd, ingalunda är du minst bland Juda furstar, ty av dig skall utgå en furste som skall vara en herde för mitt folk Israel.'»
Då kallade Herodes hemligen till sig de vise männen och utfrågade dem noga om tiden då stjärnan hade visat sig.
Sedan lät han dem fara till Betlehem och sade: »Faren åstad och forsken noga efter barnet; och när I haven funnit det, så låten mig veta detta, för att också jag må komma och giva det min hyllning.»
När de hade hört konungens ord, foro de åstad; och se, stjärnan som de hade sett i östern gick framför dem, till dess att den kom över det ställe där barnet var.
Där stannade den.
Och när de sågo stjärnan, uppfylldes de av mycket stor glädje.
Och de gingo in i huset och fingo se barnet med Maria, dess moder.
Då föllo de ned och gåvo det sin hyllning; och de togo fram sina skatter och framburo åt det skänker: guld, rökelse och myrra.
Sedan fingo de, genom en uppenbarelse i drömmen, befallning att icke återvända till Herodes; och de drogo så en annan väg tillbaka till sitt land.
Men när de hade dragit åstad, se, då visade sig i drömmen en Herrens ängel för Josef och sade: »Stå upp och tag barnet och dess moder med dig, och fly till Egypten, och bliv kvar där, till dess jag säger dig till; ty Herodes tänker söka efter barnet för att förgöra det.»
Då stod han upp och tog barnet och dess moder med sig om natten, och drog bort till Egypten.
Där blev han kvar intill Herodes' död, för att det skulle fullbordas, som var sagt av Herren genom profeten som sade: »Ut ur Egypten kallade jag min son.»
När Herodes nu såg att han hade blivit gäckad av de vise männen, blev han mycket vred.
Och han sände åstad och lät döda alla de gossebarn i Betlehem och hela området däromkring, som voro två år gamla och därunder, detta enligt den uppgift om tiden, som han hade fått genom att utfråga de vise männen.
Då fullbordades det som var sagt genom profeten Jeremias, när han sade:
»Ett rop hördes i Rama, gråt och mycken jämmer; det var Rakel som begrät sina barn, och hon ville icke låta trösta sig, eftersom de icke mer voro till.»
Men när Herodes var död, se, då visade sig i drömmen en Herrens ängel for Josef, i Egypten,
och sade: »Stå upp och tag barnet och dess moder med dig, och begiv dig till Israels land; ty de som traktade efter barnets liv äro nu döda.»
Då stod han upp och tog barnet och dess moder med sig, och kom så till Israels land.
Men när han hörde att Arkelaus regerade över Judeen; efter sin fader Herodes, fruktade han att begiva sig dit; och på grund av en uppenbarelse i drömmen drog han bort till Galileens bygder.
Och när han hade kommit dit, bosatte han sig i en stad som hette Nasaret, för att det skulle fullbordas, som var sagt genom profeterna, att han skulle kallas nasaré.
Vid den tiden uppträdde Johannes döparen och predikade i Judeens öken
och sade: »Gören bättring, ty himmelriket är nära.»
Det var om denne som profeten Esaias talade, när han sade: »Hör rösten av en som ropar i öknen: 'Bereden vägen för Herren, gören stigarna jämna för honom.'»
Och Johannes hade kläder av kamelhår och bar en lädergördel om sina länder, och hans mat var gräshoppor och vildhonung.
Och från Jerusalem och hela Judeen och hela trakten omkring Jordan gick då folket ut till honom
och lät döpa sig av honom i floden Jordan, och bekände därvid sina synder.
Men när han såg många fariséer och sadducéer komma för att låta döpa sig, sade han till dem: »I huggormars avföda, vem har ingivit eder att söka komma undan den tillstundande vredesdomen?
Bären då ock sådan frukt som tillhör bättringen.
Och menen icke att I kunnen säga vid eder själva: 'Vi hava ju Abraham till fader'; ty jag säger eder att Gud av dessa stenar kan uppväcka barn åt Abraham.
Och redan är yxan satt till roten på träden; så bliver då vart träd som icke bär god frukt avhugget och kastat i elden.
Jag döper eder i vatten till bättring, men den som kommer efter mig, han är starkare än jag, och jag är icke ens värdig att bära hans skor; han skall döpa eder i helig ande och eld.
Han har sin kastskovel i handen, och han skall noga rensa sin loge och samla in sitt vete i ladan; men agnarna skall han bränna upp i en eld som icke utsläckes.»
Därefter kom Jesus från Galileen till Johannes, vid Jordan, för att låta döpa sig av honom;
men denne ville hindra honom och sade: »Jag behövde döpas av dig, och du kommer till mig?»
Då svarade Jesus och sade till honom: »Låt det nu så ske; ty det höves oss att så uppfylla all rättfärdighet.
Då tillstadde han honom det.
Och när Jesus var döpt, steg han strax upp ur vattnet; och se, då öppnades himmelen, och han såg Guds Ande sänka sig ned såsom en duva och komma över honom.
Och från himmelen kom en röst, som sade: »Denne är min älskade Son, i vilken jag har funnit behag.»
Därefter blev Jesus av Anden förd upp i öknen, för att han skulle frestas av djävulen.
Och när han hade fastat i fyrtio dagar och fyrtio nätter, blev han omsider hungrig.
Då trädde frestaren fram och sade till honom: »Är du Guds Son, så bjud att dessa stenar bliva bröd.»
Men han svarade och sade: »Det är skrivet: 'Människan skall leva icke allenast av bröd, utan av allt det som utgår av Guds mun.'»
Därefter tog djävulen honom med sig till den heliga staden och ställde honom uppe på helgedomens mur
och sade till honom: »Är du Guds Son, så kasta dig ned; det är ju skrivet: 'Han skall giva sina änglar befallning om dig, och de skola bära dig på händerna, så att du icke stöter din fot mot någon sten.'»
Jesus sade till honom: »Det är ock skrivet: 'Du skall icke fresta Herren, din Gud.'»
Åter tog djävulen honom med sig, upp på ett mycket högt berg, och visade honom alla riken i världen och deras härlighet
och sade till honom: »Allt detta vill jag giva dig, om du faller ned och tillbeder mig.»
Då sade Jesus till honom: »Gå bort, Satan; ty det är skrivet: 'Herren, din Gud, skall du tillbedja, och honom allena skall du tjäna.'»
Då lämnade djävulen honom; och se, änglar trädde fram och betjänade honom.
Men när han hörde att Johannes hade blivit satt i fängelse, drog han sig tillbaka till Galileen.
Och han lämnade Nasaret och begav sig till Kapernaum, som ligger vid sjön, på Sabulons och Neftalims område, och bosatte sig där,
för att det skulle fullbordas, som var sagt genom profeten Esaias, när han sade:
»Sabulons land och Neftalims land, trakten åt havet till, landet på andra sidan Jordan, hedningarnas Galileen --
det folk som där satt i mörker fick se ett stort ljus; ja, de som sutto i dödens ängd och skugga, för dem gick upp ett ljus.»
Från den tiden begynte Jesus predika och säga: »Gören bättring, ty himmelriket är nära.»
Då han nu vandrade utmed Galileiska sjön, fick han se två bröder, Simon, som kallas Petrus, och Andreas, hans broder, kasta ut nät i sjön, ty de voro fiskare.
Och han sade till dem: »Följen mig så skall jag göra eder till människofiskare.»
Strax lämnade de näten och följde honom.
När han hade gått därifrån ett stycke längre fram, fick han se två andra bröder, Jakob, Sebedeus' son, och Johannes, hans broder, där de jämte sin fader Sebedeus sutto i båten och ordnade sina nät; och han kallade dem till sig.
Och strax lämnade de båten och sin fader och följde honom.
Och han gick omkring i hela Galileen och undervisade i deras synagogor och predikade evangelium om riket och botade alla slags sjukdomar och allt slags skröplighet bland folket.
Och ryktet om honom gick ut över hela Syrien, och man förde till honom alla sjuka som voro hemsökta av olika slags lidanden och plågor, alla som voro besatta eller månadsrasande eller lama; och han botade dem.
Och honom följde mycket folk ifrån Galileen och Dekapolis och Jerusalem och Judeen och från landet på andra sidan Jordan.
När han nu såg folket, gick han upp på berget; och sedan han hade satt sig ned, trädde hans lärjungar fram till honom.
Då öppnade han sin mun och undervisade dem och sade:
»Saliga äro de som äro fattiga i anden, ty dem hör himmelriket till.
Saliga äro de som sörja, ty de skola bliva tröstade.
Saliga äro de saktmodiga, ty de skola besitta jorden.
Saliga äro de som hungra och törsta efter rättfärdighet, ty de skola bliva mättade.
Saliga äro de barmhärtiga, ty dem skall vederfaras barmhärtighet.
Saliga äro de renhjärtade, ty de skola se Gud.
Saliga äro de fridsamma, ty de skola kallas Guds barn.
Saliga äro de som lida förföljelse för rättfärdighets skull, ty dem hör himmelriket till.
Ja, saliga ären I, när människorna för min skull smäda och förfölja eder och sanningslöst säga allt ont mot eder.
Glädjens och fröjden eder, ty eder lön är stor i himmelen.
Så förföljde man ju ock profeterna, som voro före eder.
I ären jordens salt; men om saltet mister sin sälta, varmed skall man då giva det sälta igen?
Till intet annat duger det än till att kastas ut och trampas ned av människorna.
I ären världens ljus.
Icke kan en stad döljas, som ligger uppe på ett berg?
Ej heller tänder man ett ljus och sätter det under skäppan, utan man sätter det på ljusstaken, så att det lyser för alla dem som äro i huset.
På samma sätt må ock edert ljus lysa inför människorna, så att de se edra goda gärningar och prisa eder Fader, som är i himmelen.
I skolen icke mena att jag har kommit för att upphäva lagen eller profeterna.
Jag har icke kommit för att upphäva, utan för att fullborda.
Ty sannerligen säger jag eder: Intill dess himmel och jord förgås, skall icke den minsta bokstav, icke en enda prick av lagen förgås, förrän det allt har fullbordats.
Därför, den som upphäver ett av de minsta bland dessa bud och lär människorna så, han skall räknas för en av de minsta i himmelriket; men den som håller dem och lär människorna så, han skall räknas för stor i himmelriket.
Ty jag säger eder, att om eder rättfärdighet icke övergår de skriftlärdes och fariséernas, så skolen I icke komma in i himmelriket.
I haven hört att det är sagt till de gamle: 'Du skall icke dräpa; och den som dräper, han är hemfallen åt Domstolens dom.'
Men jag säger eder: Var och en som vredgas på sin broder, han är hemfallen åt Domstolens dom; men den som säger till sin broder: 'Du odåga', han är hemfallen åt Stora rådets dom; och den som säger: 'Du dåre', han är hemfallen åt det brinnande Gehenna.
Därför, om du kommer med din gåva till altaret, och där drager dig till minnes att din broder har något emot dig,
så lägg ned din gåva där framför altaret, och gå först bort och förlik dig med din broder, och kom sedan och bär fram din gåva.
Var villig till snar förlikning med din motpart, medan du ännu är med honom på vägen, så att din motpart icke drager dig inför domaren, och domaren överlämnar dig åt rättstjänaren, och du bliver kastad i fängelse.
Sannerligen säger jag dig: Du skall icke slippa ut därifrån, förrän du har betalt den yttersta skärven.
I haven hört att det är sagt: 'Du skall icke begå äktenskapsbrott.'
Men jag säger eder: Var och en som med begärelse ser på en annans hustru, han har redan begått äktenskapsbrott med henne i sitt hjärta.
Om nu ditt högra öga är dig till förförelse, så riv ut det och kasta det ifrån dig; ty det är bättre för dig att en av dina lemmar fördärvas, än att hela din kropp kastas i Gehenna.
Och om din högra hand är dig till förförelse, så hugg av den och kasta den ifrån dig; ty det är bättre för dig att en av dina lemmar fördärvas, än att hela din kropp kommer till Gehenna.
Det är ock sagt: 'Den som vill skilja sig från sin hustru han skall giva henne skiljebrev.'
Men jag säger eder: Var och en som skiljer sig från sin hustru för någon annan saks skull än för otukt, han bliver orsak till att äktenskapsbrott begås med henne.
Och den som tager en frånskild kvinna till hustru, han begår äktenskapsbrott.
Ytterligare haven I hört att det är sagt till de gamle: 'Du skall icke svärja falskt' och 'Du skall hålla din ed inför Herren.'
Men jag säger eder att I alls icke skolen svärja, varken vid himmelen, ty den är 'Guds tron',
ej heller vid jorden, ty den är 'hans fotapall', ej heller vid Jerusalem, ty det är 'den store Konungens stad';
ej heller må du svärja vid ditt huvud, ty du kan icke göra ett enda hår vare sig vitt eller svart;
utan sådant skall edert tal vara, att ja är ja, och nej är nej.
Vad därutöver är, det är av ondo.
I haven hört att det är sagt: 'Öga för öga och tand för tand.'
Men jag säger eder att I icke skolen stå emot en oförrätt; utan om någon slår dig på den högra kinden, så vänd ock den andra till åt honom;
och om någon vill gå till rätta med dig för att beröva dig din livklädnad, så låt honom få manteln med;
och om någon tvingar dig att till hans tjänst gå med en mil, så gå två med honom.
Giv åt den som beder dig, och vänd dig icke bort ifrån den som vill låna av dig.
I haven hört att det är sagt: 'Du skall älska din nästa och hata din ovän.'
Men jag säger eder: Älsken edra ovänner, och bedjen för dem som förfölja eder,
och varen så eder himmelske Faders barn; han låter ju sin sol gå upp över både onda och goda och låter det regna över både rättfärdiga och orättfärdiga.
Ty om I älsken dem som älska eder, vad lön kunnen I få därför?
Göra icke publikanerna detsamma?
Och om I visen vänlighet mot edra bröder allenast, vad synnerligt gören I därmed?
Göra icke hedningarna detsamma?
Varen alltså I fullkomliga, såsom eder himmelske Fader är fullkomlig.»
»Tagen eder till vara för att öva eder rättfärdighet inför människorna, för att bliva sedda av dem; annars haven I ingen lön hos eder Fader, som är i himmelen.
Därför, när du giver en allmosa, så låt icke stöta i basun för dig, såsom skrymtarna göra i synagogorna och på gatorna, för att de skola bliva prisade av människorna.
Sannerligen säger jag eder: De hava fått ut sin lön.
Nej, när du giver en allmosa, låt då din vänstra hand icke få veta vad den högra gör,
så att din allmosa gives i det fördolda.
Då skall din Fader, som ser i det fördolda, vedergälla dig.
Och när I bedjen, skolen I icke vara såsom skrymtarna, vilka gärna stå i synagogorna och i gathörnen och bedja, för att bliva sedda av människorna.
Sannerligen säger jag eder: De hava fått ut sin lön.
Nej, när du vill bedja, gå då in i din kammare, och stäng igen din dörr, och bed till din Fader i det fördolda.
Då skall din Fader, som ser i det fördolda, vedergälla dig.
Men i edra böner skolen I icke hopa tomma ord såsom hedningarna, vilka mena att de skola bliva bönhörda för sina många ords skull.
Så varen då icke lika dem; eder Fader vet ju vad I behöven, förrän I bedjen honom.
I skolen alltså bedja sålunda: 'Fader vår, som är i himmelen!
Helgat varde ditt namn;
tillkomme ditt rike; ske din vilja, såsom i himmelen, så ock på jorden;
vårt dagliga bröd giv oss i dag;
och förlåt oss våra skulder, såsom ock vi förlåta dem oss skyldiga äro;
och inled oss icke i frestelse, utan fräls oss ifrån ondo.'
Ty om I förlåten människorna deras försyndelser, så skall ock eder himmelske Fader förlåta eder;
men om I icke förlåten människorna, så skall ej heller eder Fader förlåta edra försyndelser.
Och när I fasten, skolen I icke visa en bedrövad uppsyn såsom skrymtarna, vilka vanställa sina ansikten för att bliva sedda av människorna med sin fasta.
Sannerligen säger jag eder: De hava fått ut sin lön.
Nej, när du fastar, smörj då ditt huvud och två ditt ansikte,
för att du icke må bliva sedd av människorna med din fasta, utan allenast av din Fader, som är i det fördolda.
Då skall din Fader, som ser i det fördolda, vedergälla dig.
Samlen eder icke skatter på jorden, där mott och mal förstöra, och där tjuvar bryta sig in och stjäla,
utan samlen eder skatter i himmelen, där mott och mal icke förstöra, och där inga tjuvar bryta sig in och stjäla.
Ty där din skatt är, där kommer ock ditt hjärta att vara.
Ögat är kroppens lykta.
Om nu ditt öga är friskt, så får hela din kropp ljus.
Men om ditt öga är fördärvat, då bliver hela din kropp höljd i mörker.
Är det nu så, att ljuset, som du har i dig, är mörker, huru djupt bliver då icke mörkret!
Ingen kan tjäna två herrar; ty antingen kommer han då att hata den ene och älska den andre, eller kommer han att hålla sig till den förre och förakta den senare.
I kunnen icke tjäna både Gud och Mamon.
Därför säger jag eder: Gören eder icke bekymmer för edert liv, vad I skolen äta eller dricka, ej heller för eder kropp, vad I skolen kläda eder med.
Är icke livet mer än maten, och kroppen mer än kläderna?
Sen på fåglarna under himmelen: de så icke, ej heller skörda de, ej heller samla de in i lador; och likväl föder eder himmelske Fader dem.
Ären I icke mycket mer än de?
Vilken av eder kan, med allt sitt bekymmer, lägga en enda aln till sin livslängd?
Och varför bekymren I eder för kläder?
Beskåden liljorna på marken, huru de växa: de arbeta icke, ej heller spinna de;
och likväl säger jag eder att icke ens Salomo i all sin härlighet var så klädd som en av dem.
Kläder nu Gud så gräset på marken, vilket i dag står och i morgon kastas i ugnen, skulle han då icke mycket mer kläda eder, I klentrogne?
Så gören eder nu icke bekymmer, och sägen icke: 'Vad skola vi äta?' eller: 'Vad skola vi dricka?' eller: 'Vad skola vi kläda oss med?'
Efter allt detta söka ju hedningarna, och eder himmelske Fader vet att I behöven allt detta.
Nej, söken först efter hans rike och hans rättfärdighet, så skall också allt detta andra tillfalla eder.
Gören eder alltså icke bekymmer för morgondagen, ty morgondagen skall själv bära sitt bekymmer.
Var dag har nog av sin egen plåga.»
»Dömen icke, på det att I icke mån bliva dömda;
ty med den dom varmed I dömen skolen I bliva dömda, och med det mått som I mäten med skall ock mätas åt eder.
Huru kommer det till, att du ser grandet i din broders öga, men icke bliver varse bjälken i ditt eget öga?
Eller huru kan du säga till din broder: 'Låt mig taga ut grandet ur ditt öga', du som har en bjälke i ditt eget öga?
Du skrymtare, tag först ut bjälken ur ditt eget öga; därefter må du se till, att du kan taga ut grandet ur din broders öga.
Given icke åt hundarna vad heligt är, och kasten icke edra pärlor för svinen, på det att dessa icke må trampa dem under fötterna och sedan vända sig om och sarga eder.
Bedjen, och eder skall varda givet; söken, och I skolen finna; klappen, och för eder skall varda upplåtet.
Ty var och en som beder, han får; och den som söker, han finner; och för den som klappar skall varda upplåtet.
Eller vilken är den man bland eder, som räcker sin son en sten, när han beder honom om bröd,
eller som räcker honom en orm, när han beder om fisk?
Om nu I, som ären onda, förstån att giva edra barn goda gåvor, huru mycket mer skall icke då eder Fader, som är i himmelen, giva vad gott är åt dem som bedja honom!
Därför, allt vad I viljen att människorna skola göra eder, det skolen I ock göra dem; ty detta är lagen och profeterna.
Gån in genom den trånga porten.
Ty vid och bred är den väg som leder till fördärvet, och många äro de som gå fram på den;
och den port är trång och den väg är smal, som leder till livet, och få äro de som finna den.
Tagen eder till vara för falska profeter, som komma till eder i fårakläder, men invärtes äro glupande ulvar.
Av deras frukt skolen I känna dem.
Icke hämtar man väl vindruvor från törnen, eller fikon från tistlar?
Så bär vart och ett gott träd god frukt, men ett dåligt träd bär ond frukt.
Ett gott träd kan icke bära ond frukt, ej heller kan ett dåligt träd bära god frukt.
Vart träd som icke bär god frukt bliver avhugget och kastat i elden.
Alltså skolen I känna dem av deras frukt. --
Icke kommer var och en in i himmelriket, som säger till mig: 'Herre, Herre', utan den som gör min himmelske Faders vilja.
Många skola på 'den dagen' säga till mig: 'Herre, Herre, hava vi icke profeterat i ditt namn och genom ditt namn drivit ut onda andar och genom ditt namn gjort många kraftgärningar?'
Men då skall jag betyga för dem: 'Jag har aldrig känt eder; gån bort ifrån mig, I ogärningsmän.'
Därför, var och en som hör dessa mina ord och gör efter dem, han må liknas vid en förståndig man som byggde sitt hus på hälleberget.
Och slagregn föll, och vattenströmmarna kommo, och vindarna blåste och kastade sig mot det huset; och likväl föll det icke omkull, eftersom det var grundat på hälleberget.
Men var och en som hör dessa mina ord och icke gör efter dem, han må liknas vid en oförståndig man som byggde sitt hus på sanden.
Och slagregn föll, och vattenströmmarna kommo, och vindarna blåste och slogo mot det huset; och det föll omkull, och dess fall var stort.»
När Jesus hade slutat detta tal, häpnade folket över hans förkunnelse;
ty han förkunnade sin lära för dem med makt och myndighet, och icke såsom deras skriftlärde.
Sedan han hade kommit ned från berget, följde honom mycket folk.
Då trädde en spetälsk man fram och föll ned för honom och sade: »Herre, vill du, så kan du göra mig ren.»
Då räckte han ut handen och rörde vid honom och sade: »Jag vill; bliv ren.»
Och strax blev han ren från sin spetälska.
Och Jesus sade till honom: »Se till, att du icke säger detta för någon; men gå bort och visa dig för prästen, och frambär den offergåva som Moses har påbjudit, till ett vittnesbörd för dem.»
När han därefter kom in i Kapernaum, trädde en hövitsman fram till honom och bad honom
och sade: »Herre, min tjänare ligger därhemma lam och lider svårt.»
Han sade till honom: »Skall då jag komma och bota honom?»
Hövitsmannen svarade och sade: »Herre, jag är icke värdig att du går in under mitt tak.
Men säg allenast ett ord, så bliver min tjänare frisk.
Jag är ju själv en man som står under andras befäl: jag har ock krigsmän under mig, och om jag säger till en av dem: 'Gå', så går han, eller till en annan: 'Kom', så kommer han; och om jag säger till min tjänare: 'Gör det', då gör han så.»
När Jesus hörde detta, förundrade han sig och sade till dem som följde honom: »Sannerligen säger jag eder: I Israel har jag icke hos någon funnit så stor tro.
Och jag säger eder: Många skola komma från öster och väster och få vara med Abraham, Isak och Jakob till bords i himmelriket,
men rikets barn skola bliva utkastade i mörkret därutanför; där skall vara gråt och tandagnisslan.»
Och Jesus sade till hövitsmannen: »Gå; såsom du tror, så må det ske dig.»
Och i samma stund blev tjänaren frisk.
När Jesus sedan kom in i Petrus' hus, fick han se hans svärmoder ligga sjuk i feber.
Då rörde han vid hennes hand, och febern lämnade henne; och hon stod upp och betjänade honom.
Men när det hade blivit afton, förde man till honom många som voro besatta; och han drev ut andarna med sitt blotta ord, och alla som voro sjuka botade han,
för att det skulle fullbordas, som var sagt genom profeten Esaias, när han sade: »Han tog på sig våra krankheter, och våra sjukdomar bar han.»
Då nu Jesus såg mycket folk omkring sig, bjöd han att man skulle fara över till andra stranden.
Och en skriftlärd kom fram och sade till honom: »Mästare, jag vill följa dig varthelst du går.»
Då svarade Jesus honom: »Rävarna hava kulor, och himmelens fåglar hava nästen; men Människosonen har ingen plats där han kan vila sitt huvud.»
Och en annan av hans lärjungar sade till honom: »Herre, tillstäd mig att först gå bort och begrava min fader.»
Då svarade Jesus honom: »Följ du mig, och låt de döda begrava sina döda.»
Och han steg i båten, och hans lärjungar följde honom.
Och se, då uppstod en häftig storm på sjön, så att vågorna slogo över båten; men han låg och sov.
Då gingo de fram och väckte honom och sade: »Herre, hjälp oss; vi förgås.»
Han sade till dem: »I klentrogne, varför rädens I?»
Därefter stod han upp och näpste vindarna och sjön, och det blev alldeles lugnt.
Och människorna förundrade sig och sade: »Vad är denne för en, eftersom både vindarna och sjön äro honom lydiga?»
När han så hade kommit över till gadarenernas land på andra stranden, kommo två besatta emot honom, ut från gravarna där.
Och de voro mycket våldsamma, så att ingen kunde färdas den vägen fram.
Dessa ropade då och sade: »Vad har du med oss att göra, du Guds Son?
Har du kommit hit för att plåga oss, förrän tid är?»
Nu gick där långt ifrån dem en stor svinhjord i bet.
Och de onda andarna bådo honom och sade: »Om du vill driva ut oss så låt oss fara in i svinhjorden.»
Då sade han till dem: »Faren åstad.»
Och de gåvo sig åstad och foro in i svinen.
Och se, då störtade sig hela hjorden utför branten ned i sjön och omkom i vattnet.
Men herdarna flydde; och när de hade kommit in i staden, omtalade de alltsammans, och särskilt vad som hade skett med de besatta.
Då gick hela staden ut för att möta Jesus; och när de fingo se honom, bådo de att han skulle begiva sig bort ifrån deras område.
Och han steg i en båt och for över och kom till sin egen stad.
Då förde de till honom en lam man, som låg på en säng.
När Jesus såg deras tro sade han till den lame: »Var vid gott mod, min son; dina synder förlåtas dig.»
Då sade några av de skriftlärde vid sig själva: »Denne hädar.»
Men Jesus förstod deras tankar och sade: »Varför tänken I i edra hjärtan vad ont är?
Vilket är lättare, att säga: 'Dina synder förlåtas dig' eller att säga: 'Stå upp och gå'?
Men för att I skolen veta att Människosonen har makt här på jorden att förlåta synder, så stå upp» -- sade han nu till den lame -- »och tag din säng och gå hem.»
Då stod han upp och gick hem.
När folket såg detta, blevo de häpna och prisade Gud, som hade givit sådan makt åt människor.
När Jesus därifrån gick vidare fram, fick han se en man, som hette Matteus, sitta vid tullhuset.
Och han sade till denne: »Följ mig.»
Då stod han upp och följde honom.
När han därefter låg till bords i hans hus, kommo många publikaner och syndare dit och voro bordsgäster där, jämte Jesus och hans lärjungar.
Men då fariséerna sågo detta, sade de till hans lärjungar: »Huru kan eder mästare äta med publikaner och syndare?»
När han hörde detta, sade han: »Det är icke de friska som behöva läkare, utan de sjuka.
Men gån I åstad och lären eder vad de orden betyda: 'Jag har behag till barmhärtighet, och icke till offer.'
Ty jag har icke kommit för att kalla rättfärdiga, utan för att kalla syndare.»
Därefter kommo Johannes' lärjungar till honom och sade: »Varför fasta icke dina lärjungar då vi och fariséerna ofta fasta?»
Jesus svarade dem: »Icke kunna väl bröllopsgästerna sörja, så länge brudgummen är hos dem?
Men den tid skall komma, då brudgummen tages ifrån dem, och då skola de fasta. --
Ingen sätter en lapp av okrympt tyg på en gammal mantel, ty det isatta stycket skulle riva bort ännu mer av manteln, och hålet skulle bliva värre.
Ej heller slår man nytt vin I gamla skinnläglar; om någon så gjorde, skulle läglarna sprängas sönder och vinet spillas ut, jämte det att läglarna fördärvades.
Nej, man slår nytt vin i nya läglar, så bliva båda delarna bevarade.»
Medan han talade detta till dem, trädde en synagogföreståndare fram och föll ned för honom och sade: »Min dotter har just nu dött, men kom och lägg din hand på henne, så bliver hon åter levande.»
Då stod Jesus upp och följde honom med sina lärjungar.
Men en kvinna, som i tolv år hade lidit av blodgång, närmade sig honom bakifrån och rörde vid hörntofsen på hans mantel.
Ty hon sade vid sig själv: »Om jag allenast får röra vid hans mantel, så bliver jag hulpen.»
Då vände Jesus sig om, och när han fick se henne, sade han: »Var vid gott mod, min dotter; din tro har hjälpt dig.»
Och kvinnan var hulpen från den stunden.
När Jesus sedan kom in i föreståndarens hus och fick se flöjtblåsarna och folket som höjde klagolåt,
sade han: »Gån bort härifrån; ty flickan är icke död, hon sover.»
Då hånlogo de åt honom.
Men sedan folket hade blivit utvisat, gick han in och tog flickan vid handen.
Då stod hon upp.
Och ryktet härom gick ut över hela det landet.
När Jesus gick därifrån, följde honom två blinda som ropade och sade: »Davids son, förbarma dig över oss.»
Och då han kom hem, trädde de blinda fram till honom; och Jesus frågade dem: »Tron I att jag kan göra detta?»
De svarade honom: »Ja, Herre.»
Då rörde han vid deras ögon och sade: »Ske eder efter eder tro.»
Och deras ögon öppnades.
Och Jesus tillsade dem strängeligen att se till, att ingen finge veta detta.
Men de gingo åstad och utspridde ryktet om honom över hela det landet.
När dessa voro på väg ut, förde man till honom en dövstum som var besatt.
Och när den onde anden hade blivit utdriven, talade den dövstumme.
Och folket förundrade sig och sade: »Sådant har aldrig förut varit sett i Israel.»
Men fariséerna sade: »Det är med de onda andarnas furste som han driver ut de onda andarna.»
Och Jesus gick omkring i alla städer och byar och undervisade i deras synagogor och predikade evangelium om riket och botade alla slags sjukdomar och allt slags skröplighet.
Och när han såg folkskarorna, ömkade han sig över dem, eftersom de voro så illa medfarna och uppgivna, »lika får som icke hava någon herde.»
Därför sade han till sina lärjungar: »Skörden är mycken, men arbetarna äro få.
Bedjen fördenskull skördens Herre att han sänder ut arbetare till sin skörd.»
Och han kallade till sig sina tolv lärjungar och gav dem makt över orena andar, till att driva ut dem, så ock makt att bota alla slags sjukdomar och allt slags skröplighet.
Och dessa äro de tolv apostlarnas namn: först Simon, som kallas Petrus, och Andreas, hans broder; vidare Jakob, Sebedeus' son, och Johannes, hans broder;
Filippus och Bartolomeus; Tomas och Matteus, publikanen; Jakob, Alfeus' son, och Lebbeus;
Simon ivraren och Judas Iskariot, densamme som förrådde honom.
Dessa tolv sände Jesus ut; och han bjöd dem och sade: »Ställen icke eder färd till hedningarna, och gån icke in i någon samaritisk stad,
utan gån hellre till de förlorade fåren av Israels hus.
Och där I gån fram skolen I predika och säga: 'Himmelriket är nära.'
Boten sjuka, uppväcken döda, gören spetälska rena, driven ut onda andar.
I haven fått för intet; så given ock för intet.
Skaffen eder icke guld eller silver eller koppar i edra bälten,
icke någon ränsel för eder färd, ej heller dubbla livklädnader, ej heller skor eller stav; ty arbetaren är värd sin mat.
Men när I haven kommit in i någon stad eller by, så utforsken vilken därinne som är värdig, och stannen hos honom, till dess I lämnen den orten.
Och när I kommen in i ett hus, så hälsen det.
Om då det huset är värdigt, så må den frid I tillönsken det komma däröver; men om det icke är värdigt, då må den frid I tillönsken det vända tillbaka till eder.
Och om man på något ställe icke tager emot eder och icke hör på edra ord, så gån ut ur det huset eller den staden, och skudden stoftet av edra fötter.
Sannerligen säger jag eder: För Sodoms och Gomorras land skall det på domens dag bliva drägligare än för den staden.
Se, jag sänder eder åstad såsom får mitt in ibland ulvar.
Varen fördenskull kloka såsom ormar och menlösa såsom duvor.
Tagen eder till vara för människorna; ty de skola draga eder inför domstolar, och i sina synagogor skola de gissla eder;
och I skolen föras fram också inför landshövdingar och konungar, för min skull, till ett vittnesbörd för dem och för hedningarna.
Men när man drager eder inför rätta, gören eder då icke bekymmer för huru eller vad I skolen tala; ty vad I skolen tala skall bliva eder givet i den stunden.
Det är icke I som skolen tala, utan det är eder Faders Ande som skall tala i eder.
Och den ene brodern skall då överlämna den andre till att dödas, ja ock fadern sitt barn; och barn skola sätta sig upp mot sina föräldrar och skola döda dem.
Och I skolen bliva hatade av alla, för mitt namns skull.
Men den som är ståndaktig intill änden, han skall bliva frälst. --
När de nu förfölja eder i en stad, så flyn till en annan; och om de också där förfölja eder, så flyn till ännu en annan.
Ty sannerligen säger jag eder: I skolen icke hava hunnit igenom alla Israels städer, förrän Människosonen kommer.
Lärjungen är icke förmer än sin mästare, ej heller är tjänaren förmer än sin herre.
Det må vara lärjungen nog, om det går honom såsom hans mästare, och tjänaren, om det går honom såsom hans herre.
Om de hava kallat husbonden för Beelsebul, huru mycket mer skola de icke så kalla hans husfolk!
Frukten alltså icke för dem; ty intet är förborgat, som icke skall bliva uppenbarat, och intet är fördolt, som icke skall bliva känt.
Vad jag säger eder i mörkret, det skolen säga i ljuset, och vad I hören viskas i edert öra, det skolen I predika på taken.
Och frukten icke för dem som väl kunna dräpa kroppen, men icke hava makt att dräpa själen, utan frukten fastmer honom som har makt att förgöra både själ och kropp i Gehenna. --
Säljas icke två sparvar för en skärv?
Och icke en av dem faller till jorden utan eder Faders vilja.
Men på eder äro till och med huvudhåren allasammans räknade.
Frukten alltså icke; I ären mer värda än många sparvar.
Därför, var och en som bekänner mig inför människorna, honom skall ock jag kännas vid inför min Fader, som är i himmelen.
Men den som förnekar mig inför människorna, honom skall ock jag förneka inför min Fader, som är i himmelen.
I skolen icke mena att jag har kommit för att sända frid på jorden.
Jag har icke kommit för att sända frid, utan svärd.
Ja, jag har kommit för att uppväcka söndring, så att 'sonen sätter sig upp mot sin fader och dottern mot sin moder och sonhustrun mot sin svärmoder,
och envar får sitt eget husfolk till fiender'.
Den som älskar fader eller moder mer än mig, han är mig icke värdig, och den som älskar son eller dotter mer än mig, han är mig icke värdig;
och den som icke tager sitt kors på sig och efterföljer mig, han är mig icke värdig.
Den som finner sitt liv, han skall mista det, och den som mister sitt liv, för min skull, han skall finna det. --
Den som tager emot eder, han tager emot mig, och den som tager emot mig, han tager emot honom som har sänt mig.
Den som tager emot en profet, därför att det är en profet, han skall få en profets lön; och den som tager emot en rättfärdig man, därför att det är en rättfärdig man, han skall få en rättfärdig mans lön.
Och den som giver en av dessa små allenast en bägare friskt vatten att dricka, därför att det är en lärjunge -- sannerligen säger jag eder: Han skall ingalunda gå miste om sin lön.»
När Jesus hade givit sina tolv lärjungar alla dessa bud, gick han därifrån vidare, för att undervisa och predika i deras städer.
Men när Johannes i sitt fängelse fick höra om Kristi gärningar, sände han bud med sina lärjungar
och lät fråga honom: »Är du den som skulle komma, eller skola vi förbida någon annan?»
Då svarade Jesus och sade till dem: »Gån tillbaka och omtalen för Johannes vad I hören och sen:
blinda få sin syn, halta gå, spetälska bliva rena, döva höra, döda uppstå, och 'för fattiga förkunnas glädjens budskap'.
Och salig är den för vilken jag icke bliver en stötesten.»
När dessa sedan gingo bort, begynte Jesus tala till folket om Johannes: »Varför var det I gingen ut i öknen?
Var det för att se ett rör som drives hit och dit av vinden?
Eller varför gingen I ut?
Var det för att se en människa klädd i fina kläder?
De som bära fina kläder, dem finnen I ju i konungapalatsen.
Varför gingen I då ut?
Var det för att se en profet?
Ja, jag säger eder: Ännu mer än en profet är han.
Han är den om vilken det är skrivet: 'Se, jag sänder ut min ängel framför dig, och han skall bereda vägen för dig.'
Sannerligen säger jag eder: Bland dem som äro födda av kvinnor har ingen uppstått, som har varit större än Johannes döparen; men den som är minst i himmelriket är likväl större än han.
Och från Johannes döparens dagar intill denna stund tränger himmelriket fram med storm, och människor storma fram och rycka det till sig.
Ty alla profeterna och lagen hava profeterat intill Johannes;
och om I viljen tro det: han är Elias, den som skulle komma.
Den som har öron, han höre.
Men vad skall jag likna detta släkte vid?
Det är likt barn som sitta på torgen och ropa till andra barn
och säga: 'Vi hava spelat för eder, och I haven icke dansat; vi hava sjungit sorgesång, och I haven icke jämrat eder.'
Ty Johannes kom, och han varken äter eller dricker, och så säger man: 'Han är besatt av en ond ande.'
Människosonen kom, och han både äter och dricker, och nu säger man: 'Se vilken frossare och vindrinkare han är, en publikaners och syndares vän!'
Men Visheten har fått rätt av sina barn.»
Därefter begynte han tala bestraffande ord till de städer i vilka han hade utfört så många av sina kraftgärningar, och förehålla dem att de icke hade gjort bättring:
»Ve dig, Korasin!
Ve dig, Betsaida!
Ty om de kraftgärningar som äro gjorda i eder hade blivit gjorda i Tyrus och Sidon, så skulle de för länge sedan hava gjort bättring i säck och aska.
Men jag säger eder: För Tyrus och Sidon skall det på domens dag bliva drägligare än för eder.
Och du, Kapernaum, skall väl du bliva upphöjt till himmelen?
Nej, ned till dödsriket måste du fara.
Ty om de kraftgärningar som äro gjorda i dig hade blivit gjorda i Sodom, så skulle det hava stått ännu i dag.
Men jag säger eder att det för Sodoms land skall på domens dag bliva drägligare än för dig.»
Vid den tiden talade Jesus och sade: »Jag prisar dig, Fader, du himmelens och jordens Herre, för att du väl har dolt detta för de visa och kloka, men uppenbarat det för de enfaldiga.
Ja, Fader; så har ju varit ditt behag.
Allt har av min Fader blivit förtrott åt mig.
Och ingen känner Sonen utom Fadern, ej heller känner någon Fadern utom Sonen och den för vilken Sonen vill göra honom känd. --
Kommen till mig, I alla som arbeten och ären betungade, så skall jag giva eder ro.
Tagen på eder mitt ok och lären av mig, ty jag är saktmodig och ödmjuk i hjärtat; 'så skolen I finna ro för edra själar'.
Ty mitt ok är milt, och min börda är lätt.»
Vid den tiden tog Jesus på sabbaten vägen genom ett sädesfält; och hans lärjungar blevo hungriga och begynte rycka av ax och äta.
När fariséerna sågo detta, sade de till honom: »Se, dina lärjungar göra vad som icke är lovligt att göra på en sabbat.»
Han svarade dem: »Haven I icke läst vad David gjorde, när han och de som följde honom blevo hungriga:
huru han då gick in i Guds hus, och huru de åto skådebröden, fastän det ju varken för honom eller för dem som följde honom var lovligt att äta sådant bröd, utan allenast för prästerna?
Eller haven I icke läst i lagen att prästerna på sabbaten bryta sabbaten i helgedomen, och likväl äro utan skuld?
Men jag säger eder: Här är vad som är förmer än helgedomen.
Och haden I förstått vad det är: 'Jag har behag till barmhärtighet, och icke till offer', så skullen I icke hava dömt dem skyldiga, som äro utan skuld.
Ty Människosonen är herre över sabbaten.»
Och han gick därifrån vidare och kom in i deras synagoga.
Och se, där var en man som hade en förvissnad hand.
Då frågade de honom och sade: »Är det lovligt att bota sjuka på sabbaten?»
De ville nämligen få något att anklaga honom för.
Men han sade till dem: »Om någon bland eder har ett får, och detta på sabbaten faller i en grop, fattar han icke då i det och drager upp det?
Huru mycket mer värd är nu icke en människa än ett får!
Alltså är det lovligt att på sabbaten göra vad gott är.»
Därefter sade han till mannen: »Räck ut din hand.»
Och han räckte ut den, och den blev frisk igen och färdig såsom den andra. --
Då gingo fariséerna bort och fattade det beslutet om honom, att de skulle förgöra honom.
Men när Jesus fick veta detta, gick han bort därifrån; och många följde honom, och han botade dem alla,
men förbjöd dem strängeligen att utbreda ryktet om honom.
Ty det skulle fullbordas, som var sagt genom profeten Esaias, när han sade:
»Se, över min tjänare, som jag har utvalt, min älskade, i vilken min själ har funnit behag, över honom skall jag låta min Ande komma, och han skall förkunna rätten bland folken.
Han skall icke kiva eller skria, och hans röst skall man icke höra på gatorna,
Ett brutet rör skall han icke sönderkrossa, och en rykande veke skall han icke utsläcka, intill dess att han har fört rätten fram till seger.
Och till hans namn skola folken sätta sitt hopp.»
Då förde man till honom en besatt, som var blind och dövstum.
Och han botade honom, så att den dövstumme talade och såg.
Och allt folket uppfylldes av häpnad och sade: »Månne icke denne är Davids son?»
Men när fariséerna hörde detta, sade de: »Det är allenast med Beelsebul, de onda andarnas furste, som denne driver ut de onda andarna.»
Men han förstod deras tankar och sade till dem: »Vart rike som har kommit i strid med sig självt bliver förött, och intet samhälle eller hus som har kommit i strid med sig självt kan hava bestånd.
Om nu Satan driver ut Satan, så har han kommit i strid med sig själv.
Huru kan då hans rike hava bestånd?
Och om det är med Beelsebul som jag driver ut de onda andarna, med vem driva då edra egna anhängare ut dem?
De skola alltså vara edra domare.
Om det åter är med Guds Ande som jag driver ut de onda andarna, så har ju Guds rike kommit till eder. --
Eller huru kan någon gå in i en stark mans hus och beröva honom hans bohag, såframt han icke förut har bundit den starke?
Först därefter kan han plundra hans hus.
Den som icke är med mig, han är emot mig, och den som icke församlar med mig, han förskingrar.
Därför säger jag eder: All annan synd och hädelse skall bliva människorna förlåten, men hädelse mot Anden skall icke bliva förlåten.
Ja, om någon säger något mot Människosonen, så skall det bliva honom förlåtet; men om någon säger något mot den helige Ande, så skall det icke bliva honom förlåtet, varken i denna tidsåldern eller i den tillkommande.
I måsten döma så: antingen är trädet gott, och då måste dess frukt vara god; eller är trädet dåligt, och då måste dess frukt vara dålig.
Ty av frukten känner man trädet.
I huggormars avföda, huru skullen I kunna tala något gott, då I själva ären onda?
Vad hjärtat är fullt av, det talar ju munnen.
En god människa bär ur sitt goda förråd fram vad gott är, och en ond människa bär ur sitt onda förråd fram vad ont är.
Men jag säger eder, att för vart fåfängligt ord som människorna tala skola de göra räkenskap på domens dag.
Ty efter dina ord skall du dömas rättfärdig, och efter dina ord skall du dömas skyldig.»
Då togo några av de skriftlärde och fariséerna till orda och sade till honom: »Mästare, vi skulle vilja se något tecken av dig.»
Men han svarade och sade till dem: »Ett ont och trolöst släkte är detta!
Det åstundar ett tecken, men intet annat tecken skall givas det än profeten Jonas' tecken.
Ty likasom Jonas tre dagar och tre nätter var i den stora fiskens buk, så skall ock Människosonen tre dagar och tre nätter vara i jordens sköte.
Ninevitiska män skola vid domen träda fram tillsammans med detta släkte och bliva det till dom.
Ty de gjorde bättring vid Jonas' predikan; och se, här är vad som är mer än Jonas.
Drottningen av Söderlandet skall vid domen träda fram tillsammans med detta släkte och bliva det till dom.
Ty hon kom från jordens ända för att höra Salomos visdom; och se, här är vad som är mer än Salomo.
När en oren ande har farit ut ur en människa, vandrar han omkring i ökentrakter och söker efter ro, men finner ingen.
Då säger han: 'Jag vill vända tillbaka till mitt hus, som jag gick ut ifrån.'
Och när han kommer dit och finner det stå ledigt och vara fejat och prytt,
då går han åstad och tager med sig sju andra andar, som äro värre än han själv, och de gå ditin och bo där; och så bliver för den människan det sista värre än det första.
Så skall det ock gå med detta onda släkte.»
Medan han ännu talade till folket, kommo hans moder och hans bröder och stannade därutanför och ville tala med honom.
Då sade någon till honom: »Se, din moder och dina bröder stå härutanför och vilja tala med dig.»
Men han svarade och sade till den som omtalade detta för honom: »Vilken är min moder, och vilka äro mina bröder?»
Och han räckte ut handen mot sina lärjungar och sade: »Se här är min moder, och här äro mina bröder!
Ty var och en som gör min himmelske Faders vilja, den är min broder och min syster och min moder.»
Samma dag gick Jesus ut från huset där han bodde och satte sig vid sjön.
Då församlade sig mycket folk omkring honom.
Därför steg han i en båt; och han satt i den, medan allt folket stod på stranden.
Och han talade till dem mycket i liknelser; han sade: »En såningsman gick ut för att så.
Och när han sådde, föll somt vid vägen, och fåglarna kommo och åto upp det.
Och somt föll på stengrund, där det icke hade mycket jord, och det kom strax upp, eftersom det icke hade djup jord;
men när solen hade gått upp, förbrändes det, och eftersom det icke hade någon rot, torkade det bort.
Och somt föll bland törnen, och törnena sköto upp och förkvävde det.
Men somt föll i god jord, och det gav frukt, dels hundrafalt, dels sextiofalt, dels trettiofalt.
Den som har öron, han höre.»
Då trädde lärjungarna fram och sade till honom: »Varför talar du till dem i liknelser?»
Han svarade och sade: »Eder är givet att lära känna himmelrikets hemligheter, men dem är det icke givet.
Ty den som har, åt honom skall varda givet, så att han får över nog; men den som icke har, från honom skall tagas också det han har.
Därför talar jag till dem i liknelser, eftersom de med seende ögon intet se, och med hörande öron intet höra, och intet heller förstå.
Så fullbordas på dem Esaias' profetia, den som säger: 'Med hörande öron skolen I höra, och dock alls intet förstå, och med seende ögon skolen I se, och dock alls intet förnimma.
Ty detta folks hjärta har blivit förstockat, och med öronen höra de illa, och sina ögon hava de tillslutit, så att de icke se med sina ögon, eller höra med sina öron, eller förstå med sina hjärtan, och omvända sig och bliva helade av mig.
Men saliga äro edra ögon, som se, och edra öron, som höra.
Ty sannerligen säger jag eder: Många profeter och rättfärdiga män åstundade att se det som I sen, men fingo dock icke se det, och att höra det som I hören, men fingo dock icke höra det.
Hören alltså I vad som menas med liknelsen om såningsmannen.
När någon hör ordet om riket, men icke förstår det, då kommer den onde och river bort det som såddes i hans hjärta.
Om en sådan människa kan det sägas att säden såddes vid vägen.
Och att den såddes på stengrunden, det är sagt om den som väl hör ordet och strax tager emot det med glädje,
men som icke har någon rot i sig, utan bliver beståndande allenast till en tid, och när bedrövelse eller förföljelse påkommer för ordets skull, då kommer han strax på fall.
Och att den såddes bland törnena, det är sagt om den som väl hör ordet, men låter tidens omsorger och rikedomens bedrägliga lockelse förkväva det, så att han bliver utan frukt.
Men att den såddes i den goda jorden, det är sagt om den som både hör ordet och förstår det, och som jämväl bär frukt och giver dels hundrafalt, dels sextiofalt, dels trettiofalt.»
En annan liknelse framställde han för dem; han sade: »Med himmelriket är det, såsom när en man sådde god säd i sin åker;
men när folket sov, kom hans ovän och sådde ogräs mitt ibland vetet och gick sedan sin väg.
När nu säden sköt upp och satte frukt, så visade sig ock ogräset.
Då trädde husbondens tjänare fram och sade till honom: 'Herre, du sådde ju god säd i din åker; varifrån har den då fått ogräs?
Han svarade dem: 'En ovän har gjort detta.'
Tjänarna sade till honom: 'Vill du alltså att vi skola gå åstad och samla det tillhopa?'
Men han svarade: 'Nej; ty då kunden I rycka upp vetet jämte ogräset, när I samlen detta tillhopa.
Låten båda slagen växa tillsammans intill skördetiden; och när skördetiden är inne, vill jag säga till skördemännen: 'Samlen först tillhopa ogräset, och binden det i knippor till att brännas upp, och samlen sedan in vetet i min lada.'»
En annan liknelse framställde han för dem; han sade: »Himmelriket är likt ett senapskorn som en man tager och lägger ned i sin åker.
Det är minst av alla frön, men när det har växt upp, är det störst bland kryddväxter; ja, det bliver ett träd, så att himmelens fåglar komma och bygga sina nästen på dess grenar.»
En annan liknelse framställde han för dem: »Himmelriket är likt en surdeg som en kvinna tager och blandar in i tre skäppor mjöl, till dess alltsammans bliver syrat.»
Allt detta talade Jesus i liknelser till folket, och utan liknelser talade han intet till dem.
Ty det skulle fullbordas, som var sagt genom profeten som sade: »Jag vill öppna min mun till liknelser, uppenbara vad förborgat har varit från världens begynnelse.»
Därefter lät han folket gå och gick själv hem.
Och hans lärjungar trädde fram till honom och sade: »Uttyd för oss liknelsen om ogräset i åkern.»
Han svarade och sade: »Den som sår den goda säden är Människosonen.
Åkern är världen.
Den goda säden, det är rikets barn, men ogräset är ondskans barn.
Ovännen, som sådde det, är djävulen.
Skördetiden är tidens ände.
Skördemännen är änglar.
Såsom nu ogräset samlas tillhopa och brännes upp i eld, så skall det ock ske vid tidens ände.
Människosonen skall då sända ut sina änglar, och de skola samla tillhopa och föra bort ur hans rike alla dem som äro andra till fall, och dem som göra vad orätt är,
och skola kasta dem i den brinnande ugnen; där skall vara gråt och tandagnisslan.
Då skola de rättfärdiga lysa såsom solen, i sin Faders rike.
Den som har öron, han höre.
Himmelriket är likt en skatt som har blivit gömd i en åker.
Och en man finner den, men håller det hemligt; och i sin glädje går han bort och säljer allt vad han äger och köper den åkern.
Ytterligare är det med himmelriket, såsom när en köpman söker efter goda pärlor;
och då han har funnit en dyrbar pärla, går han bort och säljer vad han äger och köper den.
Ytterligare är det med himmelriket, såsom när en not kastas i havet och samlar tillhopa fiskar av alla slag.
När den så bliver full, drager man upp den på stranden och sätter sig ned och samlar de goda i kärl, men de dåliga kastar man bort. --
Så skall det ock ske vid tidens ände: änglarna skola gå ut och skilja de onda från de rättfärdiga
och kasta dem i den brinnande ugnen; där skall vara gråt och tandagnisslan.
Haven I förstått allt detta?»
De svarade honom: »Ja.»
Då sade han till dem: »Så är nu var skriftlärd, som har blivit en lärjunge för himmelriket, lik en husbonde som ur sitt förråd bär fram nytt och gammalt.»
När Jesus hade framställt alla dessa liknelser, drog han bort därifrån.
Och han kom till sin fädernestad, och där undervisade han folket i deras synagoga, så att de häpnade och sade: »Varifrån har han fått denna vishet?
Och hans kraftgärningar, varifrån komma de?
Är då denne icke timmermannens son?
Heter icke hans moder Maria, och heta icke hans bröder Jakob och Josef och Simon och Judas?
Och hans systrar, bo de icke alla hos oss?
Varifrån har han då fått allt detta?»
Så blev han för dem en stötesten.
Men Jesus sade till dem: »En profet är icke föraktad utom i sin fädernestad och i sitt eget hus.»
Och för deras otros skull gjorde han där icke många kraftgärningar.
Vid den tiden fick Herodes, landsfursten, höra ryktet om Jesus.
Då sade han till sina tjänare: »Det är Johannes döparen.
Han har uppstått från de döda, och därför verka dessa krafter i honom.»
Herodes hade nämligen låtit gripa Johannes och binda honom och sätta honom i fängelse, för Herodias', sin broder Filippus' hustrus, skull.
Ty Johannes hade sagt till honom: »Det är icke lovligt för dig att hava henne.»
Och han hade velat döda honom, men han fruktade för folket, eftersom de höllo honom för en profet.
Men så kom Herodes' födelsedag.
Då dansade Herodias' dotter inför dem; och hon behagade Herodes så mycket,
att han med en ed lovade att giva henne vad helst hon begärde.
Hon sade då, såsom hennes moder ingav henne: »Giv mig här på ett fat Johannes döparens huvud.»
Då blev konungen bekymrad, men för edens och för bordsgästernas skull bjöd han att man skulle giva henne det,
och sände åstad och lät halshugga Johannes i fängelset.
Och hans huvud blev framburet på ett fat och givet åt flickan; och hon bar det till sin moder.
Men hans lärjungar kommo och togo hans döda kropp och begrovo honom.
Sedan gingo de och omtalade det för Jesus.
Då Jesus hörde detta, for han i en båt därifrån bort till en öde trakt, där de kunde vara allena.
Men när folket fick höra härom, kommo de landvägen efter honom från städerna.
Och då han steg i land, fick han se att där var mycket folk; och han ömkade sig över dem och botade deras sjuka.
Men när det led mot aftonen, trädde hans lärjungar fram till honom och sade: »Trakten är öde, och tiden är redan framskriden.
Låt folket skiljas åt, så att de kunna gå bort i byarna och köpa sig mat.»
Men Jesus sade till dem: »De behöva icke gå bort; given I dem att äta.»
De svarade honom: »Vi hava här icke mer än fem bröd och två fiskar.»
Då sade han: »Bären dem hit till mig.»
Därefter tillsade han folket att lägga sig ned i gräset.
Och han tog de fem bröden och de två fiskarna och såg upp till himmelen och välsignade dem.
Och han bröt bröden och gav dem åt lärjungarna, och lärjungarna gåvo åt folket.
Och de åto alla och blevo mätta Sedan samlade man upp de överblivna styckena, tolv korgar fulla.
Men de som hade ätit voro vid pass fem tusen män, förutom kvinnor och barn.
Strax därefter nödgade han sina lärjungar att stiga i båten och före honom fara över till andra stranden, medan han tillsåg att folket skildes åt.
Och sedan detta hade skett, gick han upp på berget för att vara allena och bedja.
När det så hade blivit afton, var han där ensam.
Båten var då redan många stadier från land och hårt ansatt av vågorna, ty vinden låg emot.
Men under fjärde nattväkten kom Jesus till dem, gående fram över sjön.
När då lärjungarna fingo se honom gå på sjön, blevo de förfärade och sade: »Det är en vålnad», och ropade av förskräckelse.
Men Jesus begynte strax tala till dem och sade: »Varen vid gott mod; det är jag, varen icke förskräckta.»
Då svarade Petrus honom och sade: »Herre, är det du, så bjud mig att komma till dig på vattnet.»
Han sade: »Kom.»
Då steg Petrus ut ur båten och begynte gå på vattnet och kom till Jesus.
Men när han såg huru stark vinden var, blev han förskräckt; och då han nu begynte sjunka, ropade han och sade: »Herre, hjälp mig.»
Och strax räckte Jesus ut handen och fattade i honom och sade till honom: »Du klentrogne, varför tvivlade du?»
När de sedan hade kommit upp i båten, lade sig vinden.
Men de som voro i båten föllo ned för honom och sade: »Förvisso är du Guds Son.»
När de hade farit över, kommo de till Gennesarets land.
Då nu folket där på orten kände igen honom, sände de ut bud i hela trakten däromkring, och man förde till honom alla som voro sjuka.
Och de bådo honom att allenast få röra vid hörntofsen på hans mantel; och alla som rörde vid den blevo hulpna.
Härefter kommo fariséer och skriftlärde från Jerusalem till Jesus och sade:
»Varför överträda dina lärjungar de äldstes stadgar?
De två ju icke sina händer, när de skola äta.»
Men han svarade och sade till dem: »Varför överträden I själva Guds bud, för edra stadgars skull?
Gud har ju sagt: 'Hedra din fader och din moder' och: 'Den som smädar sin fader eller sin moder, han skall döden dö.'
Men I sägen, att om någon säger till sin fader eller sin moder: 'Vad du av mig kunde hava fått till hjälp, det giver jag i stället såsom offergåva', då behöver han alls icke hedra sin fader eller sin moder.
I haven så gjort Guds budord om intet, för edra stadgars skull.
I skrymtare, rätt profeterade Esaias om eder, när han sade:
'Detta folk ärar mig med sina läppar, men deras hjärtan äro långt ifrån mig;
och fåfängt dyrka de mig, eftersom de läror de förkunna äro människobud.'»
Och han kallade folket till sig och sade till dem: »Hören och förstån.
Icke vad som går in i munnen orenar människan, men vad som går ut ifrån munnen, det orenar människan.»
Då trädde hans lärjungar fram och sade till honom: »Vet du, att när fariséerna hörde det du nu sade, var det för dem en stötesten?»
Men han svarade och sade: »Var planta som min himmelske Fader icke har planterat skall ryckas upp med rötterna.
Frågen icke efter dem.
De äro blinda ledare; och om en blind leder en blind, så falla de båda i gropen.»
Då tog Petrus till orda och sade till honom: »Uttyd för oss detta bildliga tal.»
Han sade: »Ären då också I ännu utan förstånd?
Insen I icke att allt som går in i munnen, det går ned i buken och har sin naturliga utgång?
Men vad som går ut ifrån munnen, det kommer från hjärtat, och det är detta som orenar människan.
Ty från hjärtat komma onda tankar, mord, äktenskapsbrott, otukt, tjuveri, falskt vittnesbörd, hädelse.
Det är detta som orenar människan; men att äta med otvagna händer, det orenar icke människan.»
Och Jesus begav sig bort därifrån och drog sig undan till trakten av Tyrus och Sidon.
Då kom en kananeisk kvinna från det området och ropade och sade: »Herre, Davids son, förbarma dig över mig.
Min dotter plågas svårt av en ond ande.»
Men han svarade henne icke ett ord.
Då trädde hans lärjungar fram och bådo honom och sade: »Giv henne besked; hon förföljer oss ju med sitt ropande.»
Han svarade och sade: »Jag är icke utsänd till andra än till de förlorade fåren av Israels hus.»
Men hon kom fram och föll ned för honom och sade: »Herre, hjälp mig.»
Då svarade han och sade: »Det är otillbörligt att taga brödet från barnen och kasta det åt hundarna.»
Hon sade: »Ja, Herre.
Också äta ju hundarna allenast av de smulor som falla ifrån deras herrars bord.»
Då svarade Jesus och sade till henne: »O kvinna, din tro är stor.
Ske dig såsom du vill.»
Och hennes dotter var frisk ifrån den stunden.
Men Jesus gick därifrån vidare och kom till Galileiska sjön.
Och han gick upp på berget och satte sig där.
Då kom mycket folk till honom, och de hade med sig halta, blinda, dövstumma, lytta och många andra; dem lade de ned för hans fötter, och han botade dem,
så att folket förundrade sig, när de funno dövstumma tala, lytta vara friska och färdiga, halta gå och blinda se.
Och man prisade Israels Gud.
Och Jesus kallade sina lärjungar till sig och sade: »Jag ömkar mig över folket, ty det är redan tre dagar som de hava dröjt kvar hos mig, och de hava intet att äta; och jag vill icke låta dem gå ifrån mig fastande, för att de icke skola uppgivas på vägen.»
Då sade lärjungarna till honom: »Varifrån skola vi här, i en öken, få så mycket bröd, att vi kunna mätta så mycket folk?»
Jesus frågade dem: »Huru många bröd haven I?»
De svarade: »Sju, och därtill några få småfiskar.»
Då tillsade han folket att lägra sig på marken.
Och han tog de sju bröden, så ock fiskarna, och tackade Gud och bröt bröden och gav åt lärjungarna, och lärjungarna gåvo åt folket.
Så åto de alla och blevo mätta.
Och de överblivna styckena samlade man sedan upp, sju korgar fulla.
Men de som hade ätit voro fyra tusen män, förutom kvinnor och barn.
Sedan lät han folket skiljas åt och steg i båten och for till Magadans område.
Och fariséerna och sadducéerna kommo dit och ville sätta honom på prov; de begärde att han skulle låta dem se något tecken från himmelen.
Men han svarade och sade till dem: »Om aftonen sägen I: 'Det bliver klart väder, ty himmelen är röd',
och om morgonen: 'Det bliver oväder i dag, ty himmelen är mulen och röd.'
Ja, om himmelens utseende förstån I att döma, men om tidernas tecken kunnen I icke döma.
Ett ont och trolöst släkte är detta!
Det åstundar ett tecken, men intet annat tecken skall givas det än Jonas' tecken.»
Och så lämnade han dem och gick sin väg.
När sedan lärjungarna foro åstad, över till andra stranden, hade de förgätit att taga med sig bröd.
Och Jesus sade till dem: »Sen till, att I tagen eder till vara för fariséernas och sadducéernas surdeg.»
Då talade de med varandra och sade: »Det är därför att vi icke hava tagit med oss bröd.»
Men när Jesus märkte detta, sade han: »I klentrogne, varför talen I eder emellan om att I icke haven bröd med eder?
Förstån I ännu ingenting?
Och kommen I icke ihåg de fem bröden åt de fem tusen, och huru många korgar I då togen upp?
Ej heller de sju bröden åt de fyra tusen, och huru många korgar I då togen upp?
Huru kommer det då till, att I icke förstån att det ej var om bröd som jag talade till eder?
Tagen eder till vara för fariséernas och sadducéernas surdeg.»
Då förstodo de att det icke var för surdeg i bröd som han hade bjudit dem att taga sig till vara, utan för fariséernas och sadducéernas lära.
Men när Jesus kom till trakten av Cesarea Filippi, frågade han sina lärjungar och sade: »Vem säger folket Människosonen vara?»
De svarade: »Somliga säga Johannes döparen, andra Elias, andra åter Jeremias eller en annan av profeterna.»
Då frågade han dem: »Vem sägen då I mig vara?»
Simon Petrus svarade och sade: »Du är Messias, den levande Gudens Son.»
Då svarade Jesus och sade till honom: »Salig är du, Simon, Jonas' son; ty kött och blod har icke uppenbarat detta för dig, utan min Fader, som är i himmelen.
Så säger ock jag dig att du är Petrus; och på denna klippa skall jag bygga min församling, och dödsrikets portar skola icke bliva henne övermäktiga.
Jag skall giva dig himmelrikets nycklar: allt vad du binder på jorden, det skall vara bundet i himmelen; och allt vad du löser på jorden, det skall vara löst i himmelen.»
Därefter förbjöd han lärjungarna att för någon säga att han var Messias.
Från den tiden begynte Jesus förklara för sina lärjungar, att han måste gå till Jerusalem och lida mycket av de äldste och översteprästerna och de skriftlärde, och att han skulle bliva dödad, men att han på tredje dagen skulle uppstå igen.
Då tog Petrus honom avsides och begynte ivrigt motsäga honom och sade: »Bevare dig Gud, Herre!
Ingalunda får detta vederfaras dig.»
Men han vände sig om och sade till Petrus: »Gå bort, Satan, och stå mig icke i vägen; du är för mig en stötesten, ty dina tankar äro icke Guds tankar, utan människotankar.»
Därefter sade Jesus till sina lärjungar: »Om någon vill efterfölja mig, så försake han sig själv och tage sitt kors på sig: så följe han mig.
Ty den som vill bevara sitt liv, han skall mista det; men den som mister sitt liv, för min skull, han skall finna det.
Och vad hjälper det en människa, om hon vinner hela världen, men förlorar sin själ?
Eller vad kan en människa giva till lösen för sin själ?
Människosonen skall komma i sin Faders härlighet med sina änglar, och då skall han vedergälla var och en efter hans gärningar.
Sannerligen säger jag eder: Bland dem som här stå finnas några som icke skola smaka döden, förrän de få se Människosonen komma i sitt rike.»
Sex dagar därefter tog Jesus med sig Petrus och Jakob och Johannes, Jakobs broder, och förde dem upp på ett högt berg, där de voro allena.
Och hans utseende förvandlades inför dem: hans ansikte sken såsom solen, och hans kläder blevo vita såsom ljuset.
Och se, för dem visade sig Moses och Elias, i samtal med honom.
Då tog Petrus till orda och sade till Jesus: »Herre, här är oss gott att vara; vill du, så skall jag här göra tre hyddor, åt dig en och åt Moses en och åt Elias en.»
Och se, medan han ännu talade, överskyggade dem en ljus sky, och ur skyn kom en röst som sade: »Denne är min älskade Son, i vilken jag har funnit behag; hören honom.»
När lärjungarna hörde detta, föllo de ned på sina ansikten i stor förskräckelse.
Men Jesus gick fram och rörde vid dem och sade: »Stån upp, och varen icke förskräckta.»
När de då lyfte upp sina ögon, sågo de ingen utom Jesus allena.
Då de sedan gingo ned från berget, bjöd Jesus dem och sade: »Omtalen icke för någon denna syn, förrän Människosonen har uppstått från de döda.»
Men lärjungarna frågade honom och sade: »Huru kunna då de skriftlärde säga att Elias först måste komma?»
Han svarade och sade: »Elias måste visserligen komma och upprätta allt igen;
men jag säger eder att Elias redan har kommit.
Men de ville icke veta av honom, utan förforo mot honom alldeles såsom de ville.
Sammalunda skall ock Människosonen få lida genom dem.»
Då förstodo lärjungarna att det var om Johannes döparen som han talade till dem.
När de därefter kommo till folket, trädde en man fram till honom och föll på knä för honom
och sade: »Herre, förbarma dig över min son ty han är månadsrasande och plågas svårt; ofta faller han i elden och ofta i vattnet.
Och jag förde honom till dina lärjungar, men de kunde icke bota honom.»
Då svarade Jesus och sade: »O du otrogna och vrånga släkte, huru länge måste jag vara bland eder?
Huru länge måste jag härda ut med eder?
Fören honom hit till mig.»
Och Jesus tilltalade honom strängt, och den onde anden for ut ur honom; och gossen var botad från den stunden.
Sedan, när de voro allena, trädde lärjungarna fram till Jesus och frågade: »Varför kunde icke vi driva ut honom?»
Han svarade dem: »För eder otros skull.
Ty sannerligen säger jag eder: Om I haven tro, vore den ock blott såsom ett senapskorn, så skolen I kunna säga till detta berg: 'Flytta dig härifrån dit bort', och det skall flytta sig; ja, intet skall då vara omöjligt för eder.»
237910
Medan de nu tillsammans vandrade omkring i Galileen, sade Jesus till dem: »Människosonen skall bliva överlämnad i människors händer,
och man skall döda honom, men på tredje dagen skall han uppstå igen.»
Då blevo de mycket bedrövade.
Och när de hade kommit till Kapernaum, trädde de som uppburo tempelskatten fram till Petrus och sade: »Plägar icke eder mästare betala tempelskatt?»
Han svarade: »Jo.»
När han sedan hade kommit hem, förekom honom Jesus med frågan: »Vad synes dig, Simon?
Av vilka taga jordens konungar tull eller skatt, av sina söner eller av andra människor?»
Han svarade: »Av andra människor.»
Då sade Jesus till honom: »Alltså äro då sönerna fria.
Men för att vi icke skola bliva dem till en stötesten, så gå ned till sjön och kasta ut en krok.
Tag så den första fisk som du drager upp, och när du öppnar munnen på den skall du där finna en silverpenning.
Tag den, och giv den åt dem for mig och dig.»
I samma stund trädde lärjungarna fram till Jesus och frågade: »Vilken är den störste i himmelriket?»
Då kallade han fram ett barn och ställde det mitt ibland dem
och sade: »Sannerligen säger jag eder: Om I icke omvänden eder och bliven såsom barn, skolen I icke komma in i himmelriket.
Den som nu så ödmjukar sig, att han bliver såsom detta barn, han är den störste i himmelriket.
Och den som tager emot ett sådant barn I mitt namn, han tager emot mig.
Men den som förför en av dessa små som tro på mig, för honom vore det bättre att en kvarnsten hängdes om hans hals och han sänktes ned i havets djup.
Ve världen för förförelsers skull!
Förförelser måste ju komma; men ve den människa genom vilken förförelsen kommer!
Om nu din hand eller din fot är dig till förförelse, så hugg av den och kasta den ifrån dig.
Det är bättre för dig att ingå i livet lytt eller halt, än att hava båda händerna eller båda fötterna i behåll och kastas i den eviga elden.
Och om ditt öga är dig till förförelse, så riv ut det och kasta det ifrån dig.
Det är bättre för dig att ingå i livet enögd, än att hava båda ögonen i behåll och kastas i det brinnande Gehenna.
Sen till, att I icke förakten någon av dessa små; ty jag säger eder att deras änglar i himmelen alltid se min himmelske Faders ansikte.
238080
Vad synes eder?
Om en man har hundra får, och ett av dem har kommit vilse, lämnar han icke då de nittionio på bergen och går åstad och söker efter det som har kommit vilse?
Och händer det då att han finner det -- sannerligen säger jag eder: då gläder han sig mer över det fåret än över de nittionio som icke hade kommit vilse.
Så är det ej heller eder himmelske Faders vilja att någon av dessa små skall gå förlorad.
Men om din broder försyndar sig, så gå åstad och förehåll honom det enskilt.
Om han då lyssnar till dig, så har du vunnit din broder.
Men om han icke lyssnar till dig, så tag med dig ännu en eller två, för att 'var sak må avgöras efter två eller tre vittnens utsago'.
Lyssnar han icke till dem, så säg det till församlingen.
Lyssnar han ej heller till församlingen, så vare han för dig såsom en hedning och en publikan.
Sannerligen säger jag eder: Allt vad I binden på jorden, det skall vara bundet i himmelen; och allt vad I lösen på jorden, det skall vara löst i himmelen.
Ytterligare säger jag eder, att om två av eder här på jorden komma överens att bedja om något, vad det vara må, så skall det beskäras dem av min Fader, som är i himmelen.
Ty var två eller tre är församlade i mitt namn, där är jag mitt ibland dem.»
Då trädde Petrus fram och sade till honom: »Herre, huru många gånger skall jag förlåta min broder, om han försyndar sig mot mig?
Är sju gånger nog?»
Jesus svarade honom: »Jag säger dig: Icke sju gånger, utan sjuttio gånger sju gånger.
Alltså är det med himmelriket, såsom när en konung ville hålla räkenskap med sina tjänare.
Och när han begynte hålla räkenskap, förde man fram till honom en som var skyldig honom tio tusen pund.
Men då denna icke kunde betala, bjöd hans herre att han skulle säljas, så ock hans hustru och barn och allt vad han ägde, för att skulden måtte bliva betald.
Då föll tjänaren ned för hans fötter och sade: 'Hav tålamod med mig, så skall jag betala dig alltsammans.'
Och tjänarens herre ömkade sig över honom och gav honom fri och efterskänkte honom hans skuld.
Men när samme tjänare kom ut, träffade han på en av sina medtjänare, som var skyldig honom hundra silverpenningar; och han tog fast denne och grep honom vid strupen och sade: 'Betala vad du är skyldig.'
Då föll hans medtjänare ned och bad honom och sade: 'Hav tålamod med mig, så skall jag betala dig.'
Men han ville icke, utan gick åstad och lät sätta honom i fängelse, till dess han hade betalt vad han var skyldig.
Då nu hans medtjänare sågo det som skedde, togo de mycket illa vid sig och gingo och berättade för sin herre allt som hade skett.
Då kallade hans herre honom till sig och sade till honom: 'Du onde tjänare, allt vad du var skyldig efterskänkte jag dig, eftersom du bad mig därom.
Borde då icke också du hava förbarmat dig över din medtjänare, såsom jag förbarmade mig över dig?'
Och i sin vrede överlämnade hans herre honom i fångknektarnas våld, intill dess han hade betalt allt vad han var skyldig.
Så skall ock min himmelske Fader göra med eder, om I icke av hjärtat förlåten var och en sin broder.»
När Jesus hade slutat detta tal, drog han bort ifrån Galileen och begav sig, genom landet på andra sidan Jordan, till Judeens område.
Och mycket folk följde honom, och han botade där de sjuka.
Då ville några fariséer snärja honom och trädde fram till honom och sade: »Är det lovligt att skilja sig från sin hustru av vilken orsak som helst?»
Men han svarade och sade: »Haven I icke läst att Skaparen redan i begynnelsen 'gjorde dem till man och kvinna'
och sade: 'Fördenskull skall en man övergiva sin fader och sin moder och hålla sig till sin hustru, och de tu skola varda ett kött'?
Så äro de icke mer två, utan ett kött.
Vad nu Gud har sammanfogat, det må människan icke åtskilja.»
Då sade de till honom: »Huru kunde då Moses bjuda att man skulle giva hustrun skiljebrev och så skilja sig från henne?»
Han svarade dem: »För edra hjärtans hårdhets skull tillstadde Moses eder att skiljas från edra hustrur, men från begynnelsen har det icke varit så.
Och jag säger eder: Den som för någon annan orsaks skull än för otukt skiljer sig från sin hustru och tager sig en annan hustru, han begår äktenskapsbrott.»
Då sade lärjungarna till honom: »Är det så med mannens ställning till hustrun, då är det icke rådligt att gifta sig.»
Men han svarade dem: »Icke alla kunna taga emot det ordet, utan allenast de åt vilka sådant är givet.
Ty visserligen finnas somliga som genom födelsen, allt ifrån moderlivet, äro oskickliga till äktenskap, andra åter som av människor hava gjorts oskickliga därtill, men somliga finnas ock, som för himmelrikets skull självmant hava gjort sig oskickliga därtill.
Den som kan taga emot detta, han tage emot det.»
Därefter buros barn fram till honom, för att han skulle lägga händerna på dem och bedja; men lärjungarna visade bort dem.
Då sade Jesus: »Låten barnen vara, och förmenen dem icke att komma till mig; ty himmelriket hör sådana till.»
Och han lade händerna på dem och gick sedan därifrån.
Då trädde en man fram till honom och sade: »Mästare, vad gott skall jag göra för att få evigt liv?»
Han sade till honom: »Varför frågar du mig om vad som är gott?
En finnes som är god.
Men vill du ingå i livet, så håll buden.»
Han frågade: »Vilka?»
Jesus svarade: »'Du skall icke dräpa', 'Du skall icke begå äktenskapsbrott', 'Du skall icke stjäla', 'Du skall icke bära falskt vittnesbörd',
'Hedra din fader och din moder' och 'Du skall älska din nästa såsom dig själv.'»
Då sade den unge mannen till honom: »Allt detta har jag hållit.
Vad fattas mig ännu?»
Jesus svarade honom: »Vill du vara fullkomlig, så gå bort och sälj vad du äger och giv åt de fattiga; då skall du få en skatt i himmelen.
Och kom sedan och följ mig.»
Men när den unge mannen hörde detta, gick han bedrövad bort, ty han hade många ägodelar.
Då sade Jesus till sina lärjungar: »Sannerligen säger jag eder: För den som är rik är det svårt att komma in i himmelriket.
Ja, jag säger eder: Det är lättare för en kamel att komma in genom ett nålsöga, än för den som är rik att komma in i Guds rike.»
När lärjungarna hörde detta, blevo de mycket häpna och sade: »Vem kan då bliva frälst?»
Men Jesus såg på dem och sade till dem: »För människor är detta omöjligt, men för Gud är allting möjligt.»
Då tog Petrus till orda och sade till honom: »Se, vi hava övergivit allt och följt dig; vad skola vi få därför?»
Jesus svarade dem: »Sannerligen säger jag eder: När världen födes på nytt, då när Människosonen sätter sig på sin härlighets tron, då skolen också I, som haven efterföljt mig, få sitta på tolv troner såsom domare över Israels tolv stammar.
Och var och en som har övergivit hus, eller bröder eller systrar, eller fader eller moder, eller barn, eller jordagods, för mitt namns skull, han skall få mångfaldigt igen, och skall få evigt liv till arvedel.
Men många som äro de första skola bliva de sista, och många som äro de sista skola bliva de första.»
»Ty med himmelriket är det, såsom när en husbonde bittida om morgonen gick ut för att leja åt sig arbetare till sin vingård.
Och när han hade kommit överens med arbetarna om en viss dagspenning, sände han dem till sin vingård.
När han sedan gick ut vid tredje timmen, fick han se några andra stå sysslolösa på torget;
och han sade till dem: 'Gån ock I till min vingård, så skall jag giva eder vad skäligt är.'
Och de gingo.
Åter gick han ut vid sjätte timmen och vid nionde och gjorde sammalunda.
Också vid elfte timmen gick han ut och fann då några andra stå där; och han sade till dem: 'Varför stån I här hela dagen sysslolösa?'
De svarade honom: 'Därför att ingen har lejt oss.'
Då sade han till dem: 'Gån ock I till min vingård.'
När det så hade blivit afton, sade vingårdens herre till sin förvaltare: 'Kalla fram arbetarna och giv dem deras lön, men begynn med de sista och gå så tillbaka ända till de första.'
Då nu de kommo fram, som voro lejda vid elfte timmen, fick var och en av dem full dagspenning.
När sedan de första kommo, trodde de att de skulle få mer, men också var och en av dem fick samma dagspenning.
När de så fingo, knorrade de mot husbonden.
och sade: 'Dessa sista hava arbetat allenast en timme, och du har ändå ställt dem lika med oss, som hava burit dagens tunga och solens hetta?'
Då svarade han en av dem och sade: 'Min vän, jag gör dig ingen orätt.
Kom du icke överens med mig om den dagspenningen?
Tag vad dig tillkommer och gå.
Men åt denne siste vill jag giva lika mycket som åt dig.
Har jag icke lov att göra såsom jag vill med det som är mitt?
Eller skall du med onda ögon se på att jag är så god?' --
Så skola de sista bliva de första, och de första bliva de sista.»
Då nu Jesus ville gå upp till Jerusalem, tog han till sig de tolv, så att de voro allena; och under vägen sade han till dem:
»Se, vi gå nu upp till Jerusalem, och Människosonen skall bliva överlämnad åt översteprästerna och de skriftlärde, och de skola döma honom till döden
och överlämna honom åt hedningarna till att begabbas och gisslas och korsfästas; men på tredje dagen skall han uppstå igen.»
Då trädde Sebedeus' söners moder fram till honom med sina söner och föll ned för honom och ville begära något av honom.
Han frågade henne: »Vad vill du?»
Hon svarade honom: »Säg att i ditt rike den ene av dessa mina två söner skall få sitta på din högra sida, och den andre på din vänstra.»
Men Jesus svarade och sade: »I veten icke vad I begären.
Kunnen I dricka den kalk som jag skall dricka?»
De svarade honom: »Det kunna vi.»
Då sade han till dem: »Ja, väl skolen I få dricka min kalk, men platsen på min högra sida och platsen på min vänstra tillkommer det icke mig att bortgiva, utan de skola tillfalla dem för vilka så är bestämt av min Fader.»
När de tio andra hörde detta, blevo de misslynta på de två bröderna.
Då kallade Jesus dem till sig och sade: »I veten att furstarna uppträda mot sina folk såsom herrar, och att de mäktige låta folken känna sin myndighet.
Så är det icke bland eder; utan den som vill bliva störst bland eder, han vare de andras tjänare,
och den som vill vara främst bland eder, han vare de andras dräng,
likasom Människosonen har kommit, icke för att låta tjäna sig, utan för att tjäna och giva sitt liv till lösen för många.»
När de sedan gingo ut ifrån Jeriko, följde honom mycket folk.
Och se, två blinda sutto där vid vägen.
När dessa hörde att det var Jesus som gick där fram, ropade de och sade: »Herre, förbarma dig över oss, du Davids son.»
Och folket tillsade dem strängeligen att de skulle tiga; men de ropade dess mer och sade: »Herre, förbarma dig över oss, du Davids son.»
Då stannade Jesus och kallade dem till sig och sade: »Vad viljen I att jag skall göra eder?»
De svarade honom: »Herre, låt våra ögon bliva öppnade.»
Då förbarmade sig Jesus över dem och rörde vid deras ögon, och strax fingo de sin syn och följde honom.
När de nu nalkades Jerusalem och kommo till Betfage vid Oljeberget, då sände Jesus åstad två lärjungar
och sade till dem: »Gån in i byn som ligger mitt framför eder, så skolen I strax finna en åsninna stå där bunden och en fåle bredvid henne; lösen dem och fören dem till mig.
Och om någon säger något till eder, så skolen I svara: 'Herren behöver dem'; då skall han strax släppa dem.»
Detta har skett, för att det skulle fullbordas, som var sagt genom profeten som sade:
»Sägen till dottern Sion: 'Se, din konung kommer till dig, saktmodig, ridande på en åsna, på en arbetsåsninnas fåle.'»
Och lärjungarna gingo åstad och gjorde såsom Jesus hade befallt dem
och ledde till honom åsninnan och fålen; och de lade sina mantlar på denne, och han satte sig därovanpå.
Och folkskaran, som var mycket stor, bredde ut sina mantlar på vägen; men somliga skuro kvistar av träden och strödde på vägen.
Och folket, både de som gingo före honom och de som följde efter, ropade och sade: »Hosianna Davids son!
Välsignad vare han som kommer, i Herrens namn.
Hosianna i höjden!»
När han så drog in i Jerusalem, kom hela staden i rörelse, och man frågade: »Vem är denne?»
Och folket sade: »Det är Jesus, profeten, från Nasaret i Galileen.»
Och Jesus gick in i helgedomen.
Och han drev ut alla dem som sålde och köpte i helgedomen, och han stötte omkull växlarnas bord och duvomånglarnas säten.
Och han sade till dem: »Det är skrivet: 'Mitt hus skall kallas ett bönehus.'
Men I gören det till en rövarkula.»
Och blinda och halta kommo fram till honom i helgedomen, och han botade dem.
Men när översteprästerna och de skriftlärde sågo de under som han gjorde, och sågo barnen som ropade i helgedomen och sade: »Hosianna Davids son!», då förtröt detta dem;
och de sade till honom: »Hör du vad dessa säga?»
Då svarade Jesus dem: »Ja; haven I aldrig läst: 'Av barns och spenabarns mun har du berett dig lov'?»
Därefter lämnade han dem och gick ut ur staden till Betania och stannade där över natten.
När han sedan på morgonen gick in till staden igen, blev han hungrig.
Och då han fick se ett fikonträd vid vägen, gick han fram till det, men fann intet därpå, utom allenast löv.
Då sade han till det: »Aldrig någonsin mer skall frukt växa på dig.»
Och strax förtorkades fikonträdet.
När lärjungarna sågo detta, förundrade de sig och sade: »Huru kunde fikonträdet så i hast förtorkas?»
Då svarade Jesus och sade till dem: »Sannerligen säger jag eder: Om I haven tro och icke tvivlen, så skolen I icke allenast kunna göra sådant som skedde med fikonträdet, utan I skolen till och med kunna säga till detta berg: 'Häv dig upp och kasta dig i havet', och det skall ske.
Och allt vad I med tro bedjen om i eder bön, det skolen I få.»
När han därefter hade kommit in i helgedomen, trädde översteprästerna och folkets äldste fram till honom, där han undervisade; och de sade: »Med vad myndighet gör du detta?
Och vem har givit dig sådan myndighet?»
Jesus svarade och sade till dem: »Också jag vill ställa en fråga till eder; om I svaren mig på den, så skall ock jag säga eder med vad myndighet jag gör detta».
Johannes' döpelse, varifrån var den: från himmelen eller från människor?»
Då överlade de med varandra och sade: »Om vi svara: 'Från himmelen', så frågar han oss: 'Varför trodden I honom då icke?'
Men om vi svara: 'Från människor', då måste vi frukta för folket, ty alla hålla de Johannes för en profet.»
De svarade alltså Jesus och sade: »Vi veta det icke.»
Då sade ock han till dem: »Så säger icke heller jag eder med vad myndighet jag gör detta.
Men vad synes eder?
En man hade två söner.
Och han kom till den förste och sade: 'Min son, gå i dag och arbeta i vingården.'
Han svarade och sade: 'Jag vill icke'; men efteråt ångrade han sig och gick.
Och han kom till den andre och sade sammalunda.
Då svarade denne och sade: 'Ja, herre'; men han gick icke,
Vilken av de två gjorde vad fadern ville?»
De svarade: »Den förste.»
Jesus sade till dem: »Ja, sannerligen säger jag eder: Publikaner och skökor skola förr gå in i Guds rike än I.
Ty Johannes kom och lärde eder rättfärdighetens väg, och I trodden honom icke, men publikaner och skökor trodde honom.
Och fastän I sågen detta, ångraden I eder icke heller efteråt, så att I trodden honom.
Hören nu en annan liknelse: En husbonde planterade en vingård, och han satte stängsel omkring den och högg ut ett presskar därinne och byggde ett vakttorn; därefter lejde han ut den åt vingårdsmän och for utrikes.
När sedan frukttiden nalkades, sände han sina tjänare till vingårdsmännen för att uppbära frukten åt honom.
Men vingårdsmännen togo fatt på hans tjänare, och en misshandlade de, en annan dräpte de, en tredje stenade de.
Åter sände han åstad andra tjänare, flera än de förra, men de gjorde med dem sammalunda.
Slutligen sände han till dem sin son, ty han tänkte: 'De skola väl hava försyn för min son.'
Men när vingårdsmännen fingo se hans son, sade de till varandra: 'Denne är arvingen; kom, låt oss dräpa honom, så få vi hans arv.'
Och de togo fatt på honom och förde honom ut ur vingården och dräpte honom.
När nu vingårdens herre kommer, vad skall han då göra med de vingårdsmännen?»
De svarade honom: »Eftersom de hava illa gjort, skall han illa förgöra dem, och vingården skall han lämna åt andra vingårdsmän, som giva honom frukten, när tiden därtill är inne.»
Jesus sade till dem: »Ja, haven I aldrig läst i skrifterna: 'Den sten som byggningsmännen förkastade. den har blivit en hörnsten; av Herren har den blivit detta, och underbar är den i våra ögon'?
Därför säger jag eder att Guds rike skall tagas ifrån eder, och givas åt ett folk som bär dess frukt.»
239400
Då nu översteprästerna och fariséerna hörde hans liknelser, förstodo de att det var om dem som han talade.
Och de hade gärna velat gripa honom, men de fruktade för folket, eftersom man höll honom för en profet.
Och Jesus begynte åter tala till dem i liknelser och sade:
»Med himmelriket är det, såsom när en konung gjorde bröllop åt sin son.
Han sände ut sina tjänare för att kalla till bröllopet dem som voro bjudna; men de ville icke komma.
Åter sände han ut andra tjänare och befallde dem att säga till dem som voro bjudna: 'Jag har nu tillrett min måltid, mina oxar och min gödboskap äro slaktade, och allt är redo; kommen till bröllopet.'
Men de aktade icke därpå, utan gingo bort, den ene till sitt jordagods, den andre till sin köpenskap.
Och de övriga grepo hans tjänare och misshandlade och dräpte dem.
Då blev konungen vred och sände ut sitt krigsfolk och förgjorde dråparna och brände upp deras stad.
Därefter sade han till sina tjänare: 'Bröllopet är tillrett, men de som voro bjudna voro icke värdiga.
Gån därför ut till vägskälen och bjuden till bröllopet alla som I träffen på.'
Och tjänarna gingo ut på vägarna och samlade tillhopa alla som de träffade på, både onda och goda, och bröllopssalen blev full av bordsgäster.
Men när konungen nu kom in för att se på gästerna, fick han där se en man som icke var klädd i bröllopskläder.
Då sade han till honom: 'Min vän, huru har du kommit hitin, då du icke bär bröllopskläder?'
Och han kunde intet svara.
Då sade konungen till tjänarna: 'Gripen honom vid händer och fötter, och kasten honom ut i mörkret härutanför.'
Där skall vara gråt och tandagnisslan.
Ty många äro kallade, men få utvalda.»
Därefter gingo fariséerna bort och fattade det beslutet att de skulle söka snärja honom genom något hans ord.
Och de sände till honom sina lärjungar, tillika med herodianerna, och läto dem säga: »Mästare, vi veta att du är sannfärdig och lär om Guds väg vad sant är, utan att fråga efter någon; ty du ser icke till personen.
Så säg oss då: Vad synes dig?
Är det lovligt att giva kejsaren skatt, eller är det icke lovligt?»
Men Jesus märkte deras ondska och sade: »Varför söken I att snärja mig, I skrymtare?
Låten mig se skattepenningen.»
Då lämnade de fram till honom en penning.
Därefter frågade han dem: »Vems bild och överskrift är detta?»
De svarade: »Kejsarens.»
Då sade han till dem: »Så given då kejsaren vad kejsaren tillhör, och Gud vad Gud tillhör.»
När de hörde detta, förundrade de sig.
Och de lämnade honom och gingo sin väg.
Samma dag trädde några sadducéer fram till honom och ville påstå att det icke gives någon uppståndelse; de frågade honom
och sade: »Mästare, Moses har sagt: 'Om någon dör barnlös, så skall hans broder i hans ställe äkta hans hustru och skaffa avkomma åt sin broder.'
Nu voro hos oss sju bröder.
Den förste tog sig hustru och dog, och eftersom han icke hade någon avkomma, lämnade han sin hustru efter sig åt sin broder.
Sammalunda ock den andre och den tredje, allt intill den sjunde.
Sist av alla dog hustrun.
Vilken av de sju skall då vid uppståndelsen få henne till hustru?
De hade ju alla äktat henne.»
Jesus svarade och sade till dem: »I faren vilse, ty I förstån icke skrifterna, ej heller Guds kraft.
Vid uppståndelsen taga män sig icke hustrur, ej heller givas hustrur åt män, utan de äro då såsom änglarna i himmelen.
Men vad nu angår de dödas uppståndelse, haven I icke läst vad eder är sagt av Gud:
'Jag är Abrahams Gud och Isaks Gud och Jakobs Gud'?
Han är en Gud icke för döda, utan för levande.»
När folket hörde detta, häpnade de över hans undervisning.
Men när fariséerna fingo höra att han hade stoppat munnen till på sadducéerna, samlade de sig tillhopa;
och en av dem, som var lagklok, ville snärja honom och frågade:
»Mästare, vilket är det yppersta budet i lagen?»
Då svarade han honom: »'Du skall älska HERREN, din Gud, av allt ditt hjärta och av all din själ och av allt ditt förstånd.'
Detta är det yppersta och förnämsta budet.
Därnäst kommer ett som är detta likt: 'Du skall älska din nästa såsom dig själv.'
På dessa två bud hänger hela lagen och profeterna.»
Men då nu fariséerna voro församlade, frågade Jesus dem
och sade: »Vad synes eder om Messias, vems son är han?»
De svarade honom: »Davids.»
Då sade han till dem: »Huru kan då David, genom andeingivelse, kalla honom 'herre'?
Han säger ju:
'Herren sade till min herre: Sätt dig på min högra sida, till dess jag har lagt dina fiender under dina fötter.'
Om nu David kallar honom 'herre', huru kan han då vara hans son?»
Och ingen förmådde svara honom ett ord.
Ej heller dristade sig någon från den dagen att vidare ställa någon fråga till honom.
Därefter talade Jesus till folket och till sina lärjungar
och sade: »På Moses' stol hava de skriftlärde och fariséerna satt sig.
Därför, allt vad de säga eder, det skolen I göra och hålla, men efter deras gärningar skolen I icke göra; ty de säga, men göra icke.
De binda ihop tunga bördor och lägga dem på människornas skuldror, men själva vilja de icke röra ett finger för att flytta dem.
Och alla sina gärningar göra de för att bliva sedda av människorna.
De göra sina böneremsor breda och hörntofsarna på sina mantlar stora.
De vilja gärna hava de främsta platserna vid gästabuden och sitta främst i synagogorna
och vilja gärna bliva hälsade på torgen och av människorna kallas 'rabbi'.
Men I skolen icke låta kalla eder 'rabbi', ty en är eder Mästare, och I ären alla bröder.
Ej heller skolen I kalla någon på jorden eder 'fader', ty en är eder Fader, han som är i himmelen.
Ej heller skolen I låta kalla eder 'läromästare', ty en är eder läromästare, Kristus.
Den som är störst bland eder, han vare de andras tjänare.
Men den som upphöjer sig, han skall bliva förödmjukad, och den som ödmjukar sig, han skall bliva upphöjd.
Ve eder, I skriftlärde och fariséer, I skrymtare, som tillsluten himmelriket för människorna!
Själva kommen I icke ditin, och dem som vilja komma dit tillstädjen I icke att komma in.
240020
Ve eder, I skriftlärde och fariséer, I skrymtare, som faren omkring över vatten och land för att göra en proselyt, och när någon har blivit det, gören I honom till ett Gehennas barn, dubbelt värre än I själva ären!
Ve eder, I blinde ledare, som sägen: 'Om någon svär vid templet, så betyder det intet; men om någon svär vid guldet i templet, då är han bunden av sin ed'!
I dåraktige och blinde, vilket är då förmer, guldet eller templet, som har helgat guldet?
Så ock: 'Om någon svär vid altaret, så betyder det intet; men om någon svär vid offergåvan som ligger därpå, då är han bunden av sin ed.'
I blinde, vilket är då förmer, offergåvan eller altaret, som helgar offergåvan?
Den som svär vid altaret, han svär alltså både vid detta och vid allt som ligger därpå.
Och den som svär vid templet, han svär både vid detta och vid honom som bor däri.
Och den som svär vid himmelen, han svär både vid Guds tron och vid honom som sitter därpå.
Ve eder, I skriftlärde och fariséer.
I skrymtare, som given tionde av mynta och dill och kummin, men underlåten det som är viktigast i lagen, nämligen rätten och barmhärtigheten och troheten!
Det ena borden I göra, men icke underlåta det andra.
I blinde ledare, som silen bort myggan och sväljen kamelen!
Ve eder, I skriftlärde och fariséer, I skrymtare, som gören det yttre av bägaren och fatet rent, medan de inuti äro fulla av vad I haven förvärvat genom rofferi och omättlig ondska!
Du blinde farisé, gör först insidan av bägaren ren, för att sedan också dess utsida må bliva ren.
Ve eder, I skriftlärde och fariséer, I skrymtare, som ären lika vitmenade gravar, vilka väl utanpå synas prydliga, men inuti äro fulla av de dödas ben och allt slags orenlighet!
Så synens ock I utvärtes för människorna rättfärdiga, men invärtes ären I fulla av skrymteri och orättfärdighet.
Ve eder, I skriftlärde och fariséer, I skrymtare, som byggen upp profeternas gravar och pryden de rättfärdigas grifter
och sägen: 'Om vi hade levat på våra fäders tid, så skulle vi icke hava varit delaktiga med dem i profeternas blod'!
Så vittnen I då om eder själva, att I ären barn av dem som dräpte profeterna.
Nåväl, uppfyllen då I edra fäders mått.
I ormar, I huggormars avföda, huru skullen I kunna söka undgå att dömas till Gehenna?
Se, därför sänder jag till eder profeter och vise och skriftlärde.
Somliga av dem skolen I dräpa och korsfästa, och somliga av dem skolen I gissla i edra synagogor och förfölja ifrån den ena staden till den andra.
Och så skall över eder komma allt rättfärdigt blod som är utgjutet på jorden, ända ifrån den rättfärdige Abels blod intill Sakarias', Barakias' sons blod, hans som I dräpten mellan templet och altaret.
Sannerligen säger jag eder: Allt detta skall komma över detta släkte.
Jerusalem, Jerusalem, du som dräper profeterna och stenar dem som äro sända till dig!
Huru ofta har jag icke velat församla dina barn, likasom hönan församlar sina kycklingar under sina vingar!
Men I haven icke velat.
Se, edert hus skall komma att stå övergivet och öde.