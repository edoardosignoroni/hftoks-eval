Låt ditt ansikte lysa över din tjänare, och lär mig dina stadgar.
Vattenbäckar rinna ned från mina ögon, därför att man icke håller din lag.
HERRE, du är rättfärdig, och dina domar äro rättvisa.
Du har påbjudit dina vittnesbörd i rättfärdighet och i stor trofasthet.
Jag förtäres av nitälskan, därför att mina ovänner förgäta dina ord.
Ditt tal är väl luttrat, och din tjänare har det kärt.
Jag är ringa och föraktad, men jag förgäter icke dina befallningar.
Din rättfärdighet är en evig rättfärdighet, och din lag är sanning.
Nöd och trångmål hava träffat mig, men dina bud äro min lust.
Dina vittnesbörd äro rättfärdiga evinnerligen; giv mig förstånd, så att jag får leva.
Jag ropar av allt hjärta, svara mig, HERRE; jag vill taga dina stadgar i akt.
Jag ropar till dig, fräls mig, så vill jag hålla dina vittnesbörd.
Jag kommer tidigt i morgongryningen och ropar; jag hoppas på dina ord.
Mina ögon hasta före nattens väkter till att begrunda ditt tal.
Hör min röst efter din nåd; HERRE, behåll mig vid liv efter dina rätter.
Nära äro de som jaga efter skändlighet, de som äro långt ifrån din lag.
Nära är ock du, HERRE, och alla dina bud äro sanning.
Längesedan vet jag genom dina vittnesbörd att du har stadgat dem för evig tid.
Se till mitt lidande och rädda mig, ty jag förgäter icke din lag.
Utför min sak och förlossa mig; behåll mig vid liv efter ditt tal.
Frälsning är långt borta från de ogudaktiga, ty de fråga icke efter dina stadgar.
HERRE, din barmhärtighet är stor; behåll mig vid liv efter dina rätter.
Mina förföljare och ovänner äro många, men jag viker icke ifrån dina vittnesbörd.
När jag ser de trolösa, känner jag leda vid dem, därför att de icke hålla sig vid ditt tal.
Se därtill att jag har dina befallningar kära; HERRE, behåll mig vid liv efter din nåd.
Summan av ditt ord är sanning, och alla din rättfärdighets rätter vara evinnerligen.
Furstar förfölja mig utan sak, men mitt hjärta fruktar för dina ord.
Jag fröjdar mig över ditt tal såsom den som vinner stort byte.
Jag hatar lögnen, den skall vara mig en styggelse; men din lag har jag kär.
Jag lovar dig sju gånger om dagen för din rättfärdighets rätter.
Stor frid äga de som hava din lag kär, och intet finnes, som bringar dem på fall.
Jag väntar efter din frälsning, HERRE, och jag gör efter dina bud.
Min själ håller dina vittnesbörd, och jag har dem storligen kära.
Jag håller dina befallningar och vittnesbörd, ty du känner alla mina vägar.
HERRE, mitt rop komme inför ditt ansikte; giv mig förstånd efter ditt ord.
Min bön komme inför ditt ansikte; rädda mig efter ditt tal.
Mina läppar må flöda över av lov, ty du lär mig dina stadgar.
Min tunga sjunge om ditt ord, ty alla dina bud äro rättfärdiga.
Din hand vare mig till hjälp, ty jag har utvalt dina befallningar.
Jag längtar efter din frälsning, HERRE, och din lag är min lust.
Låt min själ leva, så skall hon lova dig; och låt dina rätter hjälpa mig.
Om jag far vilse, så uppsök din tjänare såsom ett förlorat får, ty jag förgäter icke dina bud.
En vallfartssång.
Jag ropar till HERREN i min nöd, och han svarar mig.
HERRE, rädda min själ från lögnaktiga läppar, från en falsk tunga.
Varmed bliver du lönad, både nu och allt framgent, du falska tunga?
Jo, med en våldsverkares skarpa pilar och med glödande ginstkol.
Ve mig, att jag måste dväljas i Meseks land och bo ibland Kedars hyddor!
Länge nog har min själ måst bo ibland dem som hata friden.
Jag själv håller frid, men säger jag blott ett ord, äro de redo till strid.
En vallfartssång.
Jag lyfter mina ögon upp till bergen: varifrån skall min hjälp komma?
Min hjälp kommer från HERREN, som har gjort himmel och jord.
Icke skall han låta din fot vackla, icke slumrar han som bevarar dig!
Nej, han som bevarar Israel, han slumrar icke, han sover icke.
HERREN är den som bevarar dig, HERREN är ditt skygd på din högra sida.
Solen skall icke skada dig om dagen, ej heller månen om natten.
HERREN skall bevara dig för allt ont, han skall bevara din själ.
HERREN skall bevara din utgång och din ingång, från nu och till evig tid.
En vallfartssång; av David.
Jag gladdes, när man sade till mig: »Vi skola gå till HERRENS hus.»
Våra fötter fingo träda in i dina portar, Jerusalem,
Jerusalem, du nyuppbyggda stad, där hus sluter sig väl till hus,
dit stammarna draga upp, HERRENS stammar, efter lagen för Israel, till att prisa HERRENS namn.
Ty där äro ställda domarstolar, stolar för Davids hus.
Önsken Jerusalem frid; ja, dem gånge väl, som älska dig.
Frid vare inom dina murar, välgång i dina palats!
För mina bröders och vänners skull vill jag tillsäga dig frid.
För HERRENS, vår Guds, hus' skull vill jag söka din välfärd.
En vallfartssång.
Jag lyfter mina ögon upp till dig, du som bor i himmelen.
Ja, såsom tjänares ögon skåda på deras herres hand, såsom en tjänarinnas ögon på hennes frus hand, så skåda våra ögon upp till HERREN, vår Gud, till dess han varder oss nådig.
Var oss nådig, HERRE, var oss nådig, ty vi äro rikligen mättade med förakt.
Rikligen mättad är vår själ med de säkras bespottelse, med de högmodigas förakt.
En vallfartssång; av David.
Om HERREN icke hade varit med oss -- så säge Israel --
om HERREN icke hade varit med oss, när människorna reste sig upp emot oss,
då hade de uppslukat oss levande, när deras vrede upptändes mot oss;
då hade vattnen fördränkt oss, strömmen gått över vår själ;
ja, då hade de gått över vår själ, de svallande vattnen.
Lovad vare HERREN för att han ej gav oss till rov åt deras tänder!
Vår själ kom undan såsom en fågel ur fågelfängarnas snara; snaran gick sönder, och vi kommo undan.
Vår hjälp är i HERRENS namn, hans som har gjort himmel och jord.
En vallfartssång.
De som förtrösta på HERREN, de likna Sions berg, som icke vacklar, utan förbliver evinnerligen.
Jerusalem omhägnas av berg, och HERREN omhägnar sitt folk, ifrån nu och till evig tid.
Ty ogudaktighetens spira skall icke förbliva över de rättfärdigas arvslott, på det att de rättfärdiga ej må uträcka sina händer till orättfärdighet.
Gör gott, o HERRE, mot de goda och mot dem som hava redliga hjärtan.
Men dem som vika av på vrånga vägar, dem rycke HERREN bort tillika med ogärningsmännen.
Frid vare över Israel!
En vallfartssång.
När HERREN åter upprättade Sion, då voro vi såsom drömmande.
Då blev vår mun uppfylld med löje och vår tunga med jubel; då sade man bland hedningarna: »HERREN har gjort stora ting med dem.»
Ja, HERREN hade gjort stora ting med oss; däröver voro vi glada.
HERRE, upprätta oss igen, såsom du återför bäckarna i Sydlandet.
De som så med tårar skola skörda med jubel.
De gå åstad gråtande och bära sitt utsäde; de komma åter med jubel och bära sina kärvar.
En vallfartssång; av Salomo.
Om HERREN icke bygger huset, så arbeta de fåfängt, som bygga därpå.
Om HERREN icke bevarar staden, så vakar väktaren fåfängt.
Det är fåfängt att I bittida stån upp och sent gån till vila, och äten eder bröd med vedermöda; detsamma giver han åt sina vänner, medan de sova.
Se, barn äro en HERRENS gåva, livsfrukt en lön.
Likasom pilar i en hjältes hand, så äro söner som man får vid unga år.
Säll är den man som har sitt koger fyllt av sådana.
De komma icke på skam, när de mot fiender föra sin talan i porten.
En vallfartssång.
Säll är envar som fruktar HERREN och vandrar på hans vägar.
Ja, av dina händers arbete får du njuta frukten; säll är du, och väl dig!
Lik ett fruktsamt vinträd varder din hustru, därinne i ditt hus, lika olivtelningar dina barn, omkring ditt bord.
Ty se, så varder den man välsignad, som fruktar HERREN.
HERREN välsigne dig från Sion; må du få se Jerusalems välgång i alla dina livsdagar,
och må du få se barn av dina barn.
Frid över Israel!
En vallfartssång.
Mycken nöd hava de vållat mig allt ifrån min ungdom -- så säge Israel --
mycken nöd hava de vållat mig allt ifrån min ungdom, dock blevo de mig ej övermäktiga.
På min rygg hava plöjare plöjt och dragit upp långa fåror.
Men HERREN är rättfärdig och har huggit av de ogudaktigas band.
De skola komma på skam och vika tillbaka, så många som hata Sion.
De skola bliva lika gräs på taken, som vissnar, förrän det har vuxit upp;
ingen skördeman fyller därmed sin hand, ingen kärvbindare sin famn,
och de som gå där fram kunna icke säga: »HERRENS välsignelse vare över eder!
Vi välsigna eder i HERRENS namn.»
En vallfartssång.
Ur djupen ropar jag till dig, HERRE.
Herre, hör min röst, låt dina öron akta på mina böners ljud.
Om du, HERRE, vill tillräkna missgärningar, Herre, vem kan då bestå?
Dock, hos dig är ju förlåtelse, på det att man må frukta dig.
Jag väntar efter HERREN, min själ väntar, och jag hoppas på hans ord.
Min själ väntar efter Herren mer än väktarna efter morgonen, ja, mer än väktarna efter morgonen.
Hoppas på HERREN, Israel; ty hos HERREN är nåd, och mycken förlossning är hos honom.
Och han skall förlossa Israel från alla dess missgärningar.
En vallfartssång; av David.
HERRE, mitt hjärta står icke efter vad högt är, och mina ögon se ej efter vad upphöjt är, och jag umgås icke med stora ting, med ting som äro mig för svåra.
Nej, jag har lugnat och stillat min själ; såsom ett avvant barn i sin moders famn, ja, såsom ett avvant barn, så är min själ i mig.
Hoppas på HERREN, Israel, från nu och till evig tid.
En vallfartssång.
Tänk, HERRE, David till godo, på allt vad han fick lida,
han som svor HERREN en ed och gjorde ett löfte åt den Starke i Jakob;
»Jag skall icke gå in i den hydda där jag bor, ej heller bestiga mitt viloläger,
jag skall icke unna mina ögon sömn eller mina ögonlock slummer,
förrän jag har funnit en plats åt HERREN, en boning åt den Starke i Jakob.»
Ja, vi hörde därom i Efrata, vi förnummo det i skogsbygden.
Låtom oss gå in i hans boning, tillbedja vid hans fotapall.
Stå upp, HERRE, och kom till din vilostad, du och din makts ark.
Dina präster vare klädda i rättfärdighet, och dina fromma juble.
För din tjänare Davids skull må du icke visa tillbaka din smorde.
HERREN har svurit David en osviklig ed, som han icke skall rygga: »Av ditt livs frukt skall jag sätta konungar på din tron.
Om dina barn hålla mitt förbund och hålla mitt vittnesbörd, som jag skall lära dem, så skola ock deras barn till evig tid få sitta på din tron.
Ty HERREN har utvalt Sion, där vill han hava sin boning.
Detta är min vilostad till evig tid; här skall jag bo, ty till detta ställe har jag lust.
Dess förråd skall jag rikligen välsigna, åt dess fattiga skall jag giva bröd till fyllest.
Dess präster skall jag kläda i frälsning, och dess fromma skola jubla högt.
Där skall jag låta ett horn skjuta upp åt David; där har jag rett till en lampa åt min smorde.
Hans fiender skall jag kläda i skam, men på honom skall hans krona glänsa.»
En vallfartssång; av David.
Se huru gott och ljuvligt det är att bröder bo endräktigt tillsammans.
Det är likt den dyrbara oljan på huvudet, som flyter ned i skägget, ned i Arons skägg, som flyter ned över linningen på hans kläder.
Det är likt Hermons dagg, som faller ned på Sions-bergen.
Ty där beskär HERREN välsignelse, liv till evig tid.
En vallfartssång.
Upp, välsignen HERREN, alla I HERRENS tjänare, I som stån om natten i HERRENS hus.
Lyften edra händer upp mot helgedomen och välsignen HERREN.
HERREN välsigne dig från Sion, han som har gjort himmel och jord.
Halleluja!
Loven HERRENS namn, loven det, i HERRENS tjänare,
I som stån i HERRENS hus, i gårdarna till vår Guds hus.
Loven HERREN, ty HERREN är god, lovsjungen hans namn, ty det är ljuvligt.
Se, HERREN har utvalt Jakob åt sig, Israel till sin egendom.
Ty jag vet att HERREN är stor, att vår Herre är förmer än alla gudar.
HERREN kan göra allt vad han vill, i himmelen och på jorden, i haven och i alla djup;
han som låter regnskyar stiga upp från jordens ända, han som låter ljungeldar komma med regn och för vinden ut ur dess förvaringsrum;
han som slog de förstfödda i Egypten, både människor och boskap;
han som sände tecken och under över dig, Egypten, över Farao och alla hans tjänare;
han som slog stora folk och dräpte mäktiga konungar:
Sihon, amoréernas konung, och Og, konungen i Basan, med alla Kanaans riken,
och gav deras land till arvedel, till arvedel åt sitt folk Israel.
HERRE, ditt namn varar evinnerligen, HERRE, din åminnelse från släkte till släkte.
Ty HERREN skaffar rätt åt sitt folk, och över sina tjänare förbarmar han sig.
Hedningarnas avgudar äro silver och guld, verk av människohänder.
De hava mun och tala icke, de hava ögon och se icke,
de hava öron och lyssna icke till, och ingen ande är i deras mun.
De som hava gjort dem skola bliva dem lika, ja, alla som förtrösta på dem.
I av Israels hus, loven HERREN; I av Arons hus, loven HERREN;
I av Levis hus, loven HERREN; I som frukten HERREN, loven HERREN.
Lovad vare HERREN från Sion, han som bor i Jerusalem!
Halleluja!
Tacken HERREN, ty han är god, ty hans nåd varar evinnerligen.
Tacken gudarnas Gud, ty hans nåd varar evinnerligen.
Tacken herrarnas HERRE, ty hans nåd varar evinnerligen;
honom som allena gör stora under, ty hans nåd varar evinnerligen;
honom som har gjort himmelen med förstånd, ty hans nåd varar evinnerligen;
honom som har utbrett jorden över vattnen, ty hans nåd varar evinnerligen;
honom som har gjort de stora ljusen, ty hans nåd varar evinnerligen:
solen till att råda över dagen, ty hans nåd varar evinnerligen,
månen och stjärnorna till att råda över natten, ty hans nåd varar evinnerligen;
honom som slog Egypten i dess förstfödda, ty hans nåd varar evinnerligen,
och som förde Israel ut därifrån, ty hans nåd varar evinnerligen,
med stark hand och uträckt arm, ty hans nåd varar evinnerligen;
honom som delade Röda havet itu, ty hans nåd varar evinnerligen,
och lät Israel gå mitt därigenom, ty hans nåd varar evinnerligen,
och kringströdde Farao och hans här i Röda havet, ty hans nåd varar evinnerligen;
honom som förde sitt folk genom öknen, ty hans nåd varar evinnerligen,
honom som slog stora konungar, ty hans nåd varar evinnerligen,
och dräpte väldiga konungar, ty hans nåd varar evinnerligen:
Sihon, amoréernas konung, ty hans nåd varar evinnerligen,
och Og, konungen i Basan, ty hans nåd varar evinnerligen;
och som gav deras land till arvedel, ty hans nåd varar evinnerligen,
till arvedel åt sin tjänare Israel, ty hans nåd varar evinnerligen;
honom som tänkte på oss i vår förnedring, ty hans nåd varar evinnerligen,
och som ryckte oss ur våra ovänners våld, ty hans nåd varar evinnerligen;
honom som giver mat åt allt levande, ty hans nåd varar evinnerligen.
Tacken himmelens Gud, ty hans nåd varar evinnerligen.
Vid Babels floder, där sutto vi och gräto, när vi tänkte på Sion.
I pilträden som där voro hängde vi upp våra harpor.
Ty de som höllo oss fångna bådo oss där att sjunga, och våra plågare bådo oss vara glada: »Sjungen för oss en av Sions sånger.»
Huru skulle vi kunna sjunga HERRENS sång i främmande land?
Nej, om jag förgäter dig, Jerusalem, så förgäte min högra hand sin tjänst.
Min tunga låde vid min gom, om jag upphör att tänka på dig, om jag icke låter Jerusalem vara min allra högsta glädje.
Tänk, HERRE, på Jerusalems dag, och straffa Edoms barn, dem som ropade: »Riven ned, riven ned det ända till grunden.»
Dotter Babel, du ödeläggelsens stad, säll är den som får vedergälla dig allt vad du har gjort oss.
Säll är den som får gripa dina späda barn och krossa dem mot klippan.
Av David.
Jag vill tacka dig av allt mitt hjärta; inför gudarna vill jag lovsjunga dig.
Jag vill tillbedja, vänd mot ditt heliga tempel, och prisa ditt namn för din nåd och sanning, ty du har gjort ditt löftesord stort utöver allt vad ditt namn hade sagt.
När jag ropade, svarade du mig; du gav mig frimodighet, och min själ fick kraft.
HERRE, alla jordens konungar skola tacka dig, när de få höra din muns tal.
De skola sjunga om HERRENS vägar, ty HERRENS ära är stor.
Ja, HERREN är hög, men han ser till det låga, och han känner den högmodige fjärran ifrån.
Om ock min väg går genom nöd, så behåller du mig vid liv; du räcker ut din hand till värn mot mina fienders vrede, och din högra hand frälsar mig.
HERREN skall fullborda sitt verk för mig.
HERRE, din nåd varar evinnerligen; övergiv icke dina händers verk.
För sångmästaren; av David; en psalm.
HERRE, du utrannsakar mig och känner mig.
Evad jag sitter eller uppstår, vet du det; du förstår mina tankar fjärran ifrån.
Evad jag går eller ligger, utforskar du det, och med alla mina vägar är du förtrogen.
Ty förrän ett ord är på min tunga, se, så känner du, HERRE, det till fullo.
Du omsluter mig på alla sidor och håller mig i din hand.
En sådan kunskap är mig alltför underbar; den är mig för hög, jag kan icke begripa den.
Vart skall jag gå för din Ande, och vart skall jag fly för ditt ansikte?
Fore jag upp till himmelen, så är du där, och bäddade jag åt mig i dödsriket, se, så är du ock där.
Toge jag morgonrodnadens vingar, gjorde jag mig en boning ytterst i havet,
så skulle också där din hand leda mig och din högra hand fatta mig.
Och om jag sade: »Mörker må betäcka mig och ljuset bliva natt omkring mig»,
så skulle själva mörkret icke vara mörkt för dig, natten skulle lysa såsom dagen: ja, mörkret skulle vara såsom ljuset.
Ty du har skapat mina njurar, du sammanvävde mig i min moders liv.
Jag tackar dig för att jag är danad så övermåttan underbart; ja, underbara äro dina verk, min själ vet det väl.
Benen i min kropp voro icke förborgade för dig, när jag bereddes i det fördolda, när jag bildades i jordens djup.
Dina ögon sågo mig, när jag ännu knappast var formad; alla mina dagar blevo uppskrivna i din bok, de voro bestämda, förrän någon av dem hade kommit.
Huru outgrundliga äro icke för mig dina tankar, o Gud, huru stor är icke deras mångfald!
Skulle jag räkna dem, så vore de flera än sanden; när jag uppvaknade, vore jag ännu hos dig.
Gud, o att du ville dräpa de ogudaktiga!
Ja, måtte de blodgiriga vika bort ifrån mig,
de som tala om dig med ränker i sinnet, de som hava bragt dina städer i fördärv!
Skulle jag icke hata dem som hata dig, HERRE?
Skulle jag icke känna leda vid dem som stå dig emot?
Jag hatar dem med starkaste hat; ja, mina fiender hava de blivit.
Utrannsaka mig, Gud, och känn mitt hjärta; pröva mig och känn mina tankar,
och se till, om jag är stadd på en olycksväg, och led mig på den eviga vägen.
För sångmästaren; en psalm av David.
Rädda mig, HERRE, från onda människor, bevara mig från våldets män,
för dem som uttänka ont i sina hjärtan och dagligen rota sig samman till strid.
De vässa sina tungor likasom ormar, huggormsgift är inom deras läppar.
Sela.
Bevara mig, HERRE, för de ogudaktigas händer, beskydda mig för våldets män, som uttänka planer för att bringa mig på fall.
Stolta människor lägga ut för mig snaror och garn; de breda ut nät invid vägens rand, giller sätta de för mig.
Sela.
Jag säger till HERREN: »Du är min Gud.»
Lyssna, o HERRE, till mina böners ljud.
HERRE, Herre, du min starka hjälp, du beskärmar mitt huvud, på stridens dag.
Tillstäd icke, HERRE; vad de ogudaktiga begära; låt deras anslag ej lyckas, de skulle eljest förhäva sig.
Sela.
Över de mäns huvuden, som omringa mig, må den olycka komma, som deras läppar bereda.
Eldsglöd må regna över dem; må de kastas i eld, i djup som de ej komma upp ur.
En förtalets man skall ej bestå i landet; en ond våldsman skall jagas, med slag på slag.
Jag vet att HERREN skall utföra den betrycktes sak och skaffa de fattiga rätt.
Ja, de rättfärdiga skola prisa ditt namn och de redliga bo inför ditt ansikte.
En psalm av David.
HERRE, jag ropar till dig, skynda till mig; lyssna till min röst, då jag nu ropar till dig.
Min bön gälle inför dig såsom ett rökoffer, mina händers upplyftande såsom ett aftonoffer.
Sätt, o HERRE, en vakt för min mun, bevaka mina läppars dörr.
Låt icke mitt hjärta vika av till något ont, till att öva ogudaktighetens gärningar tillsammans med män som göra vad orätt är; av deras läckerheter vill jag icke äta.
Må den rättfärdige slå mig i kärlek och straffa mig; det är såsom olja på huvudet, och mitt huvud skall icke försmå det.
Ty ännu en tid, så skall min bön uppfyllas, genom att det går dem illa;
deras ledare skola störtas ned utför klippan, och man skall då höra att mina ord äro ljuvliga.
Såsom när man har plöjt och ristat upp jorden, så ligga våra ben kringströdda vid dödsrikets rand.
Ja, till dig, HERRE, Herre, se mina ögon; till dig tager jag min tillflykt, förkasta icke min själ.
Bevara mig för de snaror som de lägga ut på min väg och för ogärningsmännens giller.
De ogudaktiga falle i sina egna garn, medan jag går oskadd förbi.
En sång av David; en bön, när han var i grottan.
Jag höjer min röst och ropar till HERREN, jag höjer min röst och beder till HERREN.
Jag utgjuter inför honom mitt bekymmer, min nöd kungör jag för honom.
När min ande försmäktar i mig, är du den som känner min stig.
På den väg där jag skall gå hava de lagt ut snaror för mig.
Skåda på min högra sida och se: där finnes ingen som kännes vid mig.
Ingen tillflykt återstår för mig, ingen finnes, som frågar efter min själ.
Jag ropar till dig, o HERRE, jag säger: »Du är min tillflykt, min del i de levandes land.»
Akta på mitt rop, ty jag är i stort elände; rädda mig från mina förföljare, ty de äro mig övermäktiga.
För min själ ut ur fängelset, så att jag får prisa ditt namn.
Omkring mig skola de rättfärdiga församlas, när du gör väl mot mig.
En psalm av David.
HERRE, hör min bön, lyssna till min åkallan, svara mig i din rättfärdighet, för din trofasthets skull.
Och gå icke till doms med din tjänare, ty inför dig är ingen levande rättfärdig.
Se, fienden förföljer min själ, han trampar mitt liv till jorden; han lägger mig i mörker såsom de längesedan döda.
Och min ande försmäktar i mig, mitt hjärta är stelnat i mitt bröst.
Jag tänker på forna dagar, jag begrundar alla dina gärningar, dina händers verk eftersinnar jag.
Jag uträcker mina händer till dig; såsom ett törstigt land längtar min själ efter dig.
Sela.
HERRE, skynda att svara mig, ty min ande förgås; dölj icke ditt ansikte för mig, må jag ej varda lik dem som hava farit ned i graven.
Låt mig bittida förnimma din nåd, ty jag förtröstar på dig.
Kungör mig den väg som jag bör vandra, ty till dig upplyfter jag min själ.
Rädda mig från mina fiender, HERRE; hos dig söker jag skygd.
Lär mig att göra din vilja, ty du är min Gud; din gode Ande lede mig på jämn mark.
HERRE, behåll mig vid liv för ditt namns skull; tag min själ ut ur nöden för din rättfärdighets skull.
Utrota mina fiender för din nåds skull, och förgör alla dem som tränga min själ; ty jag är din tjänare.
Av David.
Lovad vare HERREN, min klippa, han som lärde mina armar att kriga, mina händer att strida;
min nåds Gud och min borg, mitt värn och min räddare, min sköld och min tillflykt, han som lägger mitt folk under mig.
HERRE, vad är en människa, att du vill veta av henne, en människoson, att du tänker på honom?
En människa är lik en fläkt, hennes dagar såsom en försvinnande skugga.
HERRE, sänk din himmel och far ned, rör vid bergen, så att de ryka.
Låt ljungeldar ljunga och skingra dem, skjut dina pilar och förvirra dem.
Räck ut dina händer från höjden, fräls mig och rädda mig ur de stora vattnen, ur främlingarnas hand,
vilkas mun talar lögn och vilkas högra hand är en falskhetens hand.
Gud, en ny sång vill jag sjunga till din ära, till tiosträngad psaltare vill jag lovsjunga dig,
dig som giver seger åt konungarna, dig som frälste din tjänare David från det onda svärdet.
Fräls mig och rädda mig ur främlingarnas hand, vilkas mun talar lögn, och vilkas högra hand är en falskhetens hand.
När våra söner stå i sin ungdom såsom högväxta plantor, våra döttrar lika hörnstoder, huggna såsom för palatser;
när våra visthus äro fulla och skänka förråd på förråd; när våra får öka sig tusenfalt, ja, tiotusenfalt på våra utmarker;
när våra oxar gå rikt lastade; när ingen rämna har brutits i muren och ingen nödgas draga ut såsom fånge, när intet klagorop höres på våra gator --
saligt är det folk som det så går; ja, saligt är det folk vars Gud HERREN är.
En lovsång av David.
Jag vill upphöja dig, min Gud, du konung, och lova ditt namn alltid och evinnerligen.
Jag vill dagligen lova dig och prisa ditt namn alltid och evinnerligen.
Stor är HERREN och högtlovad, ja, hans storhet är outrannsaklig.
Det ena släktet prisar för det andra dina verk, de förkunna dina väldiga gärningar.
Ditt majestäts härlighet och ära vill jag begrunda och dina underfulla verk.
Man skall tala om dina fruktansvärda gärningars makt; dina storverk skall jag förtälja.
Man skall utbreda ryktet om din stora godhet och jubla över din rättfärdighet.
Nådig och barmhärtig är HERREN, långmodig och stor i mildhet.
HERREN är god mot alla och förbarmar sig över alla sina verk.
Alla dina verk, HERRE, skola tacka dig, och dina fromma skola lova dig.
De skola tala om ditt rikes ära, och din makt skola de förkunna.
Så skola de kungöra för människors barn dina väldiga gärningar och ditt rikes ära och härlighet.
Ditt rike är ett rike för alla evigheter, och ditt herradöme varar från släkte till släkte.
HERREN uppehåller alla dem som äro på väg att falla, och han upprättar alla nedböjda.
Allas ögon vänta efter dig, och du giver dem deras mat i rätt tid.
Du upplåter din hand och mättar allt levande med nåd.
HERREN är rättfärdig i alla sina vägar och nådig i alla sina verk.
HERREN är nära alla dem som åkalla honom, alla dem som åkalla honom uppriktigt.
Han gör vad de gudfruktiga begära och hör deras rop och frälsar dem.
HERREN bevarar alla dem som älska honom, men alla ogudaktiga skall han förgöra.
Min mun skall uttala HERREN lov, och allt kött skall prisa hans heliga namn alltid och evinnerligen.
Halleluja!
Lova HERREN, min själ.
Jag vill lova HERREN, så länge jag lever, jag vill lovsjunga min Gud, så länge jag är till.
Förliten eder icke på furstar, icke på en människoson, han kan icke hjälpa.
Hans ande måste sin väg, han vänder tillbaka till den jord varav han är kommen; då varda hans anslag om intet.
Säll är den vilkens hjälp är Jakobs Gud, den vilkens hopp står till HERREN, hans Gud,
till honom som har gjort himmelen och jorden och havet och allt vad i dem är, till honom som håller tro evinnerligen,
som skaffar rätt åt de förtryckta, som giver bröd åt de hungrande.
HERREN löser de fångna,
HERREN öppnar de blindas ögon, HERREN upprättar de nedböjda, HERREN älskar de rättfärdiga,
HERREN bevarar främlingar, faderlösa och änkor uppehåller han; men de ogudaktigas väg vänder han i villa.
HERREN är konung evinnerligen, din Gud, Sion, från släkte till släkte.
Halleluja!
Halleluja!
Ja, det är gott att lovsjunga vår Gud, ja, det är ljuvligt; lovsång höves oss.
HERREN är den som bygger upp Jerusalem, Israels fördrivna samlar han tillhopa.
Han helar dem som hava förkrossade hjärtan, och deras sår förbinder han.
Han bestämmer stjärnornas mängd, han nämner dem alla vid namn.
Vår Herre är stor och väldig i kraft, hans förstånd har ingen gräns.
HERREN uppehåller de ödmjuka, men de ogudaktiga slår han till jorden.
Höjen sång till HERREN med tacksägelse, lovsjungen vår Gud till harpa,
honom som betäcker himmelen med moln, honom som bereder regn åt jorden, honom som låter gräs skjuta upp på bergen,
honom som giver föda åt djuren, åt korpens ungar som ropa.
Han har icke sin lust i hästens styrka, hans behag står ej till mannens snabbhet.
HERRENS behag står till dem som frukta honom, till dem som hoppas på hans nåd.
Jerusalem, prisa HERREN; Sion, lova din Gud.
Ty han har gjort bommarna för dina portar fasta; han har välsignat dina barn i dig.
Han skaffar dina gränser frid, han mättar dig med bästa vete.
Han låter sitt tal gå ut till jorden, hans ord löper åstad med hast.
Han låter snö falla såsom ull, rimfrost strör han ut såsom aska.
Han kastar sitt hagel såsom smulor; vem kan bestå för hans frost?
Åter sänder han sitt ord, då smälter det frusna; sin vind låter han blåsa, då strömmar vatten.
Han har förkunnat för Jakob sitt ord, för Israel sina stadgar och rätter.
Så har han icke gjort för något hednafolk; och hans rätter, dem känna de icke.
Halleluja!
Halleluja!
Loven HERREN från himmelen, loven honom i höjden.
Loven honom, alla hans änglar, loven honom, all hans här.
Loven honom, sol och måne, loven honom, alla lysande stjärnor.
Loven honom, I himlars himlar och I vatten ovan himmelen.
Ja, de må lova HERRENS namn, ty han bjöd, och de blevo skapade.
Och han gav dem deras plats för alltid och för evigt; han gav dem en lag, och ingen överträder den.
Loven HERREN från jorden, I havsdjur och alla djup,
eld och hagel, snö och töcken, du stormande vind, som uträttar hans befallning,
I berg och alla höjder, I fruktträd och alla cedrar,
I vilda djur och all boskap, I kräldjur och bevingade fåglar,
I jordens konungar och alla folk, I furstar och alla domare på jorden,
I ynglingar, så ock I jungfrur, I gamle med de unga.
Ja, de må lova HERRENS namn, ty hans namn allena är högt, hans majestät når över jorden och himmelen.
Och han har upphöjt ett horn åt sitt folk -- ett ämne till lovsång för alla hans fromma, för Israels barn, det folk som står honom nära.
Halleluja!
Halleluja!
Sjungen till HERRENS ära en ny sång, hans lov i de frommas församling.
Israel glädje sig över sin skapare, Sions barn fröjde sig över sin konung.
Må de lova hans namn under dans, till puka och harpa må de lovsjunga honom.
Ty HERREN har behag till sitt folk, han smyckar de ödmjuka med frälsning.
De fromma fröjde sig och give honom ära, de juble på sina läger.
Guds lov skall vara i deras mun och ett tveeggat svärd i deras hand,
för att utkräva hämnd på hedningarna och hemsöka folken med tuktan,
för att binda deras konungar med kedjor och deras ädlingar med järnbojor,
för att utföra på dem den dom som är skriven.
En härlighet bliver det för alla hans fromma.
Halleluja!
Halleluja!
Loven Gud i hans helgedom, loven honom i hans makts fäste.
Loven honom för hans väldiga gärningar, loven honom efter hans stora härlighet
Loven honom med basunklang, loven honom med psaltare och harpa.
Loven honom med puka och dans, loven honom med strängaspel och pipa.
Loven honom med ljudande cymbaler, loven honom med klingande cymbaler.
Allt vad anda har love HERREN.
Halleluja!
Detta är Salomos ordspråk, Davids sons, Israels konungs.
Av dem kan man lära vishet och tukt,
så ock att förstå förståndigt tal.
Av dem kan man undfå tuktan till insikt och lära rättfärdighet, rätt och redlighet.
De kunna giva åt de fåkunniga klokhet, åt den unge kunskap och eftertänksamhet.
Genom att höra på dem förökar den vise sin lärdom och förvärvar den förståndige rådklokhet.
Av dem lär man förstå ordspråk och djupsinnigt tal, de vises ord och deras gåtor.
HERRENS fruktan är begynnelsen till kunskap; vishet och tuktan föraktas av oförnuftiga.
Hör, min son, din faders tuktan, och förkasta icke din moders undervisning.
Ty sådant är en skön krans för ditt huvud och en kedja till prydnad för din hals.
Min son, om syndare locka dig, så följ icke.
Om de säga: »Kom med oss; vi vilja lägga oss på lur efter blod, sätta försåt för de oskyldiga, utan sak;
såsom dödsriket vilja vi uppsluka dem levande, friska och sunda, såsom fore de ned i graven;
allt vad dyrbart är skola vi vinna, vi skola fylla våra hus med byte;
dela du med oss vår lott, alla skola vi hava samma pung» --
då, min son, må du ej vandra samma väg som de.
Nej, håll din fot ifrån deras stig,
ty deras fötter hasta till vad ont är, och äro snara, när det gäller att utgjuta blod.
Ty väl är det fåfängt, då man vill fånga fåglar, att breda ut nätet i hela flockens åsyn.
Men dessa ligga på lur efter sitt eget blod, de sätta försåt för sina egna liv.
Så går det envar som söker orätt vinning: sin egen herre berövar den livet.
Visheten höjer sitt rop på gatan, på torgen låter hon höra sin röst.
I bullrande gathörn predikar hon; där portarna i staden öppna sig, där talar hon sina ord:
Huru länge, I fåkunnige, skolen I älska fåkunnighet?
Huru länge skola bespottarna hava sin lust i bespottelse och dårarna hata kunskap?
Vänden om och akten på min tillrättavisning; se, då skall jag låta min ande flöda för eder jag skall låta eder förnimma mina ord.
Eftersom I icke villen höra, när jag ropade, eftersom ingen aktade på, när jag räckte ut min hand,
eftersom I läten allt mitt råd fara och icke villen veta av min tillrättavisning
därför skall ock jag le vid eder ofärd och bespotta, när det kommer, som I frukten,
ja, när det I frukten kommer såsom ett oväder, när ofärden nalkas eder såsom en storm och över eder kommer nöd och ångest.
Då skall man ropa till mig, men jag skall icke svara, man skall söka mig, men icke finna mig.
Därför att de hatade kunskap och icke funno behag i HERRENS fruktan,
ej heller ville följa mitt råd, utan föraktade all min tillrättavisning,
därför skola de få äta sina gärningars frukt och varda mättade av sina egna anslag.
Ty av sin avfällighet skola de fåkunniga dräpas. och genom sin säkerhet skola dårarna förgås.
Men den som hör mig, han skall bo i trygghet och vara säker mot olyckans skräck.
Min son, om du tager emot mina ord och gömmer mina bud inom dig,
så att du låter ditt öra akta på visheten och böjer ditt hjärta till klokheten,
ja, om du ropar efter förståndet och höjer din röst till att kalla på klokheten,
Om du söker efter henne såsom efter silver och letar efter henne såsom efter en skatt,
då skall du förstå HERRENS fruktan, och Guds kunskap skall du då finna.
Ty HERREN är den som giver vishet; från hans mun kommer kunskap och förstånd.
Åt de redliga förvarar han sällhet, han är en sköld för dem som vandra i ostrafflighet,
ty han beskyddar det rättas stigar, och sina frommas väg bevarar han.
Då skall du förstå rättfärdighet och rätt och redlighet, ja, det godas alla vägar.
Ty visheten skall draga in i ditt hjärta och kunskapen kännas ljuvlig för din själ,
eftertänksamheten skall vaka över dig, klokheten skall beskydda dig.
Så skall hon rädda dig från de ondas väg, från män som tala vad vrångt är,
från dem som hava övergivit det rättas stigar. för att färdas på mörkrets vägar,
från dem som glädjas att göra om och fröjda sig åt ondskans vrånga väsen,
från dem som gå på krokiga stiga och vandra på förvända vägar.
Så skall hon rädda dig ifrån främmande kvinnor, från din nästas hustru, som talar hala ord,
från henne som har övergivit sin ungdoms vän och förgätit sin Guds förbund.
Ty en sådan sjunker med sitt hus ned i döden, och till skuggornas boning leda hennes stigar.
Ingen som har gått in till henne vänder åter Och hittar tillbaka till livets vägar.
Ja, så skall du vandra på de godas väg och hålla dig på de rättfärdigas stigar.
Ty de redliga skola förbliva boende i landet och de ostraffliga få stanna kvar däri.
Men de ogudaktiga skola utrotas ur landet och de trolösa ryckas bort därur.
Min son, förgät icke min undervisning, och låt ditt hjärta bevara mina bud.
Ty långt liv och många levnadsår och frid, mer och mer, skola de bereda dig.
Låt godhet och sanning ej vika ifrån dig; bind dem omkring din hals, skriv dem på ditt hjärtas tavla;
så skall du finna nåd och få gott förstånd, i Guds och i människors ögon.
Förtrösta på HERREN av allt ditt hjärta, och förlita dig icke på ditt förstånd.
På alla dina vägar må du akta på honom, så skall han göra dina stigar jämna.
Håll dig icke själv för vis; frukta HERREN, och fly det onda.
Det skall vara ett hälsomedel för din kropp och en vederkvickelse för benen däri.
Ära HERREN med dina ägodelar! och med förstlingen av all din gröda,
så skola dina lador fyllas med ymnighet, och av vinmust skola dina pressar flöda över.
Min son, förkasta icke HERRENS tuktan, och förargas icke, när du agas av honom.
Ty den HERREN älskar, den agar han, likasom en fader sin son, som han har kär.
Säll är den människa som har funnit visheten, den människa som undfår förstånd.
Ty bättre är att förvärva henne än att förvärva silver, och den vinning hon giver är bättre än guld.
Dyrbarare är hon än pärlor; allt vad härligt du äger går ej upp emot henne.
Långt liv bär hon i sin högra hand, i sin vänstra rikedom och ära.
Hennes vägar äro ljuvliga vägar, och alla hennes stigar äro trygga.
Ett livets träd är hon för dem som få henne fatt, och sälla må de prisa, som hålla henne kvar.
Genom vishet har HERREN lagt jordens grund, himmelen har han berett med förstånd.
Genom hans insikt bröto djupens vatten fram, och genom den låta skyarna dagg drypa ned.
Min son, låt detta icke vika ifrån dina ögon, tag klokhet och eftertänksamhet i akt;
så skola de lända din själ till liv bliva ett smycke för din hals.
Då skall du vandra din väg fram i trygghet, och din fot skall du då icke stöta.
När du lägger dig, skall intet förskräcka dig, och sedan du har lagt dig, skall du sova sött.
Du behöver då ej frukta för plötslig skräck, ej för ovädret, när det kommer över de ogudaktiga.
Ty HERREN skall då vara ditt hopp, och han skall bevara din fot för snaran.
Neka icke den behövande din hjälp, är det står i din makt att giva den.
Säg icke till din nästa: »Gå din väg och kom igen; i morgon vill jag giva dig», fastän du kunde strax.
Stämpla intet ont mot din nästa, när han menar sig bo trygg i din närhet.
Tvista icke med någon utan sak, då han icke har gjort dig något ont.
Avundas icke den orättrådige, och finn ej behag i någon av hans vägar.
Ty en styggelse för HERREN är den vrånge, men med de redliga har han sin umgängelse.
HERRENS förbannelse vilar över den ogudaktiges hus, men de rättfärdigas boning välsignar han.
Har han att skaffa med bespottare, så bespottar också han; men de ödmjuka giver han nåd.
De visa få ära till arvedel, men dårarna få uppbära skam.
Hören, I barn, en faders tuktan, och akten därpå, så att I lären förstånd.
Ty god lärdom giver jag eder; min undervisning mån I icke låta fara.
Ty själv har jag varit barn och haft en fader, varit späd och för min moder ende sonen.
Då undervisade han mig och sade till mig: Låt ditt hjärta hålla fast vid mina ord; bevara mina bud, så får du leva.
Sök förvärva vishet, sök förvärva förstånd, förgät icke min muns tal och vik icke därifrån.
Övergiv henne icke, så skall hon bevara dig; älska henne, så skall hon beskydda dig.
Vishetens begynnelse är: »Sök förvärva vishet»; ja, för allt ditt förvärv sök förvärva förstånd.
Akta henne högt, så skall hon upphöja dig; hon skall göra dig ärad, om du sluter henne i din famn.
Hon skall sätta på ditt huvud en skön krans; en ärekrona skall hon räcka åt dig.
Hör, min son, och tag emot mina ord, så skola dina levnadsår bliva många.
Om vishetens väg undervisar jag dig, jag leder dig på det rättas stigar.
När du går, skall sedan intet vara till hinder för dina steg, och när du löper, skall du icke falla;
håll blott oavlåtligt fast vid min tuktan; bevara henne, ty hon är ditt liv.
Träd icke in på de ogudaktigas stig, och skrid icke fram på de ondas väg.
Undfly den, gå ej in på den, vik av ifrån den och gå undan.
Ty de kunna icke sova, om de ej få göra vad ont är, sömnen förtages dem, om de ej få vålla någons fall.
Ja, ogudaktighet är det bröd som de äta, och våld är det vin som de dricka.
De rättfärdigas stig är lik gryningens ljus, som växer i klarhet, till dess dagen når sin höjd;
men de ogudaktigas väg är såsom tjocka mörkret: de märka icke det som skall vålla deras fall.
Min son, akta på mitt tal, böj ditt öra till mina ord.
Låt dem icke vika ifrån dina ögon, bevara dem i ditt hjärtas djup.
Ty de äro liv för envar som finner dem, och en läkedom för hela hans kropp.
Framför allt som skall bevaras må du bevara ditt hjärta, ty därifrån utgår livet.
Skaffa bort ifrån dig munnens vrånghet, och låt läpparnas falskhet vara fjärran ifrån dig.
Låt dina ögon skåda rätt framåt och dina blickar vara riktade rakt ut.
Akta på den stig där din fot går fram, och låt alla dina vägar vara rätta.
Vik ej av, vare sig till höger eller till vänster, vänd din fot bort ifrån vad ont är.
Min son, akta på min vishet, böj ditt öra till mitt förstånd,
så att du bevarar eftertänksamhet och låter dina läppar taga kunskap i akt.
Se, av honung drypa en trolös kvinnas läppar, och halare än olja är hennes mun.
Men på sistone bliver hon bitter såsom malört och skarp såsom ett tveeggat svärd.
Hennes fötter styra nedåt mot döden till dödsriket draga hennes steg.
Livets väg vill hon ej akta på; hennes stigar äro villostigar, fastän hon ej vet det.
Så hören mig nu, I barn, och viken icke ifrån min muns tal.
Låt din väg vara fjärran ifrån henne, och nalkas icke dörren till hennes hus.
Må du ej åt andra få offra din ära, ej dina år åt en som hämnas grymt;
må icke främmande få mätta sig av ditt gods och dina mödors frukt komma i en annans hus,
så att du själv på sistone måste sucka, när ditt hull och ditt kött är förtärt.
och säga: »Huru kunde jag så hata tuktan, huru kunde mitt hjärta så förakta tillrättavisning!
Varför lyssnade jag icke till mina lärares röst, och böjde icke mitt öra till dem som ville undervisa mig?
Föga fattas nu att jag har drabbats av allt vad ont är, mitt i församling och menighet.
Drick vatten ur din egen brunn det vatten som rinner ur din egen källa.
Icke vill du att dina flöden skola strömma ut på gatan, dina vattenbäckar på torgen?
Nej, dig allena må de tillhöra, och ingen främmande jämte dig.
Din brunn må vara välsignad, och av din ungdoms hustru må du hämta din glädje;
hon, den älskliga hinden, den täcka gasellen, hennes barm förnöje dig alltid, i hennes kärlek finne du ständig din lust.
Min son, icke skall du hava din lust i en främmande kvinna?
Icke skall du sluta din nästas hustru i din famn?
Se, för HERRENS ögon ligga var människas vägar blottade, och på alla hennes stigar giver han akt.
Den ogudaktige fångas av sina egna missgärningar och fastnar i sin egen synds snaror.
Han måste dö, därför att han icke lät tukta sig; ja, genom sin stora dårskap kommer han på fall.
Min son, om du har gått i borgen för din nästa och givit ditt handslag för en främmande,
om du har blivit bunden genom din muns tal, ja, fångad genom din muns tal,
då, min son, må du göra detta för att rädda dig, eftersom du har kommit i din nästas våld: gå och kasta dig ned för honom och ansätt honom,
unna dina ögon ingen sömn och dina ögonlock ingen slummer.
Sök räddning såsom en gasell ur jägarens våld, och såsom en fågel ur fågelfängarens våld.
Gå bort till myran, du late; se huru hon gör, och bliv vis.
Hon har ingen furste över sig, ingen tillsyningsman eller herre;
dock bereder hon om sommaren sin föda och samlar under skördetiden in sin mat.
Huru länge vill du ligga, du late?
När vill du stå upp ifrån din sömn?
Ja, sov ännu litet, slumra ännu litet, lägg ännu litet händerna i kors för att vila,
så skall fattigdomen komma över dig såsom en rövare och armodet såsom en väpnad man.
En fördärvlig människa, ja, en ogärningsman är den som går omkring med vrånghet i munnen,
som blinkar med ögonen, skrapar med fötterna, giver tecken med fingrarna.
Svek bär en sådan i sitt hjärta, ont bringar han alltid å bane, trätor kommer han åstad.
Därför skall ofärd plötsligt komma över honom; oförtänkt varder han krossad utan räddning.
Sex ting är det som HERREN hatar, ja, sju äro styggelser för hans själ
stolta ögon, en lögnaktig tunga, händer som utgjuta oskyldigt blod,
ett hjärta som hopsmider fördärvliga anslag, fötter som äro snara till att löpa efter vad ont är,
den som främjar lögn genom falskt vittnesbörd, och den som vållar trätor mellan bröder.
Min son, bevara din faders bud, och förkasta icke din moders undervisning.
Hav dem alltid bundna vid ditt hjärta, fäst dem omkring din hals.
När du går, må de leda dig, när du ligger, må de vaka över dig, och när du vaknar upp, må de tala till dig.
Ty budet är en lykta och undervisningen ett ljus, och tillrättavisningar till tukt äro en livets väg.
De kunna bevara dig för onda kvinnor, för din nästas hustrus hala tunga.
Hav icke begärelse i ditt hjärta till hennes skönhet, och låt henne icke fånga dig med sina blickar.
Ty för skökan måste du lämna din sista brödkaka, och den gifta kvinnan går på jakt efter ditt dyra liv.
Kan väl någon hämta eld i sitt mantelveck utan att hans kläder bliva förbrända?
Eller kan någon gå på glödande kol, utan att hans fötter varda svedda?
Så sker ock med den som går in till sin nästas hustru; ostraffad bliver ingen som kommer vid henne.
Föraktar man icke tjuven som stjäl för att mätta sitt begär, när han hungrar?
Och han måste ju, om han ertappas, betala sjufalt igen och giva allt vad han äger i sitt hus.
Så är ock den utan förstånd, som förför en annans hustru; ja, en självspilling är den som sådant gör.
Plåga och skam är vad han vinner, och hans smälek utplånas icke.
Ty svartsjuk är mannens vrede, och han skonar icke på hämndens dag;
lösepenning aktar han alls icke på, och bryr sig ej om att du bjuder stora skänker.
Min son, tag vara på mina ord, och göm mina bud inom dig.
Håll mina bud, så får du leva, och bevara min undervisning såsom din ögonsten.
Bind dem vid dina fingrar, skriv dem på ditt hjärtas tavla.
Säg till visheten: »Du är min syster», och kalla förståndet din förtrogna,
så att de bevara dig för främmande kvinnor, för din nästas hustru, som talar hala ord.
Ty ut genom fönstret i mitt hus, fram genom gallret där blickade jag;
då såg jag bland de fåkunniga, jag blev varse bland de unga en yngling utan förstånd.
Han gick fram på gatan invid hörnet där hon bodde, på vägen till hennes hus skred han fram,
skymningen, på aftonen av dagen, nattens dunkel, när mörker rådde
Se, då kom där en kvinna honom till mötes; hennes dräkt var en skökas, och hennes hjärta illfundigt.
Yster och lättsinnig var hon, hennes fötter hade ingen ro i hennes hus.
Än var hon på gatan, än var hon på torgen vid vart gathörn stod hon på lur.
Hon tog nu honom fatt och kysste honom och sade till honom med fräckhet i sin uppsyn:
»Tackoffer har jag haft att frambära; i dag har jag fått infria mina löften.
Därför gick jag ut till att möta dig jag ville söka upp dig, och nu ha jag funnit dig.
Jag har bäddat min säng med sköna täcken, med brokigt linne från Egypten.
Jag har bestänkt min bädd med myrra, med aloe och med kanel.
Kom, låt oss förnöja oss med kärlek intill morgonen, och förlusta oss med varandra i älskog.
Ty min man är nu icke hemma han har rest en lång väg bort.
Sin penningpung tog han med sig; först vid fullmånstiden kommer han hem.»
Så förleder hon honom med allahanda fagert tal; genom sina läppars halhet förför hon honom.
Han följer efter henne med hast, lik oxen som går för att slaktas, och lik fången som föres bort till straffet för sin dårskap;
ja, han följer, till dess pilen genomborrar hans lever, lik fågeln som skyndar till snaran, utan att förstå att det gäller dess liv.
Så hören mig nu, I barn, och given akt på min muns tal.
Låt icke ditt hjärta vika av till hennes vägar, och förvilla dig ej in på hennes stigar.
Ty många som ligga slagna äro fällda av henne, och stor är hopen av dem hon har dräpt.
Genom hennes hus gå dödsrikets vägar, de som föra nedåt till dödens kamrar.
Hör, visheten ropar, och förståndet höjer sin röst.
Uppe på höjderna står hon, vid vägen, där stigarna mötas.
Invid portarna, vid ingången till staden där man träder in genom dörrarna, höjer hon sitt rop:
Till eder, I man, vill jag ropa, och min röst skall utgå till människors barn.
Lären klokhet, I fåkunnige, och I dårar, lären förstånd.
Hören, ty om höga ting vill jag tala, och mina läppar skola upplåta sig till att säga vad rätt är.
Ja, sanning skall min mun tala, en styggelse för mina läppar är ogudaktighet.
Rättfärdiga äro alla min muns ord; i dem finnes intet falskt eller vrångt.
De äro alla sanna för den förståndige och rätta för dem som hava funnit kunskap.
Så tagen emot min tuktan hellre än silver, och kunskap hellre än utvalt guld.
Ty visheten är bättre än pärlor; allt vad härligt som finnes går ej upp emot henne.
Jag, visheten, är förtrogen med klokheten, och jag råder över eftertänksam insikt.
Att frukta HERREN är att hata det onda; ja, högfärd, högmod, en ond vandel och en ränkfull mun, det hatar jag.
Hos mig finnes råd och utväg; jag är förstånd, hos mig är makt.
Genom mig regera konungarna och stadga furstarna vad rätt är.
Genom mig härska härskarna och hövdingarna, ja, alla domare på jorden.
Jag älskar dem som älska mig, och de som söka mig, de finna mig.
Rikedom och ära vinnas hos mig, ädla skatter och rättfärdighet.
Min frukt är bättre än guld, ja, finaste guld och den vinning jag skänker bättre än utvalt silver.
På rättfärdighetens väg går jag fram, mitt på det rättas stigar,
till att giva dem som älska mig en rik arvedel och till att fylla deras förrådshus.
HERREN skapade mig såsom sitt förstlingsverk, i urminnes tid, innan han gjorde något annat.
Från evighet är jag insatt, från begynnelsen, ända ifrån jordens urtidsdagar.
Innan djupen voro till, blev jag född, innan källor ännu funnos, fyllda med vatten
Förrän bergens grund var lagd, förrän höjderna funnos, blev jag född,
när han ännu icke hade skapat land och mark, ej ens det första av jordkretsens stoft.
När han beredde himmelen, var jag tillstädes, när han spände ett valv över djupet,
när han fäste skyarna i höjden, när djupets källor bröto fram med makt,
när han satte för havet dess gräns, så att vattnet icke skulle överträda hans befallning, när han fastställde jordens grundvalar --
då fostrades jag såsom ett barn hos honom, då hade jag dag efter dag min lust och min lek inför hans ansikte beständigt;
jag hade min lek på hans jordkrets och min lust bland människors barn.
Så hören mig nu, I barn, ty saliga äro de som hålla mina vägar.
Hören tuktan, så att I bliven visa, ja, låten henne icke fara.
Säll är den människa som hör mig, så att hon vakar vid mina dörrar dag efter dag håller vakt vid dörrposterna i mina portar.
Ty den som finner mig, han finner livet och undfår nåd från HERREN.
Men den som går miste om mig han skadar sig själv; alla de som hata mig, de älska döden.
Visheten har byggt sig ett hus, hon har huggit ut sitt sjutal av pelare.
Hon har slaktat sin boskap, blandat sitt vin, hon har jämväl dukat sitt bord
Sina tjänarinnor har hon utsänt och låter ropa ut sin bjudning uppe på stadens översta höjder:
»Den som är fåkunnig, han komme hit.»
Ja, till den oförståndige säger hon så:
»Kommen och äten av mitt bröd, och dricken av vinet som jag har blandat.
Övergiven eder fåkunnighet, så att I fån leva, och gån fram på förståndets väg.
(Den som varnar en bespottare, han får skam igen, och den som tillrättavisar en ogudaktig får smälek därav.
Tillrättavisa icke bespottaren, på det att han icke må hata dig; tillrättavisa den som är vis, så skall han älska dig.
Giv åt den vise, så bliver han ännu visare; undervisa den rättfärdige, så lär han än mer.
HERRENS fruktan är vishetens begynnelse, och att känna den Helige är förstånd.)
Ty genom mig skola dina dagar bliva många och levnadsår givas dig i förökat mått.
Är du vis, så är din vishet dig själv till gagn, och är du en bespottare, så umgäller du det själv allena.»
En dåraktig, yster kvinna är fåkunnigheten, och intet förstå hon.
Hon har satt sig vid ingången till sitt hus, på sin stol, högt uppe i staden,
för att ropa ut sin bjudning till dem som färdas på vägen, dem som där vandra sin stig rätt fram:
»Den som är fåkunnig, han komme hit.»
Ja, till den oförståndige säger hon så:
»Stulet vatten är sött, bröd i lönndom smakar ljuvligt.»
han vet icke att det bär till skuggornas boning, hennes gäster hamna i dödsrikets djup. ----
Detta är Salomos ordspråk.
En vis son gör sin fader glädje, men en dåraktig son är sin moders bedrövelse.
Ogudaktighetens skatter gagna till intet men rättfärdigheten räddar från döden.
HERREN lämnar ej den rättfärdiges hunger omättad, men de ogudaktigas lystnad avvisar han.
Fattig bliver den som arbetar med lat hand, men de idogas hand skaffar rikedom.
En förståndig son samlar om sommaren, men en vanartig son sover i skördetiden.
Välsignelser komma över den rättfärdiges huvud, men de ogudaktigas mun gömmer på orätt.
Den rättfärdiges åminnelse lever i välsignelse, men de ogudaktigas namn multnar bort.
Den som har ett vist hjärta tager emot tillsägelser, men den som har oförnuftiga läppar går till sin undergång.
Den som vandrar i ostrafflighet, han vandrar trygg, men den som går vrånga vägar, han bliver röjd.
Den som blinkar med ögonen, han kommer ont åstad, och den som har oförnuftiga läppar går till sin undergång.
Den rättfärdiges mun är en livets källa, men de ogudaktigas mun gömmer på orätt.
Hat uppväcker trätor, men kärlek skyler allt som är brutet.
På den förståndiges läppar finner man vishet, men till den oförståndiges rygg hör ris.
De visa gömma på sin kunskap, men den oförnuftiges mun är en överhängande olycka.
Den rikes skatter äro honom en fast stad, men de armas fattigdom är deras olycka.
Den rättfärdiges förvärv bliver honom till liv; den ogudaktiges vinning bliver honom till synd.
Att taga vara på tuktan är vägen till livet, men den som ej aktar på tillrättavisning, han far vilse.
Den som gömmer på hat är en lögnare med sina läppar, och den som utsprider förtal, han är en dåre.
Där många ord äro bliver överträdelse icke borta; men den som styr sina läppar, han är förståndig.
Den rättfärdiges tunga är utvalt silver, men de ogudaktigas förstånd är föga värt.
Den rättfärdiges läppar vederkvicka många, men de oförnuftiga dö genom brist på förstånd.
Det är HERRENS välsignelse som giver rikedom, och egen möda lägger intet därtill
Dårens fröjd är att öva skändlighet, men den förståndiges är att vara vis.
Vad den ogudaktige fruktar, det vederfares honom, och vad de rättfärdiga önska, del varder dem givet.
När stormen kommer, är det ute med den ogudaktige; men den rättfärdige är en grundval som evinnerligen består.
Såsom syra för tänderna och såsom rök för ögonen, så är den late för den som har sänt honom åstad.
HERRENS fruktan förlänger livet men de ogudaktigas år varda förkortade.
De rättfärdigas väntan får en glad fullbordan, men de ogudaktigas hopp varder om intet.
HERRENS vägar äro den ostraffliges värn, men till olycka för ogärningsmännen.
Den rättfärdige skall aldrig vackla men de ogudaktiga skola icke förbliva boende i landet.
Den rättfärdiges mun bär vishet såsom frukt, men en vrång tunga bliver utrotad.
Den rättfärdiges läppar förstå vad välbehagligt är, men de ogudaktigas mun är idel vrånghet.
Falsk våg är en styggelse för HERREN, men full vikt behagar honom väl.
När högfärd kommer, kommer ock smälek, men hos de ödmjuka är vishet.
De redligas ostrafflighet vägleder dem, men de trolösas vrånghet är dem till fördärv.
Gods hjälper intet på vredens dag men rättfärdighet räddar från döden.
Den ostraffliges rättfärdighet gör hans väg jämn, men genom sin ogudaktighet faller den ogudaktige.
De redligas rättfärdighet räddar dem, men de trolösa fångas genom sin egen lystnad.
När en ogudaktig dör, varder hans hopp om intet; ja, ondskans väntan bliver om intet.
Den rättfärdige räddas ur nöden, och den ogudaktige får träda i hans ställe.
Genom sin mun fördärvar den gudlöse sin nästa, men genom sitt förstånd bliva de rättfärdiga räddade.
När det går de rättfärdiga väl, fröjdar sig staden, och när de ogudaktiga förgås, råder jubel.
Genom de redligas välsignelse varder en stad upphöjd, men genom de ogudaktigas mun brytes den ned.
Den är utan vett, som visar förakt för sin nästa; en man med förstånd tiger stilla.
Den som går med förtal, han förråder din hemlighet, den som har ett trofast hjärta döljer vad han får veta.
Där ingen rådklokhet finnes kommer folket på fall, där de rådvisa äro många, där går det väl.
En som går i borgen för en annan, honom går det illa, den som skyr att giva handslag, han är trygg.
En skön kvinna vinner ära, och våldsverkare vinna rikedom.
En barmhärtig man gör väl mot sig själv men den grymme misshandlar sitt eget kött.
Den ogudaktige gör en bedräglig vinst, men den som utsår rättfärdighet får en säker lön.
Den som står fast i rättfärdighet, han vinner liv, men den som far efter ont drager över sig död.
En styggelse för HERREN äro de vrånghjärtade, men de vilkas väg är ostrafflig behaga honom väl.
De onda bliva förvisso icke ostraffade, men de rättfärdigas avkomma får gå fri.
Såsom en gyllene ring i svinets tryne, så är skönhet hos en kvinna som saknar vett.
Vad de rättfärdiga önska får i allo en god fullbordan, men vad de ogudaktiga kunna hoppas är vrede.
Den ene utströr och får dock mer, den andre spar över hövan, men bliver allenast fattigare.
Den frikostige varder rikligen mättad, och den som vederkvicker andra, han bliver själv vederkvickt.
Den som håller inne sin säd, honom förbannar folket, den som lämnar ut sin säd, över hans huvud kommer välsignelse.
Den som vinnlägger sig om vad gott är, han strävar efter nåd, men den son söker vad ont är, över honom kommer ock ont.
Den som förtröstar på sin rikedom, han kommer på fall, men de rättfärdiga skola grönska likasom löv.
Den som drager olycka över sitt hus, han får vind till arvedel, och den oförnuftige bliver träl åt den som har ett vist hjärta.
Den rättfärdiges frukt är ett livets träd, och den som är vis, han vinner hjärtan.
Se, den rättfärdige får sin lön på jorden; huru mycket mer då den ogudaktige och syndaren!
Den som älskar tuktan, han älskar kunskap, men oförnuftig är den som hatar tillrättavisning.
Den gode undfår nåd av HERREN, men den ränkfulle varder av honom fördömd.
Ingen människa bliver beståndande genom ogudaktighet, men de rättfärdigas rot kan icke rubbas.
En idog hustru är sin mans krona, men en vanartig är såsom röta i hans ben.
De rättfärdigas tankar gå ut på vad rätt är, men de ogudaktigas rådklokhet går ut på svek.
De ogudaktigas ord ligga på lur efter blod, men de redliga räddas genom sin mun.
De ogudaktiga varda omstörtade och äro så icke mer, men de rättfärdigas hus består.
I mån av sitt vett varder en man prisad, men den som har ett förvänt förstånd, han bliver föraktad.
Bättre är en ringa man, som likväl har en tjänare, än den som vill vara förnäm och saknar bröd.
Den rättfärdige vet huru hans boskap känner det, men de ogudaktigas hjärtelag är grymt.
Den som brukar sin åker får bröd till fyllest, men oförståndig är den som far efter fåfängliga ting.
Den ogudaktige vill in i det nät som fångar de onda, men de rättfärdigas rot skjuter skott.
Den som är ond bliver snärjd i sina läppars synd, men den rättfärdige undkommer ur nöden
Sin muns frukt får envar njuta sig fullt till godo, och vad en människas händer hava förövat, det varder henne vedergällt.
Den oförnuftige tycker sin egen väg vara den rätta, med den som är vis lyssnar till råd.
Den oförnuftiges förtörnelse bliver kunnig samma dag, men den som är klok, han döljer sin skam
Den som talar vad rätt är, han främjar sanning, men ett falskt vittne talar svek.
Mången talar i obetänksamhet ord som stinga likasom svärd, men de visas tunga är en läkedom.
Sannfärdiga läppar bestå evinnerligen, men en lögnaktig tunga allenast ett ögonblick.
De som bringa ont å bane hava falskhet i hjärtat, men de som stifta frid, de undfå glädje.
Intet ont vederfares den rättfärdige, men över de ogudaktiga kommer olycka i fullt mått.
En styggelse för HERREN äro lögnaktiga låppar, men de som handla redligt behaga honom väl.
En klok man döljer sin kunskap, men dårars hjärtan ropa ut sitt oförnuft.
De idogas hand kommer till välde, men en lat hand måste göra trältjänst.
Sorg i en mans hjärta trycker det ned, men ett vänligt ord skaffar det glädje.
Den rättfärdige visar sin vän till rätta, men de ogudaktigas väg för dem själva vilse.
Den late får icke upp något villebråd, men idoghet är för människan en dyrbar skatt.
På rättfärdighetens väg är liv, och där dess stig går fram är frihet ifrån död.
En vis son hör på sin faders tuktan, men en bespottare hör icke på någon näpst.
Sin muns frukt får envar njuta sig till godo, de trolösa hungra efter våld.
Den som bevakar sin mun, han bevarar sitt liv, men den som är lösmunt kommer i olycka
Den late är full av lystnad, och han får dock intet, men de idogas hunger varder rikligen mättad.
Den rättfärdige skyr lögnaktigt tal, men den ogudaktige är förhatlig och skändlig.
Rättfärdighet bevarar den vilkens väg är ostrafflig, men ogudaktighet kommer syndarna på fall.
Den ene vill hållas för rik och har dock alls intet, den andre vill hållas för fattig och har dock stora ägodelar.
Den rike måste giva sin rikedom såsom lösepenning för sitt liv, den fattige hör icke av något
De rättfärdigas ljus brinner glatt, men de ogudaktigas lampa slocknar ut.
Genom övermod kommer man allenast split åstad, men hos dem som taga emot råd är vishet.
Lättfånget gods försvinner, men den som samlar efter hand får mycket.
Förlängd väntan tär på hjärtat, men en uppfylld önskan är ett livets träd.
Den som föraktar ordet hemfaller åt dess dom, men den som fruktar budet, han får vedergällning.
Den vises undervisning är en livets källa; genom den undviker man dödens snaror.
Ett gott förstånd bereder ynnest, men de trolösas väg är alltid sig lik.
Var och en som är klok går till väga med förstånd, men dåren breder ut sitt oförnuft.
En ogudaktig budbärare störtar i olycka, men ett tillförlitligt sändebud är en läkedom.
Fattigdom och skam får den som ej vill veta av tuktan, men den som tager vara på tillrättavisning, han kommer till ära.
Uppfylld önskan är ljuvlig för själen, men att fly det onda är en styggelse för dårar.
Hav din umgängelse med de visa, så varder du vis; den som giver sig i sällskap med dårar, honom går det illa.
Syndare förföljas av olycka, men de rättfärdiga få till lön vad gott är.
Den gode lämnar arv åt barnbarn, men syndarens gods förvaras åt den rättfärdige.
De fattigas nyodling giver riklig föda, men mången förgås genom sin orättrådighet.
Den som spar sitt ris, han hatar sin son, men den som älskar honom agar honom i tid.
Den rättfärdige får äta, så att hans hunger bliver mättad, men de ogudaktigas buk måste lida brist.
Genom visa kvinnor varder huset uppbyggt, men oförnuft river ned det med egna händer.
Den som fruktar HERREN, han vandrar i redlighet, men den som föraktar honom, han går krokiga vägar.
I den oförnuftiges mun är ett gissel för hans högmod, men de visa bevaras genom sina läppar.
Där inga dragare finnas, där förbliver krubban tom, men riklig vinning får man genom oxars kraft.
Ett sannfärdigt vittne ljuger icke, men ett falskt vittne främjar lögn.
Bespottaren söker vishet och finner ingen, men för den förståndige är kunskap lätt.
Gå bort ifrån den man som är dåraktig; aldrig fann du på hans läppar något förstånd.
Det är den klokes vishet, att han aktar på sin väg, men det är dårars oförnuft, att de öva svek.
De oförnuftiga bespottas av sitt eget skuldoffer, men bland de redliga råder gott behag.
Hjärtat känner självt bäst sin egen sorg, ej heller kan en främmande intränga i dess glädje.
De ogudaktigas hus förödes, men de rättsinnigas hydda blomstrar.
Mången håller sin väg för den i rätta, men på sistone leder den dock till döden.
Mitt under löjet kan hjärtat sörja, och slutet på glädjen bliver bedrövelse.
Av sina gärningars frukt varder den avfällige mättad, och den gode bliver upphöjd över honom.
Den fåkunnige tror vart ord, men den kloke aktar på sina steg.
Den vise tager sig till vara och flyr det onda, men dåren är övermodig och sorglös.
Den som är snar till vrede gör vad oförnuftigt är, och en ränkfull man bliver hatad.
De fåkunniga hava fått oförnuft till sin arvedel, men de kloka bliva krönta med kunskap.
De onda måste falla ned inför de goda, och de ogudaktiga vid den rättfärdiges portar.
Jämväl av sina närmaste är den fattige hatad, men den rike har många vänner.
Den som visar förakt för sin nästa, han begår synd, men säll är den som förbarmar sig över de betryckta.
De som bringa ont å bane skola förvisso fara vilse, men barmhärtighet och trofasthet röna de som bringa gott å bane.
Av all möda kommer någon vinning, men tomt tal är ren förlust.
De visas rikedom är för dem en krona men dårarnas oförnuft förbliver oförnuft.
Ett sannfärdigt vittne räddar liv, men den som främjar lögn, han är full av svek.
Den som fruktar HERREN har ett tryggt fäste, och hans barn få där en tillflykt.
I HERRENS fruktan är en livets källa genom dem undviker man dödens snaror
Att hava många undersåtar är en konungs härlighet, men brist på folk är en furstes olycka.
Den som är tålmodig visar gott förstånd, men den som är snar till vrede går långt i oförnuft.
Ett saktmodigt hjärta är kroppens liv, men bittert sinne är röta i benen.
Den som förtrycker den arme smädar hans skapare, men den som förbarmar sig över de fattiga, han ärar honom.
Genom sin ondska kommer de ogudaktige på fall, men den rättfärdige är frimodig in i döden.
I den förståndiges hjärta bor visheten, och i dårarnas krets gör hon sig kunnig.
Rättfärdighet upphöjer ett folk men synd är folkens vanära.
En förståndig tjänare behaga konungen väl, men över en vanartig skall han vrede komma.
Ett mjukt svar stillar vrede, men ett hårt ord kommer harm åstad.
De visas tunga meddelar god kunskap, men dårars mun flödar över av oförnuft.
HERRENS ögon äro överallt; de giva akt på både onda och goda.
En saktmodig tunga är ett livets träd, men en vrång tunga giver hjärtesår.
Den oförnuftige föraktar sin faders tuktan, men den som tager vara på tillrättavisning, han varder klok.
Den rättfärdiges hus gömmer stor rikedom, men i de ogudaktigas vinning är olycka.
De visas läppar strö ut kunskap, men dårars hjärtan äro icke såsom sig bör.
De ogudaktigas offer är en styggelse för HERREN, men de redligas bön behagar honom väl.
En styggelse för HERREN är den ogudaktiges väg, men den som far efter rättfärdighet, honom älskar han.
Svår tuktan drabbar den som övergiver vägen; den som hatar tillrättavisning, han måste dö.
Dödsriket och avgrunden ligga uppenbara inför HERREN; huru mycket mer då människornas hjärtan!
Bespottaren finner ej behag i tillrättavisning; till dem som äro visa går han icke.
Ett glatt hjärta gör ansiktet ljust, men vid hjärtesorg är modet brutet.
Den förståndiges hjärta söker kunskap, men dårars mun far med oförnuft.
Den betryckte har aldrig en glad dag, men ett gott mod är ett ständigt gästabud.
Bättre är något litet med HERRENS fruktan än en stor skatt med oro.
Bättre är ett fat kål med kärlek än en gödd oxe med hat.
En snarsticken man uppväcker träta, men en tålmodig man stillar kiv.
Den lates stig är såsom spärrad av törne, men de redliga hava en banad stig.
En vis son gör sin fader glädje, och en dåraktig människa är den som föraktar sin moder.
I oförnuft har den vettlöse sin glädje, men en förståndig man går sin väg rätt fram.
Där rådplägning fattas varda planerna om intet, men beståndande bliva de, där de rådvisa äro många.
En man gläder sig, när hans mun kan giva svar; ja, ett ord i sinom tid, det är gott.
Den förståndige vandrar livets väg uppåt, Då att han undviker dödsriket därnere.
Den högmodiges hus rycker HERREN bort, men änkans råmärke låter han stå fast.
För HERREN äro ondskans anslag en styggelse, men milda ord rena.
Den som söker orätt vinning drager olycka över sitt hus, men den som hatar mutor, han får leva.
Den rättfärdiges hjärta betänker vad svaras bör, men de ogudaktigas mun flödar över av onda ord.
HERREN är fjärran ifrån de ogudaktiga, men de rättfärdigas bön hör han.
En mild blick gör hjärtat glatt, ett gott budskap giver märg åt benen.
Den vilkens öra hör på hälsosam tillrättavisning, han skall få dväljas i de vises krets.
Den som ej vill veta av tuktan frågar icke efter sitt liv, men den som hör på tillrättavisning, han förvärvar förstånd.
HERRENS fruktan är en tuktan till vishet, och ödmjukhet går före ära.
En människa gör upp planer i sitt hjärta, men från HERREN kommer vad tungan svarar.
Var man tycker sina vägar vara goda, men HERREN är den som prövar andarna.
Befall dina verk åt HERREN, så hava dina planer framgång.
HERREN har gjort var sak för dess särskilda mål, så ock den ogudaktige för olyckans dag.
En styggelse för HERREN är var högmodig man; en sådan bliver förvisso icke ostraffad.
Genom barmhärtighet och trofasthet försonas missgärning, och genom HERRENS fruktan undflyr man det onda.
Om en mans vägar behaga HERREN väl så gör han ock hans fiender till hans vänner.
Bättre är något litet med rättfärdighet än stor vinning med orätt.
Människans hjärta tänker ut en väg, men HERREN är den som styr hennes steg.
Gudasvar är på konungens läppar, i domen felar icke hans mun.
Våg och rätt vägning äro från HERREN, alla vikter i pungen äro hans verk.
En styggelse för konungar äro ogudaktiga gärningar, ty genom rättfärdighet bliver tronen befäst.
Rättfärdiga läppar behaga konungar väl, Och den som talar vad rätt är, han bliver älskad.
Konungens vrede är dödens förebud, men en vis man blidkar den.
När konungen låter sitt ansikte lysa, är där liv, och hans välbehag är såsom ett moln med vårregn.
Långt bättre är att förvärva vishet än guld förstånd är mer värt att förvärvas än silver.
De redligas väg är att fly det onda; den som aktar på sin väg, han bevarar sitt liv.
Stolthet går före undergång, och högmod går före fall.
Bättre är att vara ödmjuk bland de betryckta än att utskifta byte med de högmodiga.
Den som aktar på ordet, han finner lycka, och säll är den som förtröstar på HERREN.
Den som har ett vist hjärta, honom kallar man förståndig, och där sötma är på läpparna hämtas mer lärdom.
En livets källa är förståndet för den som äger det, men oförnuftet är de oförnuftigas tuktan.
Den vises hjärta gör hans mun förståndig och lägger lärdom på hans läppar, allt mer och mer.
Milda ord äro honungskakor; de äro ljuvliga för själen och en läkedom för kroppen.
Mången håller sin väg för den rätta, men på sistone leder den dock till döden.
Arbetarens hunger hjälper honom att arbeta ty hans egen mun driver på honom.
Fördärvlig är den människa som gräver gropar för att skada; det är såsom brunne en eld på hennes läppar.
En vrång människa kommer träta åstad, och en örontasslare gör vänner oense.
Den orättrådige förför sin nästa och leder honom in på en väg som icke är god.
Den som ser under lugg, han umgås med vrånga tankar; den som biter ihop läpparna, han är färdig med något ont.
En ärekrona äro grå hår; den vinnes på rättfärdighetens väg.
Bättre är en tålmodig man än en stark, och bättre den som styr sitt sinne än den som intager en stad.
Lotten varder kastad i skötet, men den faller alltid vart HERREN vill.
Bättre är ett torrt brödstycke med ro än ett hus fullt av högtidsmat med kiv.
En förståndig tjänare får råda över en vanartig son, och bland bröderna får han skifta arv.
Degeln prövar silver och smältugnen guld, så prövar HERREN hjärtan.
En ond människa aktar på ondskefulla läppar, falskheten lyssnar till fördärvliga tungor.
Den som bespottar den fattige smädar hans skapare; den som gläder sig åt andras ofärd bliver icke ostraffad.
De gamlas krona äro barnbarn, och barnens ära äro deras fäder.
Stortaliga läppar hövas icke dåren, mycket mindre lögnaktiga läppar en furste.
En gåva är en lyckosten i dens ögon, som ger den; vart den än kommer bereder den framgång.
Den som skyler vad som är brutet, han vill främja kärlek, men den som river upp gammalt, han gör vänner oense.
En förebråelse verkar mer på den förståndige än hundra slag på dåren.
Upprorsmakaren vill allenast vad ont är, men en budbärare utan förbarmande skall sändas mot honom.
Bättre är att möta en björninna från vilken man har tagit ungarna, än att möta en dåre i hans oförnuft.
Den som vedergäller gott med ont, från hans hus skall olyckan icke vika.
Att begynna träta är att släppa ett vattenflöde löst; håll därför inne, förrän kivet har brutit ut.
Den som friar den skyldige och den som fäller den oskyldige, de äro båda en styggelse för HERREN.
Vartill gagna väl penningar i dårens hand?
Han kunde köpa sig vishet, men han saknar förstånd.
En väns kärlek består alltid. och en broder födes till hjälp i nöden.
En människa utan förstånd är den som giver handslag, den som går i borgen för sin nästa.
Den som älskar split, han älskar överträdelse; Men som bygger sin dörr hög, han far efter fall.
Den som har ett vrångt hjärta vinner ingen framgång, och den som har en förvänd tunga, han faller i olycka.
Den som har fött en dåraktig son får bedrövelse av honom, en dåres fader har ingen glädje.
Ett glatt hjärta är en god läkedom, men ett brutet mod tager märgen ur benen.
Den ogudaktige tager gärna skänker i lönndom, för att han skall vränga rättens vägar.
Den förståndige har sin blick på visheten, men dårens ögon äro vid jordens ända.
En dåraktig son är sin faders grämelse och en bitter sorg för henne som har fött honom.
Att pliktfälla jämväl den rättfärdige är icke tillbörligt; att slå ädla män strider mot rättvisan.
Den som har vett, han spar sina ord; och lugn till sinnes är en man med förstånd.
Om den oförnuftige tege, så aktades också han för vis; den som tillsluter sina läppar är förståndig.
Den egensinnige följer sin egen lystnad, med all makt söker han strid.
Dåren frågar ej efter förstånd, allenast efter att få lägga fram vad han har i hjärtat.
Där den ogudaktige kommer, där kommer förakt, och med skamlig vandel följer smälek.
Orden i en mans mun äro såsom ett djupt vatten, såsom en flödande bäck, en vishetens källa.
Att vara partisk för den skyldige är icke tillbörligt ej heller att vränga rätten för den oskyldige.
Dårens läppar komma med kiv, och hans mun ropar efter slag.
Dårens mun är honom själv till olycka, och hans läppar äro en snara hans liv.
Örontasslarens ord äro såsom läckerbitar och tränga ned till hjärtats innandömen.
Den som är försumlig i sitt arbete, han är allaredan en broder till rövaren.
HERRENS namn är ett starkt torn; den rättfärdige hastar dit och varder beskyddad.
Den rikes skatter äro honom en fast stad, höga murar likna de, i hans inbillning.
Före fall går högmod i mannens hjärta, och ödmjukhet går före ära.
Om någon giver svar, förrän han har hört, så tillräknas det honom såsom oförnuft och skam.
Mod uppehåller mannen i hans svaghet; men ett brutet mod, vem kan bära det?
Den förståndiges hjärta förvärvar kunskap, och de visas öron söka kunskap.
Gåvor öppna väg för en människa och föra henne fram inför de store.
Den som först lägger fram sin sak har rätt; sedan kommer vederparten och uppdagar huru det är.
Lottkastning gör en ände på trätor, den skiljer mellan mäktiga män.
En förorättad broder är svårare att vinna än en fast stad, och trätor äro såsom bommar för ett slott.
Av sin muns frukt får envar sin buk mättad, han varder mättad av sina läppars gröda.
Död och liv har tungan i sitt våld, de som gärna bruka henne få äta hennes frukt.
Den som har funnit en rätt hustru, han har funnit lycka och har undfått nåd av HERREN.
Bönfallande är den fattiges tal, men den rike svarar med hårda ord.
Den som ävlas att få vänner, han kommer i olycka; men vänner finnas, mer trogna än en broder.
Bättre är en fattig man som vandrar i ostrafflighet än en man som har vrånga läppar och därtill är en dåre.
Ett obetänksamt sinne, redan det är illa; och den som är snar på foten, han stiger miste.
En människas eget oförnuft kommer henne på fall, och dock är det på HERREN som hennes hjärta vredgas
Gods skaffar många vänner, men den arme bliver övergiven av sin vän.
Ett falskt vittne bliver icke ostraffat, och den som främjar lögn, han kommer icke undan.
Många söka en furstes ynnest, och alla äro vänner till den givmilde.
Den fattige är hatad av alla sina fränder, ännu längre draga sig hans vänner bort ifrån honom; han far efter löften som äro ett intet.
Den som förvärvar förstånd har sitt liv kärt; den som tager vara på insikt, han finner lycka
Ett falskt vittne bliver icke ostraffat, och den som främjar lögn, han skall förgås.
Det höves icke dåren att hava goda dagar, mycket mindre en träl att råda över furstar.
Förstånd gör en människa tålmodig, och det är hennes ära att tillgiva vad någon har brutit.
En konungs vrede är såsom ett ungt lejons rytande, hans nåd är såsom dagg på gräset.
En dåraktig son är sin faders fördärv, och en kvinnas trätor äro ett oavlåtligt takdropp.
Gård och gods får man i arv från sina fäder, men en förståndig hustru är en gåva från HERREN.
Lättja försänker i dåsighet, och den håglöse får lida hunger.
Den som håller budet får behålla sitt liv; den som ej aktar på sin vandel han varder dödad.
Den som förbarmar sig över den arme, han lånar åt HERREN och får vedergällning av honom för vad gott han har gjort.
Tukta din son, medan något hopp är, och åtrå icke att vålla hans död.
Den som förgår sig i vrede, han må plikta därför, ty om du vill ställa till rätta, så gör du det allenast värre.
Hör råd och tag emot tuktan, på det att du för framtiden må bliva vis.
Många planer har en man i sitt hjärta, men HERRENS råd, det bliver beståndande.
Efter en människas goda vilja räknas hennes barmhärtighet, och en fattig man är bättre än en som ljuger.
HERRENS fruktan för till liv; så får man vila mätt och hemsökes icke av något ont.
Den late sticker sin hand i fatet, men gitter icke föra den åter till munnen.
Slår man bespottaren, så bliver den fåkunnige klok; och tillrättavisar man den förståndige, så vinner han kunskap.
Den som övar våld mot sin fader eller driver bort sin moder, han är en vanartig och skändlig son.
Min son, om du icke vill höra tuktan, så far du vilse från de ord som giva kunskap.
Ett ont vittne bespottar vad rätt är, och de ogudaktigas mun är glupsk efter orätt.
Straffdomar ligga redo för bespottarna och slag för dårarnas rygg.
En bespottare är vinet, en larmare är rusdrycken, och ovis är envar som raglar därav.
Såsom ett ungt lejons rytande är den skräck en konung ingiver; den som ådrager sig hans vrede har förverkat sitt liv.
Det är en ära för en man att hålla sig ifrån kiv, den oförnuftige söker alltid strid.
När hösten kommer, vill den late icke plöja; därför söker han vid skördetiden förgäves efter frukt.
Planerna i en mans hjärta äro såsom ett djupt vatten, men en man med förstånd hämtar ändå upp dem.
Många finnas, som ropa ut var och en sin barmhärtighet; men vem kan finna en man som är att lita på?
Den som vandrar i ostrafflighet såsom en rättfärdig man, hans barn går det val efter honom.
En konung, som sitter på domarstolen, rensar med sina ögons kastskovel bort allt vad ont är.
Vem kan säga: »Jag har bevarat mitt hjärta rent, jag är fri ifrån synd»?
Två slags vikt och två slags mått, det ena som det andra är en styggelse för HERREN.
Redan barnet röjer sig i sina gärningar, om dess vandel är rättskaffens och redlig.
Örat, som hör, och ögat, som ser, det ena som det andra har HERREN gjort.
Älska icke sömn, på det att du icke må bliva fattig; håll dina ögon öppna, så får du bröd till fyllest.
»Uselt, uselt», säger köparen; men när han går sin väg, rosar han sitt köp.
Man må hava guld, så ock pärlor i myckenhet, den dyrbaraste klenoden äro dock läppar som tala förstånd.
Tag kläderna av honom, ty han har gått i borgen för en annan, och panta ut vad han har, för de främmandes skull.
Orättfånget bröd smakar mannen ljuvligt, men efteråt bliver hans mun full av stenar.
Planer hava framgång, när de äro väl överlagda, och med rådklokhet må man föra krig.
Den som går med förtal, han förråder hemligheter; med den som är lösmunt må du ej giva dig i lag.
Den som uttalar förbannelser över fader eller moder, hans lampa skall slockna ut mitt i mörkret.
Det förvärv man i förstone ävlas efter, det varder på sistone icke välsignat.
Säg icke: »Jag vill vedergälla ont med ont»; förbida HERREN, han skall hjälpa dig.
Tvåfaldig vikt är en styggelse för HERREN, och falsk våg är icke något gott.
Av HERREN bero en mans steg; ja, en människa förstår icke själv sin väg.
Det är farligt för en människa att obetänksamt helga något och att överväga sina löften, först när de äro gjorda.
En vis konung rensar bort de ogudaktiga såsom med en kastskovel och låter tröskhjulet gå över dem.
Anden i människan är en HERRENS lykta; den utrannsakar alla hjärtats innandömen.
Mildhet och trofasthet äro en konungs vakt; genom mildhet stöder han sin tron.
De ungas ära är deras kraft, och de gamlas prydnad äro deras grå hår.
Sår som svida rena från ondska, ja, tuktan renar hjärtats innandömen.
Konungars hjärtan äro i HERRENS hand såsom vattenbäckar: han leder dem varthelst han vill.
Var man tycker sin väg vara den rätta, men HERREN är den som prövar hjärtan.
Att öva rättfärdighet och rätt, det är mer värt för HERREN än offer.
Stolta ögon och högmodigt hjärta -- de ogudaktigas lykta är dem till synd.
Den idoges omtanke leder allenast till vinning, men all fikenhet allenast till förlust.
De skatter som förvärvas genom falsk tunga, de äro en försvinnande dunst och hasta till döden.
De ogudaktigas övervåld bortrycker dem själva, eftersom de icke vilja göra vad rätt är.
En oärlig mans väg är idel vrånghet, men en rättskaffens man handla redligt
Bättre är att bo i en vrå på taket än att hava hela huset gemensamt med en trätgirig kvinna.
Den ogudaktiges själ har lust till det onda; hans nästa finner ingen barmhärtighet hos honom.
Straffar man bespottaren, så bliver den fåkunnige vis: och undervisar man den vise, så inhämtar han kunskap.
Den Rättfärdige giver akt på den ogudaktiges hus, han störtar de ogudaktiga i olycka.
Den som tillsluter sitt öra för den armes rop, han skall själv ropa utan att få svar.
En hemlig gåva stillar vrede och en skänk i lönndom våldsammaste förbittring.
Det är den rättfärdiges glädje att rätt skipa, men det är ogärningsmännens skräck.
Den människa som far vilse ifrån förståndets väg, hon hamnar i skuggornas krets.
Den som älskar glada dagar varder fattig; den som älskar vin och olja bliver icke rik.
Den ogudaktige varder given såsom lösepenning för den rättfärdige, och den trolöse sättes i de redligas ställe.
Bättre är att bo i ett öde land än med en trätgirig och besvärlig kvinna.
Dyrbara skatter och salvor har den vise i sin boning, men en dåraktig människa förslösar sitt gods.
Den som far efter rättfärdighet och godhet, han finner liv, rättfärdighet och ära.
En vis man kan storma en stad full av hjältar och bryta ned det fäste som var dess förtröstan.
Den som besvarar sin mun och sin tunga han bevarar sitt liv för nöd.
Bespottare må den kallas, som är fräck och övermodig, den som far fram med fräck förmätenhet.
Den lates begärelse för honom till döden, i det att hans händer icke vilja arbeta.
Den snikne är alltid full av snikenhet; men den rättfärdige giver och spar icke.
De ogudaktigas offer är en styggelse; mycket mer, när det frambäres i skändligt uppsåt.
Ett lögnaktigt vittne skall förgås; men en man som hör på får allt framgent tala.
En ogudaktig man uppträder fräckt; men den redlige vandrar sina vägar ståndaktigt.
Ingen vishet, intet förstånd, intet råd förmår något mot HERREN.
Hästar rustas ut för stridens dag, men från HERREN är det som segern kommer.
Ett gott namn är mer värt än stor rikedom, ett gott anseende är bättre än silver och guld.
Rik och fattig få leva jämte varandra; HERREN har gjort dem båda.
Den kloke ser faran och söker skydd; men de fåkunniga löpa åstad och få plikta därför.
Ödmjukhet har sin lön i HERRENS fruktan, i rikedom, ära och liv.
Törnen och snaror ligga på den vrånges väg; den som vill bevara sitt liv håller sig fjärran ifrån dem.
Vänj den unge vid den väg han bör vandra, så viker han ej därifrån, när han bliver gammal.
Den rike råder över de fattiga, och låntagaren bliver långivarens träl.
Den som sår vad orätt är, han får skörda fördärv, och hans övermods ris får en ände.
Den som unnar andra gott, han varder välsignad, ty han giver av sitt bröd åt den arme.
Driv ut bespottaren, så upphör trätan, och tvist och smädelse få en ände.
Den som älskar hjärtats renhet, den vilkens läppar tala ljuvligt, hans vän är konungen.
HERRENS ögon bevara den förståndige; därför omstörtar han den trolöses planer.
Den late säger: »Ett lejon är på gatan; därute på torget kunde jag bliva dräpt.»
En trolös kvinnas mun är en djup grop; den som har träffats av HERRENS vrede, han faller däri.
Oförnuft låder vid barnets hjärta, men tuktans ris driver det bort.
Den som förtrycker den arme bereder honom vinning men den som giver åt den rike vållar honom allenast förlust. ----
Böj ditt öra härtill, och hör de vises ord, och lägg mina lärdomar på hjärtat.
Ty det bliver dig ljuvligt, om du bevarar dem i ditt innersta; må de alla ligga redo på dina läppar.
För att du skall sätta din förtröstan till HERREN, undervisar jag i dag just dig.
Ja, redan förut har jag ju skrivit regler för dig och meddelat dig råd och insikt,
för att lära dig tillförlitliga sanningsord, så att du rätt kan svara den som har sänt dig åstad.
Plundra icke den arme, därför att han är arm, och förtrampa icke den fattige porten.
Ty HERREN skall utföra deras sak, och dem som röva från dem skall han beröva livet.
Giv dig icke i sällskap med den som lätt vredgas eller i lag med en snarsticken man,
på det att du icke må lära dig hans vägar och bereda en snara för ditt liv.
Var icke en av dem som giva handslag, en av dem som gå i borgen för lån.
Icke vill du att man skall taga ifrån dig sängen där du ligger, om du icke har något att betala med?
Flytta icke ett gammalt råmärke, ett sådant som dina fäder hava satt upp.
Ser du en man som är väl förfaren i sin syssla, hans plats är att tjäna konungar; icke må han tjäna ringa män.
När du sitter till bords med en furste, så besinna väl vad du har framför dig,
och sätt en kniv på din strupe, om du är alltför hungrig.
Var ej lysten efter hans smakliga rätter, ty de äro en bedräglig kost.
Möda dig icke för att bliva rik; avstå från att bruka klokskap.
Låt icke dina blickar flyga efter det som ej har bestånd; ty förvisso gör det sig vingar och flyger sin väg, såsom örnen mot himmelen.
Ät icke den missunnsammes bröd, och var ej lysten efter hans smakliga rätter;
ty han förfar efter sina själviska beräkningar. »Ät och drick» kan han val säga till dig, men hans hjärta är icke med dig.
Den bit du har ätit måste du utspy, och dina vänliga ord har du förspillt.
Tala icke för en dåres öron, ty han föraktar vad klokt du säger.
Flytta icke ett gammalt råmärke, och gör icke intrång på de faderlösas åkrar.
Ty deras bördeman är stark; han skall utföra deras sak mot dig.
Vänd ditt hjärta till tuktan och dina öron till de ord som giva kunskap.
Låt icke gossen vara utan aga; ty om du slår honom med riset, så bevaras han från döden;
ja, om du slår honom med riset, så räddar du hans själ undan dödsriket.
Min son, om ditt hjärta bliver vist, så gläder sig ock mitt hjärta;
ja, mitt innersta fröjdar sig, när dina läppar tala vad rätt är.
Låt icke ditt hjärta avundas syndare, men nitälska för HERRENS fruktan beständigt.
Förvisso har du då en framtid, och ditt hopp varder icke om intet.
Hör, du min son, och bliv vis, och låt ditt hjärta gå rätta vägar.
Var icke bland vindrinkare, icke bland dem som äro överdådiga i mat.
Ty drinkare och frossare bliva fattiga, och sömnaktighet giver trasiga kläder.
Hör din fader, som har fött dig, och förakta icke din moder, när hon varder gammal.
Sök förvärva sanning, och avhänd dig henne icke, sök vishet och tukt och förstånd.
Stor fröjd har den rättfärdiges fader; den som har fått en vis son har glädje av honom.
Må då din fader och din moder få glädje, och må hon som har fött dig kunna fröjda sig.
Giv mig, min son, ditt hjärta, och låt mina vägar behaga dina ögon.
Ty skökan är en djup grop, och nästans hustru är en trång brunn.
Ja, såsom en rövare ligger hon på lur och de trolösas antal förökar hon bland människorna.
Var är ve, var är jämmer?
Var äro trätor, var är klagan?
Var äro sår utan sak?
Var äro ögon höljda i dunkel?
Jo, där man länge sitter kvar vid vinet, där man samlas för att pröva kryddade drycker.
Så se då icke på vinet, att det är så rött, att det giver sådan glans i bägaren, och att det så lätt rinner ned.
På sistone stinger det ju såsom ormen, och likt basilisken sprutar det gift.
Dina ögon få då skåda sällsamma syner, och ditt hjärta talar förvända ting.
Det är dig såsom låge du i havets djup, eller såsom svävade du uppe i en mast:
»De slå mig, men åt vållar mig ingen smärta, de stöta mig, men jag känner det icke.
När skall jag då vakna upp, så att jag återigen får skaffa mig sådant?»
Avundas icke onda människor, och hav ingen lust till att vara med dem.
Ty på övervåld tänka deras hjärtan, och deras läppar tala olycka.
Genom vishet varder ett hus uppbyggt, och genom förstånd hålles det vid makt.
Genom klokhet bliva kamrarna fyllda med allt vad dyrbart och ljuvligt är.
En vis man är stark, och en man med förstånd är väldig i kraft.
Ja, med rådklokhet skall man föra krig, och där de rådvisa äro många, där går det väl.
Sällsynt korall är visheten för den oförnuftige, i porten kan han icke upplåta sin mun.
Den som tänker ut onda anslag, honom må man kalla en ränksmidare.
Ett oförnuftigt påfund är synden, och bespottaren är en styggelse för människor.
Låter du modet falla, när nöd kommer på, så saknar du nödig kraft.
Rädda dem som släpas till döden, och bistå dem som stappla till avrättsplatsen.
Om du säger: »Se, vi visste det icke», så betänk om ej han som prövar hjärtan märker det, och om ej han som har akt på din själ vet det.
Och han skall vedergälla var och en efter hans gärningar.
Ät honung, min son, ty det är gott, och självrunnen honung är söt för din mun.
Lik sådan må du räkna visheten för din själ.
Om du finner henne, så har du en framtid, och ditt hopp varder då icke om intet.
Lura icke, du ogudaktige, på den rättfärdiges boning, öva intet våld mot hans vilostad.
Ty den rättfärdige faller sju gånger och står åter upp; men de ogudaktiga störta över ända olyckan.
Gläd dig icke, när din fiende faller, och låt ej ditt hjärta fröjda sig, när han störtar över ända,
på det att HERREN ej må se det med misshag och flytta sin vrede ifrån honom.
Harmas icke över de onda, avundas icke de ogudaktiga.
Ty den som är ond har ingen framtid; de ogudaktigas lampa skall slockna ut.
Min son, frukta HERREN och konungen; giv dig icke i lag med upprorsmän.
Ty plötsligt skall ofärd komma över dem, och vem vet när deras år få en olycklig ände? ----
Dessa ord äro ock av visa män.
Att hava anseende till personen, när man dömer, är icke tillbörligt.
Den som säger till den skyldige: »Du är oskyldig», honom skola folk förbanna, honom skola folkslag önska ofärd.
Men dem som skipa rättvisa skall det gå väl, och över dem skall komma välsignelse av vad gott är.
En kyss på läpparna är det, när någon giver ett rätt svar.
Fullborda ditt arbete på marken, gör allting redo åt dig på åkern; sedan må du bygga dig bo.
Bär icke vittnesbörd mot din nästa utan sak; icke vill du bedraga med dina läppar?
Säg icke: »Såsom han gjorde mot mig vill jag göra mot honom, jag vill vedergälla mannen efter hans gärningar.»
Jag gick förbi en lat mans åker, en oförståndig människas vingård.
Och se, den var alldeles full av ogräs, dess mark var övertäckt av nässlor, och dess stenmur låg nedriven.
Och jag betraktade det och aktade därpå, jag såg det och tog varning därav.
Ja, sov ännu litet, slumra ännu litet, lägg ännu litet händerna i kors för att vila,
så skall fattigdomen komma farande över dig, och armodet såsom en väpnad man.
Dessa ordspråk äro ock av Salomo; och Hiskias, Juda konungs, män hava gjort detta utdrag.
Det är Guds ära att fördölja en sak, men konungars ära att utforska en sak.
Himmelens höjd och jordens djup och konungars hjärtan kan ingen utrannsaka.
Skaffa slagget bort ifrån silvret, så får guldsmeden fram en klenod därav.
Skaffa de ogudaktiga bort ur konungens tjänst, så varder hans tron befäst genom rättfärdighet.
Förhäv dig icke inför konungen, och träd icke fram på de stores plats.
Ty det är bättre att man säger till dig: »Stig hitupp», än att man flyttar ned dig för någon förnämligare man, någon som dina ögon redan hava sett.
Var icke för hastig att begynna en tvist; vad vill du eljest göra längre fram, om din vederpart kommer dig på skam?
Utför din egen sak mot din vederpart, men uppenbara icke en annans hemlighet,
på det att icke envar som hör det må lasta dig och ditt rykte bliva ont för beständigt.
Gyllene äpplen i silverskålar äro ord som talas i rättan tid.
Såsom en gyllene örring passar till ett bröstspänne av fint guld, så passar en vis bestraffare till ett hörsamt öra.
Såsom snöns svalka på en skördedag, så är en pålitlig budbärare för avsändaren; sin herres själ vederkvicker han.
Såsom regnskyar och blåst, och likväl intet regn, så är en man som skryter med givmildhet, men icke håller ord.
Genom tålamod varder en furste bevekt, och en mjuk tunga krossar ben.
Om du finner honung, så ät icke mer än du tål, så att du ej bliver övermätt därav och får utspy den.
Låt din fot icke för ofta komma i din väns hus, Så att han ej bliver mätt på dig och får motvilja mot dig.
En stridshammare och ett svärd och en skarp pil är den som bär falskt vittnesbörd mot sin nästa.
Såsom en gnagande tand och såsom ett skadedjurs fot är den trolöses tillförsikt på nödens dag.
Såsom att taga av dig manteln på en vinterdag, och såsom syra på lutsalt, så är det att sjunga visor för ett sorgset hjärta.
Om din ovän är hungrig, så giv honom att äta, och om han är törstig, så giv honom att dricka;
så samlar du glödande kol på hans huvud, och HERREN skall vedergälla dig.
Nordanvind föder regn och en tasslande tunga mulna ansikten.
Bättre är att bo i en vrå på taket än att hava hela huset gemensamt med en trätgirig kvinna.
Såsom friskt vatten för den försmäktande, så är ett gott budskap ifrån fjärran land.
Såsom en grumlad källa och en fördärvad brunn, så är en rättfärdig som vacklar inför den ogudaktige.
Att äta för mycket honung är icke gott, och den som vinner ära får sin ära nagelfaren.
Såsom en stad vars murar äro nedbrutna och borta, så är en man som icke kan styra sitt sinne.
Såsom snö icke hör till sommaren och regn icke till skördetiden, så höves det ej heller att dåren får ära.
Såsom sparven far sin kos, och såsom svalan flyger bort, så far en oförtjänt förbannelse förbi.
Piskan för hästen, betslet för åsnan och riset för dårarnas rygg!
Svara icke dåren efter hans oförnuft, så att du icke själv bliver honom lik.
Svara dåren efter hans oförnuft, för att han icke må tycka sig vara vis.
Den som sänder bud med en dåre, han hugger själv av sig fötterna, och får olycka till dryck.
Lika den lames ben, som hänga kraftlösa ned, äro ordspråk i dårars mun.
Såsom att binda slungstenen fast vid slungan, så är det att giva ära åt en dåre.
Såsom när en törntagg kommer i en drucken mans hand, så är det med ordspråk i dårars mun.
En mästare gör själv allt, men dåren lejer, och lejer vem som kommer.
Lik en hund som vänder åter till i sina spyor dåre som på nytt begynner sitt oförnuft.
Ser du en man som tycker sig själv vara vis, det är mer hopp om en dåre än om honom.
Den late säger: »Ett vilddjur är på vägen, ja, ett lejon är på gatorna.
Dörren vänder sig på sitt gångjärn, och den late vänder sig i sin säng.
Den late sticker sin hand i fatet, men finner det mödosamt att föra den åter till munnen.
Den late tycker sig vara vis, mer än sju som giva förståndiga svar.
Lik en som griper en hund i öronen är den som förivrar sig vid andras kiv, där han går fram.
Lik en rasande, som slungar ut brandpilar och skjuter och dödar,
är en man som bedrager sin nästa och sedan säger: »Jag gjorde det ju på skämt.»
När veden tager slut, slocknar elden. och när örontasslaren är borta, stillas trätan.
Såsom glöd kommer av kol, och eld av ved, så upptändes kiv av en trätgirig man.
Örontasslarens ord äro såsom läckerbitar och tränga ned till hjärtats innandömen.
Såsom silverglasering på ett söndrigt lerkärl äro kärleksglödande läppar, där hjärtat är ondskefullt.
En fiende förställer sig i sitt tal, men i sitt hjärta bär han på svek.
Om han gör sin röst ljuvlig, så tro honom dock icke, ty sjufaldig styggelse är i hans hjärta.
Hatet brukar list att fördölja sig med, men den hatfulles ondska varder dock uppenbar i församlingen.
Den som gräver en grop, han faller själv däri, och den som vältrar upp en sten, på honom rullar den tillbaka.
En lögnaktig tunga hatar dem hon har krossat, och en hal mun kommer fall åstad.
Beröm dig icke av morgondagen, ty du vet icke vad en dag kan bära i sitt sköte.
Må en annan berömma dig, och icke din egen mun, främmande, och icke dina egna läppar.
Sten är tung, och sand är svår att bära, men tyngre än båda är förargelse genom en oförnuftig man.
Vrede är en grym sak och harm en störtflod, men vem kan bestå mot svartsjuka?
Bättre är öppen tillrättavisning än kärlek som hålles fördold.
Vännens slag givas i trofasthet, men ovännens kyssar till överflöd.
Den mätte trampar honung under fötterna, men den hungrige finner allt vad bittert är sött.
Lik en fågel som har måst fly ifrån sitt bo är en man som har måst fly ifrån sitt hem.
Salvor och rökelse göra hjärtat glatt, ömhet hos en vän som giver välbetänkta råd.
Din vän och din faders vän må du icke låta fara, gå icke till din broders hus, när ofärd drabbar dig; bättre är en granne som står dig nära än broder som står dig fjärran.
Bliv vis, min son, så gläder du mitt hjärta; jag kan då giva den svar, som smädar mig.
Den kloke ser faran och söker skydd; de fåkunniga löpa åstad och få plikta därför.
Tag kläderna av honom, ty han har gått i borgen för en annan, och panta ut vad han har, för den främmande kvinnans skull.
Den som välsignar sin nästa med hög röst bittida om morgonen, honom kan det tillräknas såsom en förbannelse.
Ett oavlåtligt takdropp på en regnig dag och en trätgirig kvinna, det kan aktas lika.
Den som vill lägga band på en sådan vill lägga band på vinden, och hala oljan möter hans högra hand.
Järn giver skärpa åt järn; så skärper den ena människan den andra.
Den som vårdar sitt fikonträd, han får äta dess frukt; och den som vårdar sig om sin herre, han kommer till ära.
Såsom spegelbilden i vattnet liknar ansiktet, så avspeglar den ena människans hjärta den andras.
Dödsriket och avgrunden kunna icke mättas; så bliva ej heller människans ögon mätta.
Silvret prövas genom degeln och guldet genom smältugnen, så ock en man genom sitt rykte.
Om du stötte den oförnuftige mortel med en stöt, bland grynen, så skulle hans oförnuft ändå gå ur honom.
Se väl till dina får, och hav akt på dina hjordar.
Ty rikedom varar icke evinnerligen; består ens en krona från släkte till släkte?
När ny brodd skjuter upp efter gräset som försvann, och när foder samlas in på bergen,
då äger du lamm till att bereda dig kläder och bockar till att köpa dig åker;
då giva dig getterna mjölk nog, till föda åt dig själv och ditt hus och till underhåll åt dina tjänarinnor.
De ogudaktiga fly, om ock ingen förföljer dem; men de rättfärdiga äro oförskräckta såsom unga lejon.
För sin överträdelses skull får ett land många herrar; men där folket har förstånd och inser vad rätt är, där bliver det beståndande.
En usel herre, som förtrycker de arma, är ett regn som förhärjar i stället för att giva bröd.
De som övergiva lagen prisa de ogudaktiga, men de som hålla lagen gå till strids mot dem.
Onda människor förstå icke vad rätt är, men de som söka HERREN, de förstå allt.
Bättre är en fattig man som vandrar i ostrafflighet rik som i vrånghet går dubbla vägar.
Den yngling är förståndig, som tager lagen i akt; men som giver sig i sällskap med slösare gör sin fader skam.
De som förökar sitt gods genom ocker och räntor, han samlar åt den som förbarmar sig över de arma.
Om någon vänder bort sitt öra och icke vill höra lagen, så är till och med hans bön en styggelse.
Den som leder de redliga vilse in på en ond väg, han faller själv i sin grop; men de ostraffliga få till sin arvedel vad gott är.
En rik man tycker sig vara vis, men en fattig man med förstånd uppdagar hurudan han är.
När de rättfärdiga triumfera, står allt härligt till; men när de ogudaktiga komma till makt, får man leta efter människor.
Den som fördöljer sina överträdelser, honom går det icke väl; men den som bekänner och övergiver dem, han får barmhärtighet.
Säll är den människa som ständigt tager sig till vara; men den som förhärdar sitt hjärta, han faller i olycka.
Lik ett rytande lejon och en glupande björn är en ogudaktig furste över ett fattigt folk.
Du furste utan förstånd, du som övar mycket våld, att den som hatar orätt vinning, han skall länge leva.
En människa som tryckes av blodskuld bliver en flykting ända till sin grav, och ingen må hjälpa en sådan.
Den som vandrar ostraffligt, han bliver frälst; men den som i vrånghet går dubbla vägar, han faller på en av dem.
Den som brukar sin åker får bröd till fyllest; men den som far efter fåfängliga ting får fattigdom till fyllest.
En redlig man får mycken välsignelse; men den som fikar efter att varda rik, kan bliver icke ostraffad.
Att hava anseende till personen är icke tillbörligt; men för ett stycke bröd gör sig mången till överträdare.
Den missunnsamme ävlas efter ägodelar och förstår icke att brist skall komma över honom.
Den som tillrättavisar en avfälling skall vinna ynnest, mer än den som gör sin tunga hal.
Den som plundrar sin fader eller sin moder och säger: »Det är ingen synd», han är stallbroder till rövaren.
Den som är lysten efter vinning uppväcker träta; men den som förtröstar på HERREN varder rikligen mättad.
Den som förlitar sig på sitt förstånd, han är en dåre; men den som vandrar i vishet, han bliver hulpen.
Den som giver åt den fattige, honom skall intet fattas; men den som tillsluter sina ögon drabbas av mycken förbannelse.
När de ogudaktiga komma till makt, gömma sig människorna; men när de förgås, växa de rättfärdiga till.
Den som får mycken tillrättavisning, men förbliver hårdnackad, han varder oförtänkt krossad utan räddning.
När de rättfärdiga växa till, gläder sig folket, men när den ogudaktige kommer till välde, suckar folket.
Den som älskar vishet gör sin fader glädje; men den som giver sig i sällskap med skökor förstör vad han äger.
Genom rättvisa håller en konung sitt land vid makt; men den som utpressar gärder, har fördärvar det.
Den man som smickrar sin nästa han breder ut ett nät för han fötter.
En ond människas överträdelse bliver henne en snara, men den rättfärdige får jubla och glädjas.
Den rättfärdige vårdar sig om de armas sak, men den ogudaktige förstår intet.
Bespottare uppvigla staden, men visa män stilla vreden.
När en vis man vill gå till rätta med en oförnuftig man, då vredgas denne eller ler, och har ingen ro.
De blodgiriga hata den som är ostrafflig, men de redliga söka skydda hans liv.
Dåren släpper all sin vrede lös, men den vise stillar den till slut.
Den furste som aktar på lögnaktigt tal, hans tjänare äro alla ogudaktiga.
Den fattige och förtryckaren få leva jämte varandra; av HERREN få bådas ögon sitt ljus.
Den konung som dömer de armas rätt. hans tron skall bestå evinnerligen.
Ris och tillrättavisning giver vishet, men ett oupptuktat barn drager skam över sin moder.
Där de ogudaktiga växa till, där växer överträdelsen till, men de rättfärdiga skola se deras fall med lust.
Tukta din son, så skall han bliva dig till hugnad och giva ljuvlig spis åt din själ.
Där profetia icke finnes, där bliver folket tygellöst; men säll är den som håller lagen.
Med ord kan man icke tukta en tjänare ty om han än förstår, så rättar han sig icke därefter.
Ser du en man som är snar till att tala, det är mer hopp om en dåre än om honom.
Om någon är för efterlåten mot sin tjänare i hans ungdom, så visar denne honom på sistone förakt.
En snarsticken man uppväcker träta, och den som lätt förtörnas begår ofta överträdelse.
En människas högmod bliver henne till förödmjukelse, men den ödmjuke vinner ära.
Den som skiftar rov med en tjuv hatar sitt eget liv; när han hör edsförpliktelsen, yppar han intet.
Människofruktan har med sig snaror, men den som förtröstar på HERREN, han varder beskyddad.
Många söka en furstes ynnest, men av HERREN får var och en sin rätt.
En orättfärdig man är en styggelse för de rättfärdiga, och den som vandrar i redlighet är en styggelse för den ogudaktige.
Detta är Agurs, Jakes sons, ord och utsaga.
Så talade den mannen till Itiel -- till Itiel och Ukal.
Ja, jag är för oförnuftig för att kunna räknas såsom människa, jag har icke mänskligt förstånd;
vishet har jag icke fått lära, så att jag äger kunskap om den Helige.
Vem har stigit upp till himmelen och åter farit ned?
Vem har samlat vinden i sina händer?
Vem har knutit in vattnet i ett kläde?
Vem har fastställt jordens alla gränser?
Vad heter han, och vad heter hans son -- du vet ju det?
Allt Guds tal är luttrat; han är en sköld för dem som taga sin tillflykt till honom.
Lägg icke något till hans ord, på det att han icke må beslå dig med lögn.
Om två ting beder jag dig, vägra mig dem icke, intill min död:
Låt fåfänglighet och lögn vara fjärran ifrån mig; och giv mig icke fattigdom, ej heller rikedom, men låt mig få det bröd mig tillkommer.
Jag kunde eljest, om jag bleve alltför matt, förneka dig, att jag sporde: »Vem är HERREN?» eller om jag bleve alltför fattig, kunde jag bliva en tjuv, ja, förgripa mig på min Guds namn.
Förtala icke en tjänare inför hans herre; han kunde eljest förbanna dig, så att du stode där med skam.
Ett släkte där man förbannar sin fader, och där man icke välsignar sin moder;
ett släkte som tycker sig vara rent, fastän det icke har avtvått sin orenlighet;
ett släkte -- huru stolta äro icke dess ögon, och huru fulla av högmod äro icke dess blickar!
ett släkte vars tänder äro svärd, och vars kindtänder äro knivar, så att de äta ut de betryckta ur landet och de fattiga ur människornas krets!
Blodigeln har två döttrar: »Giv hit, giv hit.»
Tre finnas, som icke kunna mättas, ja, fyra, som aldrig säga: »Det är nog»:
dödsriket och den ofruktsammas kved, jorden, som icke kan mättas med vatten, och elden, som aldrig säger: »Det är nog.»
Den som bespottar sin fader och försmår att lyda sin moder hans öga skola korparna vid bäcken hacka ut, och örnens ungar skola äta upp det.
Tre ting äro mig för underbara, ja, fyra finnas, som jag icke kan spåra:
örnens väg under himmelen, ormens väg över klippan, skeppets väg mitt i havet och en mans väg hos en ung kvinna.
Sådant är äktenskapsbryterskans sätt: hon njuter sig mätt och stryker sig så om munnen och säger: »Jag har intet orätt gjort.»
Tre finnas, under vilka jorden darrar, ja, fyra, under vilka den ej kan uthärda:
under en träl, när han bliver konung, och en dåre, när han får äta sig mätt,
under en försmådd kvinna, när hon får man och en tjänstekvinna, när hon tränger undan sin fru.
Fyra finnas, som äro små på jorden, och likväl är stor vishet dem beskärd:
myrorna äro ett svagt folk, men de bereda om sommaren sin föda;
klippdassarna äro ett folk med ringa kraft, men i klippan bygga de sig hus;
gräshopporna hava ingen konung, men i härordning draga de alla ut;
gecko-ödlan kan gripas med händerna, dock bor hon i konungapalatser.
Tre finnas, som skrida ståtligt fram, ja, fyra, som hava en ståtlig gång:
lejonet, hjälten bland djuren, som ej viker tillbaka för någon,
en stridsrustad häst och en bock och en konung i spetsen för sin här.
Om du har förhävt dig, evad det var dårskap eller det var medveten synd, så lägg handen på munnen.
Ty såsom ost pressas ut ur mjölk, och såsom blod pressas ut ur näsan, så utpressas kiv ur vrede. ----
Detta är konung Lemuels ord, vad hans moder sade, när hon förmanade honom:
Hör, min son, ja, hör, du mitt livs son, hör, du mina löftens son.
Giv icke din kraft åt kvinnor, vänd icke dina vägar till dem som äro konungars fördärv.
Ej konungar tillkommer det, Lemoel, ej konungar tillkommer det att dricka vin ej furstar att fråga efter starka drycker.
De kunde eljest under sitt drickande förgäta lagen och förvända rätten för alla eländets barn.
Nej, åt den olycklige give man starka drycker och vin åt dem som hava en bedrövad själ.
Må dessa dricka och förgäta sitt armod och höra upp att tänka på sin vedermöda.
Upplåt din mun till förmån för den stumme och till att skaffa alla hjälplösa rätt.
Ja, upplåt din mun och döm med rättvisa, och skaffa den betryckte och fattige rätt. ----
En idog hustru, var finner man en sådan?
Långt högre än pärlor står hon i pris.
På henne förlitar sig hennes mans hjärta, och bärgning kommer icke att fattas honom.
Hon gör honom vad ljuvt är och icke vad lett är, i alla sina levnadsdagar.
Omsorg har hon om ull och lin och låter sina händer arbeta med lust.
Hon är såsom en köpmans skepp, sitt förråd hämtar hon fjärran ifrån.
Medan det ännu är natt, står hon upp och sätter fram mat åt sitt husfolk, åt tjänarinnorna deras bestämda del.
Hon har planer på en åker, och hon skaffar sig den; av sina händers förvärv planterar hon en vingård.
Hon omgjordar sina länder med kraft och lägger driftighet i sina armar.
Så förmärker hon att hennes hushållning går väl; hennes lampa släckes icke ut om natten.
Till spinnrocken griper hon med sina händer, och hennes fingrar fatta om sländan.
För den betryckte öppnar hon sin hand och räcker ut sina armar mot den fattige.
Av snötiden fruktar hon intet för sitt hus, ty hela hennes hus har kläder av scharlakan.
Sköna täcken gör hon åt sig, hon har kläder av finaste linne och purpur.
Hennes man är känd i stadens portar, där han sitter bland landets äldste.
Fina linneskjortor gör hon och säljer dem, och bälten avyttrar hon till krämaren.
Kraft och heder är hennes klädnad, och hon ler mot den dag som kommer.
Sin mun upplåter hon med vishet, och har vänlig förmaning på sin tunga.
Hon vakar över ordningen i sitt hus och äter ej i lättja sitt bröd.
Hennes söner stå upp och prisa henne säll, hennes man likaså och förkunnar hennes lov:
»Många idoga kvinnor hava funnits, men du, du övergår dem allasammans.»
Skönhet är förgänglig och fägring en vindfläkt; men prisas må en hustru som fruktar HERREN.
Må hon få njuta sina gärningars frukt; hennes verk skola prisa henne i portarna.
Detta är predikarens ord, Davids sons, konungens i Jerusalem.
Fåfängligheters fåfänglighet! säger Predikaren.
Fåfängligheters fåfänglighet!
Allt är fåfänglighet!
Vad förmån har människan av all möda som hon gör sig under solen?
Släkte går, och släkte kommer, och jorden står evinnerligen kvar.
Och solen går upp, och solen går ned, och har sedan åter brått att komma till den ort där hon går upp.
Vinden far mot söder och vänder sig så mot norr; den vänder sig och vänder sig, allt under det att den far fram, och så begynner den åter sitt kretslopp.
Alla floder rinna ut i havet, och ändå bliver havet aldrig fullt; där floderna förut hava runnit, dit rinna de ständigt åter.
Alla arbetar utan rast; ingen kan utsäga det.
Ögat mättas icke av att se, och örat bliver icke fullt av att höra.
Vad som har varit är vad som kommer att vara, och vad som har hänt är vad som kommer att hända; intet nytt sker under solen.
Inträffar något varom man ville säga: »Se, detta är nytt», så har detsamma ändå skett redan förut, i gamla tider, som voro före oss.
Man kommer icke ihåg dem som levde före oss.
Och dem som skola uppstå efter oss skall man icke heller komma ihåg bland dem som leva ännu senare.
Jag, Predikaren, var konung över Israel i Jerusalem.
Och jag vände mitt hjärta till att begrunda och utrannsaka genom vishet allt vad som händer under himmelen; sådant är ett uselt besvär, som Gud har givit människors barn till att plåga sig med.
När jag nu såg på allt vad som händer under himmelen, se, då var det allt fåfänglighet och ett jagande efter vind.
Det som är krokigt kan icke bliva rakt, och det som ej finnes kan ej komma med i någon räkning.
Jag sade i mitt hjärta: »Se, jag har förvärvat mig stor vishet, och jag har förökat den, så att den övergår allas som före mig hava regerat över Jerusalem; ja, vishet och insikt har mitt hjärta inhämtat i rikt mått.»
Men när jag nu vände mitt hjärta till att förstå vishet och till att förstå oförnuft och dårskap, då insåg jag att också detta var ett jagande efter vind.
Ty där mycken vishet är, där är mycken grämelse; och den som förökar sin insikt, han förökar sin plåga.
Jag sade i mitt hjärta: »Välan, jag vill pröva huru glädje kommer dig, gör dig nu goda dagar.»
Men se, också detta var fåfänglighet.
Jag måste säga om löjet: »Det är dårskap», och om glädjen: »Vad gagnar den till?»
I mitt hjärta begrundade jag huru jag skulle pläga min kropp med vin -- allt under det att mitt hjärta ägnade sig åt vishet -- och huru jag skulle hålla fast vid dårskap, till dess jag finge se vad som vore bäst för människors barn att göra under himmelen, de dagar de leva.
Jag företog mig stora arbeten, jag byggde hus åt mig, jag planterade vingårdar åt mig.
Jag anlade åt mig lustgårdar och parker och planterade i dem alla slags fruktträd.
Jag anlade vattendammar åt mig för att ur dem vattna den skog av träd, som växte upp.
Jag köpte trälar och trälinnor, och hemfödda tjänare fostrades åt mig; jag fick ock boskap, fäkreatur och får, i större myckenhet än någon som före mig hade varit i Jerusalem.
Jag samlade mig jämväl silver och guld och allt vad konungar och länder kunna äga; jag skaffade mig sångare och sångerskor och vad som är människors lust: en hustru, ja, många.
Så blev jag stor, allt mer och mer, större än någon som före mig hade varit i Jerusalem; och under detta bevarade jag ändå min vishet.
Intet som mina ögon begärde undanhöll jag dem, och ingen glädje nekade jag mitt hjärta.
Ty mitt hjärta fann glädje i all min möda, och detta var min behållna del av all min möda.
Men när jag så vände mig till att betrakta alla de verk som mina händer hade gjort, och den möda som jag hade nedlagt på dem, se, då var det allt fåfänglighet och ett jagande efter vind.
Ja, under solen finnes intet som kan räknas för vinning.
När jag alltså vände mig till att jämföra vishet med oförnuft och dårskap -- ty vad kunna de människor göra, som komma efter konungen, annat än detsamma som man redan förut har gjort? --
då insåg jag att visheten väl har samma företräde framför dårskapen, som ljuset har framför mörkret:
Den vise har ögon i sitt huvud, men dåren vandrar i mörker.
Dock märkte jag att det går den ene som den andre.
Då sade jag i mitt hjärta: »Såsom det går dåren, så skall det ock gå mig; vad gagn har då därav att jag är förmer i vishet?»
Och jag sade i mitt hjärta att också detta var fåfänglighet.
Ty den vises minne varar icke evinnerligen, lika litet som dårens; i kommande dagar skall ju alltsammans redan vara förgätet.
Och måste icke den vise dö såväl som dåren?
Och jag blev led vid livet, ty illa behagade mig vad som händer under solen, eftersom allt är fåfänglighet och ett jagande efter vind.
Ja, jag blev led vid all den möda som jag hade gjort mig under solen, eftersom jag åt någon annan som skall komma efter mig måste lämna vad jag har gjort.
Och vem vet om denne skall vara en vis man eller en dåre?
Men ändå skall han få råda över allt det varpå jag har nedlagt min möda och min vishet under solen.
Också detta är fåfänglighet.
Så begynte jag då att åter förtvivla i mitt hjärta över all den möda som jag hade gjort mig under solen.
Ty om en människa med vishet och insikt och skicklighet har utstått sin möda, så måste hon dock lämna sin del åt en annan som icke har haft någon möda därmed.
Också detta är fåfänglighet och ett stort elände.
Ja, vad gagn har människan av all möda och hjärteoro som hon gör sig under solen?
Alla hennes dagar äro ju fulla av plåga, och det besvär hon har är fullt av grämelse; icke ens om natten får hennes hjärta någon ro.
Också detta är fåfänglighet.
Det är icke en lycka som beror av människan själv, att hon kan äta och dricka och göra sig goda dagar under sin möda.
Jag insåg att också detta kommer från Guds hand, hans som har sagt:
»Vem kan äta, och vem kan njuta, mig förutan?»
Ty åt den människa som täckes honom giver han vishet och insikt och glädje; men åt syndaren giver han besväret att samla in och lägga tillhopa, för att det sedan må tillfalla någon som täckes Gud.
Också detta är fåfänglighet och ett jagande efter vind.
Allting har sin tid, och vart företag under himmelen har sin stund.
Födas har sin tid, och dö har sin tid.
Plantera har sin tid, och rycka upp det planterade har sin tid.
Dräpa har sin tid, och läka har sin tid.
Bryta ned har sin tid, och bygga upp har sin tid.
Gråta har sin tid, och le har sin tid.
Klaga har sin tid, och dansa har sin tid.
Kasta undan stenar har sin tid, och samla ihop stenar har sin tid.
Taga i famn har sin tid, och avhålla sig från famntag har sin tid.
Söka upp har sin tid, och tappa bort har sin tid.
Förvara har sin tid, och kasta bort har sin tid.
Riva sönder har sin tid, och sy ihop har sin tid.
Tiga har sin tid, och tala har sin tid.
Älska har sin tid, och hata har sin tid.
Krig har sin tid, och fred har sin tid.
Vad förmån av sin möda har då den som arbetar?
Jag såg vilket besvär Gud har givit människors barn till att plåga sig med.
Allt har han gjort skönt för sin tid, ja, han har ock lagt evigheten i människornas hjärtan, dock så, att de icke förmå att till fullo, ifrån begynnelsen intill änden, fatta det verk som Gud har gjort.
Jag insåg att intet är bättre för dem, än att de äro glada och göra sig goda dagar, så länge de leva.
Men om någon kan äta och dricka och njuta vad gott är under all sin möda, så är också detta en Guds gåva.
Jag insåg att allt vad Gud gör skall förbliva evinnerligen; man kan icke lägga något därtill, ej heller taga något därifrån.
Och Gud har så gjort, för att man skall frukta honom.
Vad som är, det var redan förut, och vad som kommer att ske, det skedde ock redan förut; Gud söker blott fram det förgångna.
Ytterligare såg jag under solen att på domarsätet rådde orättfärdighet, och på rättfärdighetens säte orättfärdighet.
Då sade jag i mitt hjärta: Både den rättfärdige och den orättfärdige skall Gud döma; ty vart företag och allt vad man gör har sin tid hos honom.
Jag sade i mitt hjärta: För människornas skull sker detta, på det att Gud må pröva dem, och på det att de själva må inse att de äro såsom fänad.
Ty det går människors barn såsom det går fänaden, dem alla går det lika.
Såsom fänaden dör, så dö ock de; enahanda ande hava de ock alla.
Ja, människorna hava intet framför fänaden, ty allt är fåfänglighet.
Alla går de till samma mål; alla have de kommit av stoft, och alla skola de åter varda stoft.
Vem kan veta om människornas ande att den stiger uppåt, och om fänadens ande att den far ned under jorden?
Och jag såg att intet är bättre för människan, än att hon är glad under sitt arbete; ty detta är den del hon får.
Ty vem kan föra henne tillbaka, så att hon får se och hava glädje av vad som skall ske efter henne?
Och ytterligare såg jag på alla de våldsgärningar som förövas under solen.
Jag såg förtryckta fälla tårar, och ingen fanns, som tröstade dem; jag såg dem lida övervåld av sina förtryckares hand, och ingen fanns, som tröstade dem.
Då prisade jag de döda, som redan hade fått dö, lyckliga framför de levande, som ännu leva;
Men lycklig framför båda prisade jag den som ännu icke hade kommit till, den som hade sluppit att se vad ont som göres under solen.
Och jag såg att all möda och all skicklighet i vad som göres icke är annat än den enes avund mot den andre.
Också detta är fåfänglighet och ett jagande efter vind.
Dåren lägger händerna i kors och tär så sitt eget kött.
Ja, bättre är en handfull ro än båda händerna fulla med möda och med jagande efter vind.
Och ytterligare såg jag något som är fåfänglighet under solen:
mången finnes, som står ensam och icke har någon jämte sig, varken son eller broder; och likväl är det ingen ände på all hans möda, och hans ögon bliva icke mätta på rikedom.
Och för vem mödar jag mig då och nekar mig själv vad gott är?
Också detta är fåfänglighet och ett uselt besvär.
Bättre är att vara två än en, ty de två få större vinning av sin möda.
Om någondera faller, så kan ju den andre resa upp sin medbroder.
Men ve den ensamme, om han faller och icke en annan finnes, som kan resa upp honom.
Likaledes, om två ligga tillsammans, så hava de det varmt; men huru skall den ensamme bliva varm?
Och om någon kan slå ned den som är ensam, så hålla dock två stånd mot angriparen.
Och en tretvinnad tråd brister icke så snart.
Bättre är en gammal konung som är dåraktig och ej har förstånd nog att låta varna sig är en fattig yngling med vishet.
Ty ifrån fängelset gick en gång en sådan till konungavälde, fastän han var född i fattigdom inom den andres rike.
Jag såg huru alla som levde och rörde sig under solen följde ynglingen, denne nye som skulle träda i den förres ställe;
det var ingen ände på hela skaran av alla dem som han gick i spetsen för.
Men ändå hava de efterkommande ingen glädje av honom.
Ty också detta är fåfänglighet och ett jagande efter vind.
Bevara din fot, när du går till Guds hus; att komma dit för att höra är bättre än något slaktoffer som dårarna frambära; ty de äro oförståndiga och göra så vad ont är.
Var icke obetänksam med din mun, och låt icke ditt hjärta förhasta sig med att uttala något ord inför Gud.
Gud är ju i himmelen, och du är på jorden; låt därför dina ord vara få.
Ty tanklöshet har med sig mångahanda besvär, och en dåres röst har överflöd på ord.
När du har gjort ett löfte åt Gud, så dröj icke att infria det; ty till dårar har han icke behag.
Det löfte du har givit skall du infria.
Det är bättre att du intet lovar, än att du gör ett löfte och icke infriar det.
Låt icke din mun draga skuld över hela din kropp; och säg icke inför Guds sändebud att det var ett förhastande.
Icke vill du att Gud skall förtörnas för ditt tals skull, så att han fördärvar sina händers verk?
Se, där mycken tanklöshet och fåfänglighet är, där är ock en myckenhet av ord.
Ja, Gud må du frukta.
Om du ser att den fattige förtryckes, och att rätt och rättfärdighet våldföres i landet, så förundra dig icke däröver; ty på den höge vaktar en högre, och andra ännu högre vakta på dem båda.
Och vid allt detta är det en förmån för ett land att hava en konung som så styr, att marken bliver brukad.
Den som så älskar penningar bliver icke mätt på penningar, och den som älskar rikedom har ingen vinning därav.
Också detta är fåfänglighet.
När ägodelarna förökas, bliva ock de som äta av dem många; och till vad gagn äro de då för ägaren, utom att hans ögon få se dem?
Söt är arbetarens sömn, vare sig han har litet eller mycket att äta; men den rikes överflöd tillstädjer honom icke att sova.
Ett bedrövligt elände som jag har sett under solen är det att hopsparad rikedom kan bliva sin ägare till skada.
Och om rikedomen har gått förlorad för någon genom en olycka, så får hans son, om han har fött en son, alls intet därav.
Sådan som han kom ur sin moders liv måste han själv åter gå bort, lika naken som han kom, och för sin möda får han alls intet som han kan taga med sig.
Också det är ett bedrövligt elände.
Om han måste gå bort alldeles sådan som han kom, vad förmån har han då därav att han så mödar sig -- för vind?
Nej, alla sina livsdagar framlever han i mörker; och mycken grämelse har han, och plåga och förtret.
Se, vad jag har funnit vara bäst och skönast för människan, det är att hon äter och dricker och gör sig goda dagar vid den möda som hon har under solen, medan de livsdagar vara, som Gud giver henne; ty detta är den del hon får.
Och om Gud åt någon har givit rikedom och skatter, och därtill förunnat honom makt att njuta härav och att göra sig till godo sin del och att vara glad under sin möda, så är också detta en Guds gåva.
Ty man tänker då icke så mycket på sina livsdagars gång, när Gud förlänar glädje i hjärtat.
Ett elände som jag har sett under solen, och som kommer tungt över människorna är det,
när Gud åt någon har givit rikedom och skatter och ära, så att denne för sin räkning intet saknar av allt det han önskar sig, och Gud sedan icke förunnar honom makt att själv njuta därav, utan låter en främling få njuta därav; detta är fåfänglighet och en usel plåga.
Om en man än finge hundra barn och finge leva i många år, ja, om hans livsdagar bleve än så många, men hans själ icke finge njuta sig mätt av hans goda, och om han så bleve utan begravning, då säger jag: lyckligare än han är ett ofullgånget foster.
Ty såsom ett fåfängligt ting har detta kommit till världen, och i mörker går det bort, och i mörker höljes dess namn;
det fick ej ens se solen, och det vet av intet.
Ett sådant har bättre ro än han.
Ja, om han än levde i två gånger tusen år utan att få njuta något gott -- gå icke ändå alla till samma mål?
All människans möda är för hennes mun, och likväl bliver hennes hunger icke mättad.
Ty vad förmån har den vise framför dåren?
Vad båtar det den fattige, om han förstår att skicka sig inför de levande?
Bättre är att se något för ögonen än att fara efter något med begäret.
Också detta är fåfänglighet och ett jagande efter vind.
Vad som är, det var redan förut nämnt vid namn; förutbestämt var vad en människa skulle bliva.
Och hon kan icke gå till rätta med honom som är mäktigare än hon själv.
Ty om man ock ordar än så mycket och därmed förökar fåfängligheten, vad förmån har man därav?
Ty vem vet vad gott som skall hända en människa i livet, under de fåfängliga livsdagar som hon får framleva, lik en skugga?
Och vem kan säga en människa vad som efter henne skall ske under solen?
Bättre är gott namn än god salva, och bättre är dödens dag än födelsedagen.
Bättre än att gå i gästabudshus är det att gå i sorgehus; ty där är änden för alla människor, och den efterlevande må lägga det på hjärtat.
Bättre är grämelse än löje, ty av det som gör ansiktet sorgset far hjärtat väl.
De visas hjärtan äro i sorgehus, och dårarnas hjärtan i hus där man glädes.
Bättre är att höra förebråelser av en vis man än att få höra sång av dårar.
Ty såsom sprakandet av törne under grytan, så är dårarnas löje.
Också detta är fåfänglighet.
Ty vinningslystnad gör den vise till en dåre, och mutor fördärva hjärtat.
Bättre är slutet på en sak än dess begynnelse; bättre är en tålmodig man än en högmodig.
Var icke för hastig i ditt sinne till att gräma dig, ty grämelse bor i dårars bröst.
Spörj icke: »Varav kommer det att forna dagar voro bättre än våra?»
Ty icke av vishet kan du fråga så.
Jämgod med arvgods är vishet, ja, hon är förmer i värde för dom som se solen.
Ty under vishetens beskärm är man såsom under penningens beskärm, men den förståndiges förmån är att visheten behåller sin ägare vid liv.
Se på Guds verk; vem kan göra rakt vad han har gjort krokigt?
Var alltså vid gott mod under den goda dagen, och betänk under den onda dagen att Gud har gjort denna såväl som den andra, för att människan icke skall kunna utfinna något om det som skall ske, när hon är borta.
Det ena som det andra har jag sett under mina fåfängliga dagar: mången rättfärdig som har förgåtts i sin rättfärdighet, och mången orättfärdig som länge har fått leva i sin ondska.
Var icke alltför rättfärdighet, och var icke alltför mycket vis; icke vill du fördärva dig själv?
Var icke alltför orättfärdig, och var icke en dåre; icke vill du dö i förtid?
Det är bäst att du håller fast vid det ena, utan att ändå släppa det andra; ty den som fruktar Gud finner en utväg ur allt detta.
Visheten gör den vise starkare än tio väldiga i staden.
Ty ingen människa är så rättfärdig på jorden, att hon gör vad gott är och icke begår någon synd.
Akta icke heller på alla ord som man talar, eljest kunde du få höra din egen tjänare uttala förbannelser över dig.
Ditt hjärta vet ju att du själv mången gång har uttalat förbannelser över andra.
Detta allt har jag försökt att utröna genom vishet.
Jag sade: »Jag vill bliva vis», men visheten förblev fjärran ifrån mig.
Ja, tingens väsen ligger i fjärran, djupt nere i djupet; vem kan utgrunda det?
När jag vände mig med mitt hjärta till att eftersinna och begrunda, och till att söka visheten och det som är huvudsumman, och till att förstå ogudaktigheten i dess dårskap och dåraktigheten i dess oförnuft,
då fann jag något som var bittrare än döden: kvinnan, hon som själv är ett nät, och har ett hjärta som är en snara, och armar som äro bojor.
Den som täckes Gud kan undkomma henne, men syndaren bliver hennes fånge.
Se, detta fann jag, säger Predikaren, i det jag lade det ena till det andra för att komma till huvudsumman.
Något gives, som min själ beständigt har sökt, men som jag icke har funnit: väl har jag funnit en man bland tusen, men en kvinna har jag icke funnit i hela hopen.
Dock se, detta har jag funnit, att Gud har gjort människorna sådana de borde vara, men själva tänka de ut mångahanda funder.
Vem är lik den vise, och vem förstår att så uttyda en sak?
Visheten gör människans ansikte ljust, genom den förvandlas det råa i hennes uppsyn.
Jag säger er: Akta på konungens bud, ja, gör det för den eds skull som du har svurit vid Gud.
Förhasta dig icke att övergiva honom, inlåt dig ej på något som är ont; han kan ju göra allt vad han vill.
Ty en konungs ord är mäktigt, och vem kan säga till honom: »Vad gör du?»
Den som håller budet skall icke veta av något ont; och tid och sätt skall den vises hjärta lära känna.
Ty vart företag har sin tid och sitt sätt, och en människas ondska kommer tungt över henne.
Hon vet ju icke vad som kommer att ske; vem kan säga henne huru något kommer att ske?
Ingen människa har makt över vinden, till att hejda den, ej heller har någon makt över dödens dag, ej heller finnes undflykt i krig; så kan ogudaktigheten icke rädda sin man.
Allt detta såg jag, när jag gav akt på allt vad som händer under solen, i en tid då den ena människan har makt över den andra, henne till olycka.
Ock likaledes såg jag att de ogudaktiga fingo komma i sin grav och gå till vila, under det att sådana som hade gjort vad rätt var måste draga bort ifrån den Heliges boning och blevo förgätna i staden.
Också detta är fåfänglighet.
Därför att dom icke strax går över vad ont som göres, få människors barn dristighet att göra det ont är,
eftersom syndaren hundra gånger kan göra vad ont är och likväl får länge leva.
Dock vet jag ju att det skall gå de gudfruktiga väl, därför att de frukta Gud,
men att det icke skall gå den ogudaktige väl, och att hans dagar icke skola förlängas, såsom skuggan förlänges, eftersom han icke fruktar Gud.
En fåfänglighet som händer här på jorden är det att rättfärdiga finnas, vilka det går såsom hade de gjort de ogudaktigas gärningar, och att ogudaktiga finnas, vilka det går såsom hade de gjort de rättfärdigas gärningar.
Jag sade: Också detta är fåfänglighet.
Så prisade jag då glädjen och fann att intet är bättre för människan under solen, än att hon äter ock dricker och är glad, så att detta får följa henne vid hennes möda, under de livsdagar som Gud giver henne under solen.
När jag vände mitt hjärta till att förstå vishet, och till att betrakta det besvär som man gör sig på jorden utan att få sömn i sina ögon, varken dag eller natt,
då insåg jag att det är så med alla Guds verk, att människan icke förmår fatta vad som händer under solen; ty huru mycket en människa än mödar sig för att utforska det, fattar hon det ändå icke.
Och om någon vis man tänker att han skall kunna förstå det, så kommer han ändå icke att kunna fatta det.
Ja, allt detta har jag besinnat, och jag har sökt pröva allt detta, huru de rättfärdiga och de visa och deras verk äro i Guds våld.
Varken om kärlek eller hat kan en människa veta något förut; allt kan förestå henne.
Ja, allt kan vederfaras alla; det går den rättfärdige såsom den ogudaktige, den gode och rene såsom den orene, den som offrar såsom den vilken icke offrar; den gode räknas lika med syndaren, den som svär bliver lik den som har försyn för att svärja.
Ett elände vid allt som händer under solen är detta, att det går alla lika.
Därför äro ock människornas hjärtan fulla med ondska, och oförnuft är i deras hjärtan, så länge de leva; och sedan måste de ned bland de döda.
För den som utkoras att vara i de levandes skara finnes ju ännu något att hoppas; ty bättre är att vara en levande hund än ett dött lejon.
Och väl veta de som leva att de måste dö, men de döda vet alls intet, och de hava ingen vinning mer att vänta, utan deras åminnelse är förgäten.
Både deras kärlek och deras hat och deras avund hava redan nått sin ände, och aldrig någonsin få de mer någon del i vad som händer under solen.
Välan, så ät då ditt bröd med glädje, och drick ditt vin med glatt hjärta, ty Gud har redan i förväg givit sitt bifall till vad du gör.
Låt dina kläder alltid vara vita, och låt aldrig olja fattas på ditt huvud.
Njut livet med någon kvinna som du älskar, så länge de fåfängliga livsdagar vara, som förlänas dig under solen, ja, under alla dina fåfängliga dagar; ty detta är den del du får i livet vid den möda som du gör dig under solen.
Allt vad du förmår uträtta med din kraft må du söka uträtta; ty i dödsriket, dit du går, kan man icke verka eller tänka, där finnes ingen insikt eller vishet.
Ytterligare såg jag under solen att det icke beror av de snabba huru de lyckas i löpandet, icke av hjältarna huru striden utfaller, icke av de visa huru de få sitt bröd, icke av de kloka vad rikedom de förvärva, eller av de förståndiga vad ynnest de vinna, utan att allt för dem beror av tid och lägenhet.
Ty människan känner icke sin tid, lika litet som fiskarna, vilka fångas i olycksnätet, eller fåglarna, vilka fastna i snaran.
Såsom dessa, så snärjas ock människornas barn på olyckans tid, när ofärd plötsligt faller över dem.
Också detta såg jag under solen, ett visdomsverk, som tycktes mig stort:
Det fanns en liten stad med få invånare, och mot den kom en stor konung och belägrade den och byggde stora bålverk mot den.
Men därinne fanns en fattig man som var vis; och denne räddade staden genom sin vishet.
Dock, sedan tänkte ingen människa på denne fattige man.
Då sade jag: Väl är vishet bättre än styrka, men den fattiges vishet bliver icke föraktad, och hans ord varda icke hörda.
De vises ord, om de ock höras helt stilla, äro förmer än allt ropande av en dårarnas överste.
Bättre är vishet än krigsredskap; ty en enda som felar kan fördärva mycket gott.
Giftflugor vålla stank och jäsning i salvoberedarens salva; så uppväger ett grand av dårskap både vishet och ära.
Den vise har sitt hjärta åt höger, men dåren har sitt hjärta åt vänster.
Ja, varhelst dåren går kommer hans förstånd till korta, och till alla säger han ifrån, att han är en dåre.
Om hos en furste vrede uppstår mot dig, så håll dig dock stilla, ty saktmod gör stora synder ogjorda.
Ett elände gives, som jag har sett under solen, ett fel som beror av den som har makten:
att dårskap sättes på höga platser, medan förnämliga män få sitta i förnedring.
Jag har sett trälar färdas till häst och hövdingar få gå till fots såsom trälar.
Den som gräver en grop, han faller själv däri, och den som bryter ned en mur, honom stinger ormen.
Den som vältrar bort stenar bliver skadad av dem, den som hugger ved kommer i fara därvid.
Om man icke slipar eggen, när ett järn har blivit slött, så måste man anstränga krafterna dess mer; och vishet är att göra allt på bästa sätt.
Om ormen får stinga, innan han har blivit tjusad, så har besvärjaren intet gagn av sin konst.
Med sin muns ord förvärvar den vise ynnest, men dårens läppar fördärva honom själv.
Begynnelsen på hans muns ord är dårskap, och änden på hans tal är uselt oförnuft.
Och dåren är rik på ord; dock vet ingen människa vad som skall ske; vem kan säga en människa vad som efter henne skall ske?
Dårens möda bliver honom tung, ty icke ens till staden hittar han fram.
Ve dig, du land vars konung är ett barn, och vars furstar hålla måltid redan på morgonen!
Väl dig, du land vars konung är en ädling, och vars furstar hålla måltid i tillbörlig tid, med måttlighet, och icke för att överlasta sig!
Genom lättja förfalla husets bjälkar, och genom försumlighet dryper det in i huset.
Till sin förlustelse håller man gästabud, och vinet gör livet glatt; men penningen är det som förlänar alltsammans.
Uttala ej ens i din tanke förbannelser över en konung, och ej ens i din sovkammare förbannelser över en rik man; ty himmelens fåglar böra fram ditt tal, och de bevingade förkunna vad du har sagt.
Sänd ditt bröd över vattnet, ty i tidens längd får du det tillbaka.
Dela vad du har i sju delar, ja, i åtta, ty du vet icke vilken olycka som kan gå över landet.
Om molnen äro fulla av regn, så tömma de ut det på jorden; och om ett träd faller omkull, det må falla mot söder eller mot norr, så ligger det på den plats där det har fallit.
En vindspejare får aldrig så, och en molnspanare får aldrig skörda.
Lika litet som du vet vart vinden far, eller huru benen bildas i den havandes liv, lika litet förstår du Guds verk, hans som verkar alltsammans.
Så ut om morgonen din säd, och underlåt det ej heller om aftonen, ty du vet icke vilketdera som är gagneligast, eller om det ena jämte det andra är bäst.
Och ljuset är ljuvligt, och det är gott för ögonen att få se solen.
Ja, om en människa får leva än så många år, så må hon vara glad under dem alla, men betänka, att eftersom mörkrets dagar bliva så många, är ändå allt som händer fåfänglighet.
Gläd dig, du yngling, din ungdom, och låt ditt hjärta unna dig fröjd i din ungdomstid; ja, vandra de vägar ditt hjärta lyster och så, som det behagar dina ögon.
Men vet att Gud för allt detta skall draga dig till doms.
Ja, låt grämelse vika ur ditt hjärta, och håll plåga borta från din kropp.
Ty ungdom och blomstring är fåfänglighet.
Så tänk då på din Skapare i din ungdomstid, förrän de onda dagarna komma och de år nalkas, om vilka du skall säga: »Jag finner icke behag i dem»;
Ja, förrän solen bliver förmörkad, och dagsljuset och månen och stjärnorna; före den ålder då molnen komma igen efter regnet,
den tid då väktarna i huset darra och de starka männen kröka sig; då malerskorna sitta fåfänga, så få som de nu hava blivit, och skåderskorna hava det mörkt i sina fönster;
då dörrarna åt gatan stängas till, medan ljudet från kvarnen försvagas; då man står upp, när fågeln begynner kvittra, och alla sångens tärnor sänka rösten;
då man fruktar för var backe och förskräckelser bo på vägarna; då mandelträdet blommar och gräshoppan släpar sig fram och kaprisknoppen bliver utan kraft, nu då människan skall fara till sin eviga boning och gråtarna redan gå och vänta på gatan;
ja, förrän silversnöret ryckes bort och den gyllene skålen slås sönder, och förrän ämbaret vid källan krossas och hjulet slås sönder och faller i brunnen
och stoftet vänder åter till jorden, varifrån det har kommit, och anden vänder åter till Gud, som har givit den.
Fåfängligheters fåfänglighet! säger Predikaren.
Allt är fåfänglighet! ----
För övrigt är att säga att Predikaren var en vis man, som också annars lärde folket insikt och övervägde och rannsakade; många ordspråk författade han.
Predikaren sökte efter att finna välbehagliga ord, sådant som med rätt kunde skrivas, och sådant som med sanning kunde sägas.
De visas ord äro såsom uddar, och lika indrivna spikar äro deras tänkespråk.
De äro gåvor från en och samma Herde.
Och för övrigt är utom detta att säga: Min son, låt varna dig!
Ingen ände är på det myckna bokskrivandet, och mycket studerande gör kroppen trött.
Änden på talet, om vi vilja höra huvudsumman, är detta: Frukta Gud och håll hans bud, ty det hör alla människor till.
Ty Gud skall draga alla gärningar till doms, när han dömer allt vad förborgat är, evad det är gott eller ont.
Sångernas sång av Salomo.
Kyssar give han mig, kyssar av sin mun!
Ty din kärlek är mer ljuv än vin.
Ljuv är doften av dina salvor, ja, en utgjuten salva är ditt namn; fördenskull hava tärnorna dig kär.
Drag mig med dig!
Med hast vilja vi följa dig.
Ja, konungen har fört mig in i sina gemak; Vi vilja fröjdas och vara glada över dig, vi vilja prisa din kärlek högre än vin; med rätta har man dig kär. ----
Svart är jag, dock är jag täck, I Jerusalems döttrar, lik Kedars hyddor, lik Salomos tält.
Sen icke därpå att jag är så svart, att solen har bränt mig så.
Min moders söner blevo vreda på mig och satte mig till vingårdsvakterska; min egen vingård kunde jag icke vakta.
»Säg mig, du som min själ har kär: Var för du din hjord i bet?
Var låter du den vila om middagen?
Må jag slippa att gå lik en vilsekommen kvinna vid dina vänners hjordar.»
»Om du icke vet det, du skönaste bland kvinnor, så gå blott åstad i hjordens spår, och för dina killingar i bet vid herdarnas tält.» ----
»Vid ett sto i Faraos spann förliknar jag dig, min älskade.
Dina kinder äro så täcka med sina kedjehängen, din hals med sina pärlerader.
Kedjehängen av guld vilja vi skaffa åt dig med silverkulor på.»
»Medan konungen håller sin fest, sprider min nardus sin doft.
Min vän är för mig ett myrragömme, som jag bär i min barm.
Min vän är för mig en klase cyperblommor från En-Gedis vingårdar.»
»Vad du är skön, min älskade!
Vad du är skön!
Dina ögon äro duvor.»
»Vad du är skön, min vän!
Ja, ljuvlig är du, och grönskande är vårt viloläger.
Bjälkarna i vår boning äro cedrar, och cypresser vår väggpanel.»
»Jag är ett ringa blomster i Saron, en lilja i dalen.»
»Ja, såsom en lilja bland törnen, så är min älskade bland jungfrur.»
»Såsom ett äppelträd bland vildmarkens träd, så är min vän bland ynglingar; ljuvligt är mig att sitta i dess skugga, och söt är dess frukt för min mun.
I vinsalen har han fört mig in, och kärleken är hans baner över mig.
Vederkvicken mig med druvkakor, styrken mig med äpplen; ty jag är sjuk av kärlek.» ----
Hans vänstra arm vilar under mitt huvud, och hans högra omfamnar mig.
Jag besvär eder, I Jerusalems döttrar, vid gaseller och hindar på marken: Oroen icke kärleken, stören den icke, förrän den själv så vill. ----
Hör, där är min vän!
Ja, där kommer han, springande över bergen, hoppande fram på höjderna.
Lik en gasell är min vän eller lik en ung hjort.
Se, nu står han där bakom vår vägg, han blickar in genom fönstret, han skådar genom gallret.
Min vän begynner tala, han säger till mig: »Stå upp, min älskade, du min sköna, och kom hitut.
Ty se, vintern är förbi, regntiden är förliden och har gått sin kos.
Blommorna visa sig på marken, tiden har kommit, då vinträden skäras, och turturduvan låter höra sin röst i vårt land.
Fikonträdets frukter begynna att mogna, vinträden stå redan i blom, de sprida sin doft.
Stå upp, min älskade, min sköna, och kom hitut.
Du min duva i bergsklyftan, i klippväggens gömsle, låt mig se ditt ansikte, låt mig höra din röst; ty din röst är så ljuv, och ditt ansikte är så täckt.» ----
Fången rävarna åt oss, de små rävarna, vingårdarnas fördärvare, nu då våra vingårdar stå i blom. ----
Min vän är min, och jag är hans, där han för sin hjord i bet ibland liljor.
Till dess morgonvinden blåser och skuggorna fly, må du ströva omkring, lik en gasell, min vän, eller lik en ung hjort, på de kassiadoftande bergen.
5. -- Brudtåget beskrives v.
6--11.
Där jag låg på mitt läger om natten, sökte jag honom som min själ har kär; jag sökte honom, men fann honom icke.
»Jag vill stå upp och gå omkring i staden, på gatorna och på torgen; jag vill söka honom som min själ har kär.»
Jag sökte honom, men fann honom icke.
Väktarna mötte mig, där de gingo omkring i staden. »Haven I sett honom som min själ har kär?»
Knappt hade jag kommit förbi dem, så fann jag honom som min själ har kär.
Jag tog honom fatt, och jag släppte honom icke, förrän jag hade fört honom in i min moders hus, in i min fostrarinnas kammare. ----
Jag besvär eder, I Jerusalems döttrar, vid gaseller och hindar på marken: Oroen icke kärleken, stören den icke, förrän den själv så vill. ----
Vem är hon som kommer hitupp från öknen såsom i stoder av rök, kringdoftad av myrra och rökelse och alla slags köpmannakryddor?
Se, det är Salomos bärstol!
Sextio hjältar omgiva den, utvalda bland Israels hjältar.
Alla bära de svärd och äro väl förfarna i strid.
Var och en har sitt svärd vid sin länd, till värn mot nattens faror.
En praktbår är det som konung Salomo har låtit göra åt sig av virke från Libanon.
Dess sidostöd äro gjorda av silver, ryggstödet av guld, sätet belagt med purpurrött tyg.
Innantill är den prydd i kärlek av Jerusalems döttrar.
I Sions döttrar, gån ut och skåden konung Salomo med lust, skåden kransen som hans moder har krönt honom med på hans bröllopsdag, på hans hjärtefröjds dag.
Vad du är skön, min älskade, vad du är skön!
Dina ögon äro duvor, där de skymta genom din slöja.
Ditt hår är likt en hjord av getter som strömma nedför Gileads berg.
Dina tänder likna en hjord av nyklippta tackor, nyss uppkomna ur badet, allasammans med tvillingar, ofruktsam är ingen ibland dem.
Ett rosenrött snöre likna dina läppar, och täck är din mun.
Lik ett brustet granatäpple är din kind, där den skymtar genom din slöja.
Din hals är lik Davids torn, det väl befästa; tusen sköldar hänga därpå, hjältarnas alla sköldar.
Din barm är lik ett killingpar, tvillingar av en gasell, som gå i bet ibland liljor.
Till dess morgonvinden blåser och skuggorna fly, vill jag gå bort till myrraberget, till den rökelsedoftande höjden.
Du är skön alltigenom, min älskade, på dig finnes ingen fläck. ----
Kom med mig från Libanon, min brud, kom med mig från Libanon.
Stig ned från Amanas topp, från toppen av Senir och Hermon, från lejonens hemvist, från pantrarnas berg. ----
Du har tagit mitt hjärta, du min syster, min brud; du har tagit mitt hjärta med en enda blick, med en enda länk av kedjan kring din hals.
Huru skön är icke din kärlek, du min syster, min brud!
Huru ljuv är icke din kärlek!
Ja, mer ljuv än vin; och doften av dina salvor övergår all vällukt.
Av sötma drypa dina läppar, min brud; din tunga gömmer honung och mjölk, och doften av dina kläder är såsom Libanons doft. ----
»En tillsluten lustgård är min syster, min brud, en tillsluten brunn, en förseglad källa.
Såsom en park av granatträd skjuter du upp, med de ädlaste frukter, med cyperblommor och nardusplantor,
med nardus och saffran, kalmus och kanel och rökelseträd av alla slag, med myrra och aloe och de yppersta kryddor av alla slag.
Ja, en källa i lustgården är du, en brunn med friskt vatten och ett rinnande flöde ifrån Libanon.»
»Vakna upp, du nordanvind, och kom, du sunnanvind; blås genom min lustgård, låt dess vällukt strömma ut.
Må min vän komma till sin lustgård och äta dess ädla frukter.»
»Ja, jag kommer till min lustgård, du min syster, min brud; jag hämtar min myrra och mina välluktande kryddor, jag äter min honungskaka och min honung, jag dricker mitt vin och min mjölk.» ---- Äten, I kära, och dricken, ja, berusen eder av kärlek.
Jag låg och sov, dock vakade mitt hjärta.
Hör, då klappar min vän på dörren: »Öppna för mig, du min syster, min älskade, min duva, min fromma; ty mitt huvud är fullt av dagg, mina lockar av nattens droppar.»
»Jag har lagt av mina kläder; skulle jag nu åter taga dem på mig?
Jag har tvagit mina fötter; skulle jag nu orena dem?»
Min vän räckte in sin hand genom luckan; då rördes mitt hjärta över honom.
Jag stod upp för att öppna för min vän, och mina händer dröpo av myrra, mina fingrar av flytande myrra, som fuktade rigelns handtag.
Så öppnade jag för min vän, men min vän var borta och försvunnen.
Min själ blev utom sig vid tanken på hans ord.
Jag sökte honom, men fann honom icke; jag ropade på honom, men han svarade mig icke.
Väktarna mötte mig, där de gingo omkring i staden, de slogo mig, de sårade mig; de ryckte av mig min mantel, väktarna på murarna.
»Jag besvär eder, I Jerusalems döttrar, om I finnen min vän, så sägen -- ja, vad skolen I säga honom?
Att jag är sjuk av kärlek!»
»Vad är då din vän förmer än andra vänner, du skönaste bland kvinnor?
Vad är din vän förmer än andra vänner, eftersom du så besvär oss?»
»Min vän är strålande vit och röd, härlig framför tio tusen.
Hans huvud är finaste guld, hans lockar palmträdsvippor, och svarta såsom korpen.
Hans ögon likna duvor invid vattenbäckar, duvor som bada sig i mjölk och sitta invid bräddfull rand.
Hans kinder liknar välluktrika blomstersängar, skrin med doftande kryddor.
Hans läppar äro röda liljor; de drypa av flytande myrra.
Hans händer äro tenar av guld, besatta med krysoliter.
Hans midja är formad av elfenben, övertäckt med safirer.
Hans ben äro pelare av vitaste marmor, som vila på fotstycken av finaste guld.
Att se honom är såsom att se Libanon; ståtlig är han såsom en ceder.
Hans mun är idel sötma, hela hans väsende är ljuvlighet.
Sådan är min vän, ja, sådan är min älskade, I Jerusalems döttrar.»
»Vart har han då gått, din vän, du skönaste bland kvinnor?
Vart har din vän tagit vägen?
Låt oss hjälpa dig att söka honom.»
»Min vän har gått ned till sin lustgård, till sina välluktrika blomstersängar, för att låta sin hjord beta i lustgårdarna och för att plocka liljor.
Jag är min väns, och min vän är min, där han för sin hjord i bet ibland liljor.
Du är skön såsom Tirsa, min älskade, ljuvlig såsom Jerusalem, överväldigande såsom en härskara.
Vänd bort ifrån mig dina ögon, ty de hava underkuvat mig.
Ditt hår är likt en hjord av getter som strömma nedför Gilead.
Dina tänder likna en hjord av tackor, nyss uppkomna ur badet, allasammans med tvillingar, ofruktsam är ingen ibland dem.
Lik ett brustet granatäpple är din kind, där den skymtar genom din slöja. ----
Sextio äro drottningarna, och åttio bihustrurna, och tärnorna en otalig skara.
Men en enda är hon, min duva, min fromma, hon, sin moders endaste, hon, sin fostrarinnas utkorade.
När jungfrur se henne, prisa de henne säll, drottningar och bihustrur höja hennes lov. ----
Vem är hon som där blickar fram lik en morgonrodnad, skön såsom månen, strålande såsom solen, överväldigande såsom en härskara?
Till valnötslunden gick jag ned, för att glädja mig åt grönskan i dalen, för att se om vinträden hade slagit ut, om granatträden hade fått blommor.
Oförtänkt satte mig då min kärlek upp på mitt furstefolks vagnar.
»Vänd om, vänd om, du brud från Sulem, vänd om, vänd om, så att vi få se på dig.» »Vad finnen I att se hos bruden från Sulem, där hon rör sig såsom i vapendans?»
»Huru sköna äro icke dina fötter i sina skor, du ädla!
Dina höfters rundning är såsom ett bröstspännes kupor, gjorda av en konstnärs händer.
Ditt sköte är en rundad skål, må vinet aldrig fattas däri.
Din midja är en vetehög, omhägnad av liljor.
Din barm är lik ett killingpar, tvillingar av en gasell.
Din hals liknar Elfenbenstornet, dina ögon dammarna i Hesbon, vid Bat-Rabbimsporten.
Din näsa är såsom Libanonstornet, som skådar ut mot Damaskus.
Ditt huvud höjer sig såsom Karmel, och lockarna på ditt huvud hava purpurglans.
En konung är fångad i deras snara.» ----
»Huru skön och huru ljuv är du icke, du kärlek, så följd av lust!
Ja, din växt är såsom ett palmträds, och din barm liknar fruktklasar.
Jag tänker: I det palmträdet vill jag stiga upp, jag vill gripa tag i dess kvistar.
Må din barm då vara mig såsom vinträdets klasar och doften av din andedräkt såsom äpplens doft
och din mun såsom ljuvaste vin!» »Ja, ett vin som lätt glider ned i min vän och fuktar de slumrandes läppar.
Jag är min väns, och till mig står hans åtrå.» ----
Kom, min vän; låt oss gå ut på landsbygden och stanna i byarna över natten.
Bittida må vi gå till vingårdarna, för att se om vinträden hava slagit ut, om knopparna hava öppnat sig, om granatträden hava fått blommor.
Där vill jag giva min kärlek åt dig.
Kärleksäpplena sprida sin doft, och vid våra dörrar finnas alla slags ädla frukter, både nya och gamla; åt dig, min vän, har jag förvarat dem.
Ack att du vore såsom en min broder, ammad vid min moders bröst!
Om jag då mötte dig därute, så finge jag kyssa dig, och ingen skulle tänka illa om mig därför.
Jag finge då ledsaga dig, föra dig in i min moders hus, och du skulle undervisa mig; kryddat vin skulle jag giva dig att dricka, saft från mitt granatträd. ----
Hans vänstra arm vilar under mitt huvud, och hans högra omfamnar mig.
Jag besvär eder, I Jerusalems döttrar: Oroen icke kärleken, stören den icke, förrän den själv så vill.
Vem är hon som kommer hitupp från öknen, stödd på sin vän? »Där under äppelträdet väckte jag dig; där var det som din moder hade fött dig, där födde dig hon som gav dig livet.
Hav mig såsom en signetring vid ditt hjärta, såsom en signetring på din arm.
Ty kärleken är stark såsom döden, dess trängtan obetvinglig såsom dödsriket; dess glöd är såsom eldens glöd, en HERRENS låga är den.
De största vatten förmå ej utsläcka kärleken, strömmar kunna icke fördränka den.
Om någon ville giva alla ägodelar i sitt hus för kärleken, så skulle han ändå bliva försmådd.» ----
»Vi hava en syster, en helt ung, som ännu icke har någon barm.
Vad skola vi göra med vår syster, när tiden kommer, att man vill vinna henne?»
»Är hon en mur, så bygga vi på den ett krön av silver; men är hon en dörr, så bomma vi för den med en cederplanka.»
»Jag är en mur, och min barm är såsom tornen därpå; så blev jag i hans ögon en kvinna som var ynnest värd.» ----
En vingård ägde Salomo i Baal-Hamon, den vingården lämnade han åt väktare; tusen siklar silver var kunde de hämta ur dess frukt.
Men min vingård, den har jag själv i min vård.
Du, Salomo, må taga dina tusen, och två hundra må de få, som vakta dess frukt. ----
»Du lustgårdarnas inbyggerska, vännerna lyssna efter din röst; låt mig höra den.»
»Skynda åstad, min vän, lik en gasell eller lik en ung hjort, upp på de välluktrika bergen.»
Detta är Jesajas, Amos' sons, syner, vad han skådade angående Juda och Jerusalem i Ussias, Jotams, Ahas' och Hiskias, Juda konungars, tid.
Hören, I himlar, och lyssna, du jord; ty HERREN talar.
Barn har jag uppfött och fostrat, men de hava avfallit från mig.
En oxe känner sin ägare och en åsna sin herres krubba, men Israel känner intet, mitt folk förstår intet.
Ve dig, du syndiga släkte, du skuldbelastade folk, du ogärningsmäns avföda, I vanartiga barn, som haven övergivit HERREN, föraktat Israels Helige och vikit bort ifrån honom!
Var skall man mer slå eder, då I så fortgån i avfällighet?
Hela huvudet är ju krankt, och hela hjärtat är sjukt.
Ifrån fotbladet ända upp till huvudet finnes intet helt, blott sårmärken och blånader och friska sår, icke utkramade eller förbundna eller lenade med olja.
Edert land är en ödemark, edra städer äro uppbrända i eld, edra åkrar bliva i eder åsyn förtärda av främlingar; en ödeläggelse är det, såsom där främlingar hava omstörtat allt.
Allenast dottern Sion står kvar där, såsom en hydda i en vingård, såsom ett vaktskjul på ett gurkfält, såsom en inspärrad stad.
Om HERREN Sebaot icke hade lämnat en liten återstod kvar åt oss, då vore vi såsom Sodom, vi vore Gomorra lika.
Hören HERRENS ord, I Sodomsfurstar, lyssna till vår Guds lag, du Gomorra-folk.
Vad skall jag med edra många slaktoffer? säger HERREN.
Jag är mätt på brännoffer av vädurar och på gödkalvars fett, och till blod av tjurar och lamm och bockar har jag intet behag.
När I kommen för att träda fram inför mitt ansikte, vem begär då av eder det, att mina förgårdar trampas ned?
Bären ej vidare fram fåfängliga spisoffer; ångan av dem är en styggelse för mig.
Nymånader och sabbater och utlysta fester, ondska i förening med högtidsförsamlingar, sådant kan jag icke lida.
Edra nymånader och högtider hatar min själ; de hava blivit mig en börda, jag orkar ej bära den.
Ja, huru I än uträcken edra händer, så gömmer jag mina ögon för eder, och om I än mycket bedjen, så hör jag icke därpå.
Edra händer äro fulla av blod;
tvån eder då, och renen eder.
Skaffen edert onda väsende bort ifrån mina ögon.
Hören upp att göra, vad ont är.
Lären att göra vad gott är, faren efter det rätt är, visen förtryckaren på bättre vägar, skaffen den faderlöse rätt, utfören änkans sak.
Kom, låt oss gå till rätta med varandra, säger HERREN.
Om edra synder än äro blodröda, så kunna de bliva snövita, och om de äro röda såsom scharlakan, så kunna de bliva såsom vit ull.
Om I ären villiga att höra, skolen I få äta av landets goda.
Men ären I ovilliga och gensträviga, skolen I förtäras av svärd; ty så har HERRENS mun talat.
Huru har hon icke blivit en sköka, den trogna staden!
Den var full av rätt, rättfärdighet bodde därinne, men nu bo där mördare.
Ditt silver har blivit slagg, ditt ädla vin är utspätt med vatten.
Dina styresmän äro upprorsmän och tjuvars stallbröder.
Alla älskar de mutor och fara efter vinning.
Den faderlöse skaffa de icke rätt, och änkans sak kommer icke inför dem.
Därför säger Herren, HERREN Sebaot, den Starke i Israel: Ve!
Jag vill släcka min harm på mina ovänner och hämnas på mina fiender.
Jag vill vända min hand emot dig och bortrensa ditt slagg såsom med lutsalt och skaffa bort all din oädla malm.
Jag vill åter giva dig sådana domare som tillförne, och sådana rådsherrar som du förut ägde.
Därefter skall du kallas »rättfärdighetens stad», »en trogen stad».
Sion skall genom rätt bliva förlossad och dess omvända genom rättfärdighet.
Men fördärv skall drabba alla överträdare och syndare, och de som övergiva HERREN, de skola förgås.
Ja, de skola komma på skam med de terebinter som voro eder fröjd; och I skolen få blygas över de lustgårdar som I haden så kära.
Ty I skolen bliva såsom en terebint med vissnade löv och varda lika en lustgård utan något vatten.
Och de väldige skola varda såsom blår, och deras verk såsom en gnista, och de skola tillsammans brinna, och ingen skall kunna släcka.
Detta är vad Jesaja, Amos' son, skådade angående Juda och Jerusalem.
Och det skall ske i kommande dagar att det berg där HERRENS hus är skall stå där fast grundat och vara det yppersta ibland bergen och upphöjt över andra höjder; och alla hednafolk skola strömma dit,
ja, många folk skola gå åstad och skola säga: »Upp, låt oss draga åstad till HERRENS berg, upp till Jakobs Guds hus, för att han må undervisa oss om sina vägar, så att vi kunna vandra på hans stigar.»
Ty från Sion skall lag utgå, och HERRENS ord från Jerusalem.
Och han skall döma mellan hednafolken och skipa rätt åt många folk.
Då skola de smida sina svärd till plogbillar och sina spjut till vingårdsknivar.
Folken skola ej mer lyfta svärd mot varandra och icke mer lära sig att strida.
I av Jakobs hus, kommen, låtom oss vandra i HERRENS ljus.
Ty du har förskjutit ditt folk, Jakobs hus, därför att de äro fulla av Österlandets väsende och öva teckentyderi såsom filistéerna; ja, med främlingar förbinda de sig.
Deras land är fullt av silver och guld, och på deras skatter är ingen ände; deras land är fullt av hästar, och på deras vagnar är ingen ände;
deras land är ock fullt av avgudar, och sina egna händers verk tillbedja de, det som deras fingrar hava gjort.
Därför bliva människorna nedböjda och männen ödmjukade; du kan icke förlåta dem.
Fly in i klippan, och göm dig i jorden, för HERRENS fruktansvärda makt och för hans höga majestät.
Ty människornas högmodiga ögon skola bliva ödmjukade, och männens övermod skall bliva nedböjt, och HERREN allena skall vara hög på den dagen.
Ty en dag har HERREN Sebaot bestämt, som skall komma över allt stolt och övermodigt och över allt som är upphöjt, och det skall bliva ödmjukat,
ja, över alla Libanons cedrar, de höga och stolta, och över alla Basans ekar;
över alla höga berg och alla stolta höjder,
över alla höga torn och alla fasta murar,
över alla Tarsis-skepp, ja, över allt som är skönt att skåda.
Och människornas högmod skall bliva nedböjt och männens övermod nedbrutet, och HERREN allena skall vara hög på den dagen.
Men avgudarna skola alldeles förgås.
Och man skall fly in i klippgrottor och in i jordhålor, för HERRENS fruktansvärda makt och för hans höga majestät, när han står upp för att förskräcka jorden.
På den dagen skola människorna kasta bort åt mullvadar och flädermöss de avgudar av silver och de avgudar av guld, som de hava gjort åt sig för att tillbedja.
Ja, de skola fly in i klipprämnor och in i bergsklyftor, för HERRENS fruktansvärda makt och för hans höga majestät, när han står upp för att förskräcka jorden.
Så förliten eder nu ej mer på människor, i vilkas näsa är allenast en fläkt; ty huru ringa äro icke de att akta!
Ty se, Herren, HERREN Sebaot skall taga bort ifrån Jerusalem och Juda allt slags stöd och uppehälle -- all mat till uppehälle och all dryck till uppehälle --
hjältar och krigsmän, domare och profeter, spåmän och äldste,
underhövitsmän och högtuppsatta män, rådsherrar och slöjdkunnigt folk och män som äro förfarna i besvärjelsekonst.
Och jag skall giva dem ynglingar till furstar, och barnsligt självsvåld skall få råda över dem.
Av folket skall den ene förtrycka den andre, var och en sin nästa; den unge skall sätta sig upp mot den gamle, den ringe mot den högt ansedde.
När då så sker, att någon fattar tag i en annan i hans faders hus och säger: »Du äger en mantel, du skall bliva vår styresman; tag du hand om detta vacklande rike» --
då skall denne svara och säga: »Jag kan icke skaffa bot; i mitt hus finnes varken bröd eller mantel.
Mig skolen I icke sätta till styresman över folket.»
Ty Jerusalem vacklar, och Juda faller, då de nu med sitt tal och sina gärningar stå emot HERREN och äro gensträviga mot hans härlighets blickar.
Deras uppsyn vittnar emot dem; och likasom Sodoms folk bedriva de sina synder uppenbart och dölja dem icke.
Ve över deras själar, ty själva hava de berett sig olycka!
Om den rättfärdige mån I tänka att det skall gå honom väl, ty sådana skola äta sina gärningars frukt.
Men ve över den ogudaktige!
Honom skall det gå illa, ty efter hans gärningar skall hans vedergällning bliva.
Mitt folks behärskare är ett barn, och kvinnor råda över det.
Mitt folk, dina ledare föra dig vilse och fördärva den väg, som du skulle gå.
Men HERREN står redo att gå till rätta, han träder fram för att döma folken;
HERREN vill gå till doms med sitt folks äldste och med dess furstar. »I haven skövlat vingården; rov från de fattiga är i edra hus.
Huru kunnen I så krossa mitt folk och söndermala de fattiga?»
Så säger Herren, HERREN Sebaot.
Och HERREN säger: Eftersom Sions döttrar äro så högmodiga, och gå med rak hals och spela med ögonen, och gå där och trippa och pingla med sina fotringar,
därför skall Herren låta Sions döttrars hjässor bliva fulla av skorv, och HERREN skall blotta deras blygd.
På den dagen skall Herren taga bort all deras ståt: fotringar, pannband och halsprydnader,
örhängen, armband och slöjor,
huvudprydnader, fotstegskedjor, gördlar, luktflaskor och amuletter,
fingerringar och näsringar,
högtidsdräkter, kåpor, mantlar och pungar,
speglar, fina linneskjortor, huvudbindlar och flor.
Och där skall vara stank i stället för vällukt, rep i stället för bälte, skalligt huvud i stället för krusat hår, hölje av säcktyg i stället för högtidsmantel, märken av brännjärn i stället för skönhet.
Dina män skola falla för svärd och dina hjältar i krig:
hennes portar skola klaga och sörja, och övergiven skall hon sitta på marken.
Och på den tiden skola sju kvinnor fatta i en och samma man och säga: »Vi vilja själva föda oss och själva kläda oss; låt oss allenast få bära ditt namn, och tag så bort vår smälek.»
På den tiden skall det som HERREN låter växa bliva till prydnad och härlighet, och vad landet alstrar bliva till berömmelse och ära, för den räddade skaran i Israel.
Och det skall ske att den som lämnas övrig i Sion och den som bliver kvar i Jerusalem, han skall då kallas helig, var och en som är upptecknad till liv i Jerusalem --
när en gång Herren har avtvått Sions döttrars orenlighet och bortsköljt ur Jerusalem dess blodskulder genom rättens och reningens ande.
Och HERREN skall över hela Sions bergs område och över dess högtidsskaror skapa en molnsky och en rök om dagen, och skenet av en lågande eld om natten; ty ett beskärmande täckelse skall vila över all dess härlighet.
Och ett skygd skall vara däröver till skugga under dagens hetta, och till en tillflykt och ett värn mot störtskurar och regn.
Jag vill sjunga om min vän, min väns sång om hans vingård.
Min vän hade en vingård på en bördig bergskulle.
Och han hackade upp den och rensade den från stenar och planterade där ädla vinträd; han byggde ett vakttorn därinne, han högg ock ut ett presskar däri.
Så väntade han att den skulle bära äkta druvor, men den bar vilddruvor.
Och nu, I Jerusalems invånare och I Juda män, fällen nu eder dom mellan mig och min vingård.
Vad kunde mer göras för min vingård, än vad jag har gjort för den?
Varför bar den då vilddruvor, när jag väntade att den skulle bära äkta druvor?
Så vill jag nu kungöra för eder vad jag skall göra med min vingård: Jag skall taga bort dess hägnad, och den skall givas till skövling; jag skall bryta ned dess mur, och den skall bliva nedtrampad.
Jag skall i grund fördärva den, ingen skall skära den eller gräva däri.
Den skall fyllas med tistel och törne; och molnen skall jag förbjuda att sända ned regn på den.
Ty HERREN Sebaots vingård, det är Israels hus; och Juda folk är hans älsklingsplantering.
Men när han väntade laglydnad, då fann han lagbrott, och när han väntade rättfärdighet, fann han skriande orättfärdighet. --
Ve eder som läggen hus till hus och fogen åker till åker, intill dess att rum ej mer finnes och I ären de enda som bo i landet!
Från HERREN Sebaot ljuder det så i mina öron: Sannerligen, de många husen skola bliva öde; huru stora och sköna de än äro, skola de bliva tomma på invånare.
Ty en vingård på tio plogland skall giva allenast ett batmått, och en homers utsäde skall giva blott en efa.
Ve dem som stå bittida upp för att hasta till starka drycker, och som sitta intill sena natten för att upphetta sig med vin!
Harpor och psaltare, pukor och flöjter och vin hava de vid sina dryckeslag, men på HERRENS gärningar akta de icke, på hans händers verk se de icke.
Därför skall mitt folk oförtänkt föras bort i fångenskap; dess ädlingar skola lida hunger och dess larmande skaror försmäkta av törst.
Ja, därför spärrar dödsriket upp sitt gap, det öppnar sina käftar utan allt mått, och stadens yperste måste fara ditned, jämte dess larmande och sorlande skaror, envar som fröjdar sig därinne.
Så bliva människorna nedböjda och männen ödmjukade, ja, ödmjukade varda de högmodigas ögon.
Men HERREN Sebaot bliver hög genom sin dom, Gud, den helige, bevisar sig helig genom rättfärdighet.
Och lamm gå där i bet såsom på sin egen mark, och på de rikas ödetomter söka vandrande herdar sin föda.
Ve dem som draga fram missgärningsstraff med lögnens tåg och syndastraff såsom med vagnslinor,
dem som säga: »Må han hasta, må han skynda med sitt verk, så att vi få se det; må det som Israels Helige har beslutit nalkas och komma, så att vi förnimma det!»
Ve dem som kalla det onda gott, och det goda ont, dem som göra mörker till ljus, och ljus till mörker, dem som göra surt till sött, och sött till surt!
Ve dem som äro visa i sina egna ögon och hålla sig själva för kloka!
Ve dem som äro hjältar i att dricka vin och som äro tappra i att blanda starka drycker,
dem som giva den skyldige rätt för mutors skull, men beröva den oskyldige vad som är hans rätt!
Därför, såsom eldsflamman förtär strå, och såsom halm sjunker tillsammans i lågan, så skall deras rot förruttna, och deras löv skola flyga bort såsom stoft, eftersom de förkastade HERREN Sebaots lag och föraktade Israels Heliges ord.
Därför har HERRENS vrede upptänts mot hans folk, och han uträcker sin hand emot det och slår det, så att bergen darra, och så att döda kroppar ligga såsom orenlighet på gatorna.
Vid allt detta vänder hans vrede icke åter, hans hand är ännu uträckt.
Och han reser upp ett baner för hednafolken i fjärran, och lockar på dem att de skola komma från jordens ända; och se, snart och med hast komma de dit.
Ingen finnes bland dem, som är trött, ingen som är stapplande.
Ingen unnar sig slummer och ingen sömn; på ingen lossnar bältet omkring hans länder, och för ingen brister en skorem sönder.
Deras pilar äro skarpa, och deras bågar äro alla spända; deras hästars hovar äro såsom av flinta, och deras vagnshjul likna stormvinden.
Deras skriande är såsom en lejoninnas; de skria såsom unga lejon, rytande gripa de sitt rov och bära bort det, och ingen finnes, som räddar.
Ett rytande över folket höres på den dagen, likt rytandet av ett hav; och skådar man ned på jorden, se, då är där mörker och nöd, och ljuset är förmörkat genom töcken.
I det år då konung Ussia dog såg jag Herren sitta på en hög och upphöjd tron, och släpet på hans mantel uppfyllde templet.
Serafer stodo omkring honom.
Var och en av dem hade sex vingar: med två betäckte de sina ansikten, med två betäckte de sina fötter, och med två flögo de.
Och den ene ropade till den andre och sade: »Helig, helig, helig är HERREN Sebaot; hela jorden är full av hans härlighet.»
Och dörrtrösklarnas fästen darrade, när ropet ljöd; och huset blev uppfyllt av rök.
Då sade jag: »Ve mig, jag förgås!
Ty jag har orena läppar, och jag bor ibland ett folk som har orena läppar, och mina ögon hava sett Konungen, HERREN Sebaot.»
Men en av seraferna flög fram till mig, och han hade i sin hand ett glödande kol, som han med en tång hade tagit på altaret.
Och han rörde därmed vid min mun.
Därefter sade han: »Se, då nu detta har rört vid dina läppar, har din missgärning blivit tagen ifrån dig, och din synd är försonad.»
Och jag hörde Herren tala, och han sade: »Vem skall jag sända, och vem vill vara vår budbärare?»
Och jag sade: »Se, här är jag, sänd mig.»
Då sade han: »Gå åstad och säg till detta folk: 'Hören alltjämt, men förstån intet; sen alltjämt, men förnimmen intet'.
Förstocka detta folks hjärta, och tillslut dess öron, och förblinda dess ögon, så att det icke kan se med sina ögon, eller höra med sina öron, eller förstå med sitt hjärta, och omvända sig och bliva helat.»
Men jag sade: »För huru lång tid, Herre?»
Han svarade: »Till dess att städerna bliva öde och utan någon invånare, och husen utan folk, och till dess att fälten ligga öde och förhärjade.
Och när HERREN har fört folket bort i fjärran och ödsligheten bliver stor i landet,
och allenast en tiondedel ännu är kvar däri, då skall denna ytterligare förödas såsom en terebint eller en ek av vilken en stubbe har lämnats kvar, när den fälldes.
Den stubben skall vara en helig säd.»
Och i Ahas', Jotams sons, Ussias sons, Juda konungs, tid hände sig att Resin, konungen i Aram, och Peka, Remaljas son, Israels konung, drogo upp mot Jerusalem för att erövra det (vilket de likväl icke förmådde göra).
Och när det blev berättat för Davids hus att araméerna hade lägrat sig i Efraim, då skälvde hans och hans folks hjärtan, såsom skogens träd skälva för vinden.
Men HERREN sade till Jesaja: »Gå åstad med din son Sear-Jasub och möt Ahas vid ändan av Övre dammens vattenledning, på vägen till Valkarfältet,
och säg till honom: Tag dig till vara och håll dig stilla; frukta icke och var icke försagd i ditt hjärta för dessa två rykande brandstumpar, för Resin med araméerna och för Remaljas son, i deras förgrymmelse.
Eftersom Aram med Efraim och Remaljas son hava gjort upp onda planer mot dig och sagt:
'Vi vilja draga upp mot Juda och slå det med skräck och erövra det åt oss och göra Tabals son till konung där',
därför säger Herren, HERREN: Det skall icke lyckas, det skall icke ske.
Ty Damaskus är Arams huvud, och Resin är Damaskus' huvud; och om sextiofem år skall Efraim vara krossat, så att det icke mer är ett folk.
Och Samaria är Efraims huvud, och Remaljas son är Samarias huvud.
Om I icke haven tro, skolen I icke hava ro.»
Och HERREN talade ytterligare till Ahas och sade:
»Begär ett tecken från HERREN, din Gud; du må begära det vare sig nedifrån djupet eller uppifrån höjden.»
Men Ahas svarade: »Jag begär intet, jag vill icke fresta HERREN.»
Då sade han: »Så hören då, I av Davids hus: Är det eder icke nog att I sätten människors tålamod på prov?
Viljen I ock pröva min Guds tålamod?
Så skall då Herren själv giva eder ett tecken: Se, den unga kvinnan skall varda havande och föda en son, och hon skall giva honom namnet Immanuel.
Gräddmjölk och honung skall bliva hans mat inemot den tid då han förstår att förkasta vad ont är och utvälja vad gott är.
Ty innan gossen förstår att förkasta vad ont är och utvälja vad gott är, skall det land för vars båda konungar du gruvar dig vara öde.
Och över dig och över ditt folk och över din faders hus skall HERREN låta dagar komma, sådana som icke hava kommit allt ifrån den tid då Efraim skilde sig från Juda: konungen i Assyrien.
Ty på den tiden skall HERREN locka på flugorna längst borta vid Egyptens strömmar och på bisvärmarna i Assyriens land;
och de skola komma och slå ned, alla tillhopa, i bergsdälder och stenklyftor, i alla törnsnår och på alla betesmarker.
På den tiden skall HERREN med en rakkniv som tingas på andra sidan floden -- nämligen med konungen i Assyrien -- raka av allt hår både på huvudet och nedtill; ja, också skägget skall den taga bort.
På den tiden skall en kviga och två tackor vara vad en man föder upp.
Men han skall få mjölk i sådan myckenhet att han kan leva av gräddmjölk; ja, alla som finnas kvar i landet skola leva av gräddmjölk och honung.
Och det skall ske på den tiden, att där nu tusen vinträd stå, värda tusen siklar silver, där skall överallt växa tistel och törne.
Med pilar och båge skall man gå dit, ty hela landet skall vara tistel och törne.
Och alla de berg där man nu arbetar med hackan, dem skall man ej mer beträda, av fruktan för tistel och törne; de skola bliva platser dit oxar drivas, och marker som trampas ned av får.»
Och HERREN sade till mig: »Tag dig en stor tavla och skriv på den med tydlig stil Maher-salal Has-bas.
Och jag vill taga mig pålitliga vittnen: prästen Uria och Sakarja, Jeberekjas son.»
Och jag gick in till profetissan, och hon blev havande och födde en son.
Och HERREN sade till mig: »Giv honom namnet Maher-salal Has-bas.
Ty förrän gossen kan säga 'fader' och 'moder' skall man bära Damaskus' skatter och byte från Samaria fram för konungen i Assyrien.»
Och HERREN talade vidare till mig och sade:
»Eftersom detta folk föraktar Siloas vatten, som flyter så stilla, och har sin fröjd med Resin och Remaljas son,
se, därför skall HERREN låta komma över dem flodens vatten, de väldiga och stora, nämligen konungen i Assyrien med all hans härlighet.
Och den skall stiga över alla sina bräddar och gå över alla sina stränder.
Den skall tränga fram i Juda, svämma över och utbreda sig och räcka ända upp till halsen; och med sina utbredda vingar, skall den uppfylla ditt land, Immanuel, så vitt det är.»
Rasen, I folk; I skolen dock krossas.
Lyssnen, alla I fjärran länder.
Rusten eder; I skolen dock krossas.
Ja, rusten eder; I skolen dock krossas.
Gören upp planer; de varda dock om intet.
Avtalen, vad I viljen; det skall dock ej lyckas.
Ty Gud är med oss.
Ty så sade HERREN till mig, när hans hand kom över mig med makt och han varnade mig för att vandra på detta folks väg:
I skolen icke kalla för sammansvärjning allt vad detta folk kallar sammansvärjning, ej heller skolen I frukta vad det fruktar, I skolen icke förskräckas därför.
Nej, HERREN Sebaot skolen I hålla helig; honom skolen I frukta, och för honom skolen I förskräckas.
Så skall han varda för eder något heligt; men för de två Israels hus skall han bliva en stötesten och en klippa till fall och för Jerusalems invånare en snara och ett giller.
Många av dem skola stupa därpå, de skola falla och krossas, de skola snärjas och varda fångade.
Lägg vittnesbördet ombundet och lagen förseglad i mina lärjungars hjärtan.
Så vill jag förbida HERREN, då han nu döljer sitt ansikte för Jakobs hus; jag vill vänta efter honom.
Se, jag och barnen som HERREN har givit mig, vi äro tecken och förebilder i Israel, från HERREN Sebaot, som bor på Sions berg.
Och när man säger till eder: »Frågen andebesvärjare och spåmän, dem som viska och mumla», så svaren: »Skall icke ett folk fråga sin Gud?
Skall man fråga de döda för de levande?»
»Nej, hållen eder till lagen, till vittnesbördet!»
Så skola förvisso en gång de nödgas mana, för vilka nu ingen morgonrodnad finnes.
De skola draga omkring i landet, nedtryckta och hungrande, och i sin hunger skola de förbittras och skola förbanna sin konung och sin Gud.
Och de skola vända blicken uppåt, de skola ock skåda ned på jorden;
men se, där är nöd och mörker och natt av ångest.
Ja, tjockt mörker är de fördrivnas liv.
Dock, natt skall icke förbliva där nu ångest råder.
I den förgångna tiden har har han låtit Sebulons och Naftalis land vara ringa aktat, men i framtiden skall han låta det komma till ära, trakten utmed Havsvägen, landet på andra sidan Jordan, hedningarnas område.
Det folk som vandrar i mörkret skall se ett stort ljus; ja, över dem som bo i dödsskuggans land skall ett ljus skina klart.
Du skall göra folket talrikt, du skall göra dess glädje stor; inför dig skola de glädja sig, såsom man glädes under skördetiden, såsom man fröjdar sig, när man utskiftar byte.
Ty du skall bryta sönder deras bördors ok och deras skuldrors gissel och deras plågares stav, likasom i Midjans tid.
Och skon som krigaren bar i stridslarmet, och manteln som sölades i blod, allt sådant skall brännas upp och förtäras av eld.
Ty ett barn varder oss fött, en son bliver oss given, och på hans skuldror skall herradömet vila; och hans namn skall vara: Underbar i råd, Väldig Gud, Evig fader, Fridsfurste.
Så skall herradömet varda stort och friden utan ände över Davids tron och över hans rike; så skall det befästas och stödjas med rätt och rättfärdighet, från nu och till evig tid.
HERREN Sebaots nitälskan skall göra detta.
Ett ord sänder Herren mot Jakob, och det slår ned i Israel,
och allt folket får förnimma det, Efraim och Samarias invånare, de som säga i sitt övermod och i sitt hjärtas stolthet:
»Tegelmurar hava fallit, men med huggen sten bygga vi upp nya; mullbärsfikonträd har man huggit ned, men cederträd sätta vi i deras ställe.»
Och HERREN uppreser mot dem Resins ovänner och uppeggar deras fiender,
araméerna från den ena sidan och filistéerna från den andra, och de äta upp Israel med glupska gap.
Vid allt detta vänder hans vrede icke åter, hans hand är ännu uträckt.
Men folket vänder ej åter till honom som slår dem; Herren Sebaot söka de icke.
Därför avhugger HERREN på Israel både huvud och svans, han hugger av både palmtopp och sävstrå, allt på en dag --
de äldste och högst uppsatte de äro huvudet, och profeterna, de falska vägvisarna, de äro svansen.
Ty detta folks ledare föra det vilse, och de som låta leda sig gå i fördärvet.
Därför kan Herren icke glädja sig över dess unga män, ej heller hava förbarmande med dess faderlösa och änkor; ty de äro allasammans gudlösa ogärningsmän, och var mun talar dårskap.
Vid allt detta vänder hans vrede icke åter, hans hand är ännu uträckt.
Ty ogudaktigheten förbränner såsom en eld, den förtär tistel och törne; den tänder på den tjocka skogen, så att den går upp i höga virvlar av rök.
Genom HERREN Sebaots förgrymmelse har landet råkat i brand, och folket är likasom eldsmat; den ene skonar icke den andre.
Man river åt sig till höger och förbliver dock hungrig, man tager för sig till vänster och bliver dock ej mätt; envar äter köttet på sin egen arm:
Manasse äter Efraim, och Efraim Manasse, och båda tillhopa vända sig mot Juda.
Vid allt detta vänder hans vrede icke åter, hans hand är ännu uträckt.
Ve eder som stadgen orättfärdiga stadgar!
I skriven, men våldslagar skriven I
för att vränga de ringas sak och beröva de fattiga i mitt folk deras rätt, för att göra änkor till edert byte och plundra de faderlösa.
Vad viljen I göra på hemsökelsens dag, när ovädret kommer fjärran ifrån?
Till vem viljen I fly för att få hjälp, och var viljen I lämna edra skatter i förvar?
Om man ej böjer knä såsom fånge, så måste man falla bland de dräpta.
Vid allt detta vänder hans vrede icke åter, hans hand är ännu uträckt.
Ve över Assur, min vredes ris, som bär min ogunst såsom en stav i sin hand!
Mot ett gudlöst folk sänder jag honom, och mot min förgrymmelses folk bjuder jag honom gå, för att taga rov och göra byte, och för att nedtrampa det såsom orenlighet på gatorna.
Men så menar icke han, och i sitt hjärta tänker han ej så, utan hans hjärta står efter att förgöra och efter att utrota folk i mängd.
Han säger: »Äro mina hövdingar ej allasammans konungar?
Har det icke gått Kalno såsom Karkemis, och Hamat såsom Arpad, och Samaria såsom Damaskus?
Då min hand har träffat de andra gudarnas riken, vilkas beläten voro förmer än Jerusalems och Samarias,
skulle jag då ej kunna göra med Jerusalem och dess gudabilder vad jag har gjort med Samaria och dess gudar?»
Men när Herren har fullbordat allt sitt verk på Sions berg och i Jerusalem, då skall jag hemsöka den assyriske konungens hjärtas högmodsfrukt och hans stolta ögons förhävelse.
Ty han säger: »Med min hands kraft har jag utfört detta och genom min vishet, ty jag har förstånd.
Jag flyttade folkens gränser, deras förråd utplundrade jag, och i min väldighet stötte jag härskarna från tronen.
Och min hand grep efter folkens skatter såsom efter fågelnästen, och såsom man samlar övergivna ägg, så samlade jag jordens alla länder; ingen fanns, som rörde vingen eller öppnade näbben till något ljud.»
Skall då yxan berömma sig mot honom som hugger med den, eller sågen förhäva sig mot honom som sätter den i rörelse?
Som om käppen satte i rörelse honom som lyfter den, eller staven lyfte en som dock är förmer än ett stycke trä!
Så skall då Herren, HERREN Sebaot sända tärande sjukdom i hans feta kropp, och under hans härlighet skall brinna en brand likasom en brinnande eld.
Och Israels ljus skall bliva en eld och hans Helige en låga, och den skall bränna upp och förtära dess törnen och dess tistlar, allt på en dag.
Och på hans skogars och parkers härlighet skall han alldeles göra en ände; det skall vara, såsom när en sjuk täres bort.
De träd som bliva kvar i hans skog skola vara lätt räknade; ett barn skall kunna teckna upp dem.
På den tiden skall kvarlevan av Israel och den räddade skaran av Jakobs hus ej vidare stödja sig vid honom som slog dem; i trohet skola de stödja sig vid HERREN, Israels Helige.
En kvarleva skall omvända sig, en kvarleva av Jakob, till Gud, den väldige.
Ty om än ditt folk, Israel, vore såsom sanden i havet, så skall dock allenast en kvarleva där omvända sig.
Förödelsen är oryggligt besluten, den kommer med rättfärdighet såsom en flod.
Ty förstöring och oryggligt besluten straffdom skall Herren, HERREN Sebaot låta komma över hela jorden.
Därför säger Herren, HERREN Sebaot så: Frukta icke, mitt folk, du som bor i Sion, för Assur, när han slår dig med riset och upplyfter sin stav mot dig, såsom man gjorde i Egypten.
Ty ännu allenast en liten tid, och ogunsten skall hava en ände, och min vrede skall vända sig till deras fördärv.
Och HERREN Sebaot skall svänga sitt gissel över dem, såsom när han slog Midjan vid Orebsklippan; och sin stav, som han räckte ut över havet, skall han åter upplyfta, såsom han gjorde i Egypten.
På den tiden skall hans börda tagas bort ifrån din skuldra och hans ok ifrån din hals, ty oket skall brista sönder för fetmas skull.
Han kommer över Ajat, han drager fram genom Migron; i Mikmas lämnar han sin tross.
De draga fram över passet; i Geba taga de nattkvarter.
Rama bävar; Sauls Gibea flyr.
Ropa högt, du dotter Gallim.
Giv akt, du Laisa.
Arma Anatot!
Madmena flyktar; Gebims invånare bärga sitt gods.
Ännu samma dag står han i Nob; han lyfter sin hand mot dottern Sions berg, mot Jerusalems höjd.
Men se, då avhugger Herren, HERREN Sebaot den lummiga kronan, med förskräckande makt; de resliga stammarna ligga fällda, de höga träden störta ned.
Den tjocka skogen nedhugges med järnet; Libanons skogar falla för den väldige.
Men ett skott skall skjuta upp ur Isais avhuggna stam, och en telning från dess rötter skall bära frukt.
Och på honom skall HERRENS Ande vila, vishets och förstånds Ande, råds och starkhets Ande, HERRENS kunskaps och fruktans Ande.
Han skall hava sitt välbehag i HERRENS fruktan; och han skall icke döma efter som ögonen se eller skipa lag efter som öronen höra.
Utan med rättfärdighet skall han döma de arma och med rättvisa skipa lag åt de ödmjuka på jorden.
Och han skall slå jorden med sin muns stav, och med sina läppars anda döda de ogudaktiga.
Rättfärdighet skall vara bältet omkring hans länder och trofasthet bältet omkring hans höfter.
Då skola vargar bo tillsammans med lamm och pantrar ligga tillsammans med killingar; och kalvar och unga lejon och gödboskap skola sämjas tillhopa, och en liten gosse skall valla dem.
Kor och björnar skola gå och beta, deras ungar skola ligga tillhopa, och lejon skola äta halm likasom oxar.
Ett spenabarn skall leka invid en huggorms hål och ett avvant barn sträcka ut sin hand efter basiliskens öga.
Ingenstädes på mitt heliga berg skall man då göra vad ont och fördärvligt är, ty landet skall vara fullt av HERRENS kunskap, likasom havsdjupet är fyllt av vattnet.
Och det skall ske på den tiden att hednafolken skola söka telningen från Isais rot, där han står såsom ett baner för folken; och hans boning skall vara idel härlighet.
Och HERREN skall på den tiden ännu en gång räcka ut sin hand, för att förvärva åt sig kvarlevan av sitt folk, vad som har blivit räddat från Assyrien, Egypten, Patros, Etiopien, Elam, Sinear, Hamat och havsländerna.
Och han skall resa upp ett baner för hednafolken och samla Israels fördrivna män; och Juda förskingrade kvinnor skall han hämta tillhopa från jordens fyra hörn.
Då skall Efraims avund upphöra och Juda ovänskap bliva utrotad; Efraim skall ej hysa avund mot Juda, och Juda icke ovänskap mot Efraim.
Men såsom rovfåglar skola de slå ned på filistéernas skuldra västerut, tillsammans skola de taga byte av österlänningarna; Edom och Moab skola gripas av deras hand, och Ammons barn skola bliva dem hörsamma.
Och HERREN skall giva till spillo Egyptens havsvik och lyfta sin hand mot floden i förgrymmelse; och han skall klyva den i sju bäckar och göra så, att man torrskodd kan gå däröver.
Så skall där bliva en banad väg för den kvarleva av hans folk, som har blivit räddad från Assur, likasom det var för Israel på den dag då de drogo upp ur Egyptens land.
På den tiden skall du säga: »Jag tackar dig, HERRE, ty väl var du vred på mig, men din vrede har upphört, och du tröstar mig.
Se, Gud är min frälsning, jag är trygg och fruktar icke; ty HERREN, HERREN är min starkhet och min lovsång, och han blev mig till frälsning.»
Och I skolen ösa vatten med fröjd ur frälsningens källor
och skolen säga på den tiden: »Tacken HERREN, åkallen hans namn, gören hans gärningar kunniga bland folken; förtäljen att hans namn är högt.
Lovsjungen HERREN, ty han har gjort härliga ting; detta vare kunnigt över hela jorden.
Ropen av fröjd och jublen, I Sions invånare, ty Israels Helige är stor bland eder.
Detta är en utsaga om Babel, vad som uppenbarades för Jesaja, Amos' son.
Resen upp ett baner på ett kalt berg, ropen högt till dem; viften med handen att de må draga in genom de mäktiges portar.
Jag själv har bådat upp mina invigda, ja, kallat mina hjältar till mitt vredesverk, min stolta skara, som jublar.
Hör, det larmar på bergen såsom av ett stort folk.
Hör, det sorlar av riken med hopade hednafolk.
HERREN Sebaot mönstrar sin krigarskara.
Ifrån fjärran land komma de, ifrån himmelens ända, HERREN och hans vredes redskap, för att fördärva hela jorden.
Jämren eder, ty nära är HERRENS dag; såsom våld från den Allsvåldige kommer den.
Därför sjunka alla händer ned, och alla människohjärtan förfäras.
Man förskräckes, man gripes av ångest och kval, ja, våndas såsom en barnaföderska.
Häpen stirrar den ene på den andre; röda såsom eldslågor äro deras ansikten.
Se, HERRENS dag kommer, gruvlig och med förgrymmelse och med vredesglöd, för att göra jorden till en ödemark och utrota syndarna som där bo.
Ty himmelens stjärnor och stjärnbilder sända ej mer ut sitt ljus, solen går mörk upp, och månens ljus skiner icke.
Jag skall hemsöka jordens krets för dess ondska och de ogudaktiga för deras missgärning; jag skall göra slut på de fräckas övermod och slå ned våldsverkarnas högmod.
Jag skall göra en man mer sällsynt än fint guld, en människa mer sällsynt än guld från Ofir.
Därför skall jag komma himmelen att darra, och jorden skall bäva och vika från sin plats -- genom HERREN Sebaots förgrymmelse, på hans glödande vredes dag.
Och likasom jagade gaseller och en hjord som ingen samlar vända de då hem, var och en till sitt folk, och fly, var och en till sitt land.
Men envar som upphinnes bliver genomborrad, och envar som gripes faller för svärd.
Deras späda barn krossas inför deras ögon, deras hus plundras, och deras kvinnor skändas.
Ty se, jag vill uppväcka mot dem mederna, som akta silver för intet och icke fråga efter guld.
Deras bågar skola fälla de unga männen, med frukten i moderlivet hava de intet förbarmande, och barnen skona de icke.
Och det skall gå med Babel, rikenas krona, kaldéernas ära och stolthet, likasom när Gud omstörtade Sodom och Gomorra.
Aldrig mer skall det bliva bebyggt, från släkte till släkte skall det ligga obebott; ingen arab skall där slå upp sitt tält, ingen herde lägra sig där med sin hjord.
Nej, öknens djur skola lägra sig där, och dess hus skola fyllas av uvar; strutsar skola bo där, och gastar skola hoppa där.
Schakaler skola tjuta i dess palatser och ökenhundar i praktbyggnaderna.
Snart kommer dess tid; dess dagar skola ej fördröjas.
Ty HERREN skall förbarma sig över Jakob och ännu en gång utvälja Israel och låta dem komma till ro i deras land; och främlingar skola sluta sig till dem och hålla sig till Jakobs hus.
Och folk skola taga dem och föra dem hem igen; men Israels hus skall lägga dem under sig såsom sin arvedel i HERRENS land, och skall göra dem till trälar och trälinnor.
Så skola de få sina fångvaktare till fångar och råda över sina plågare.
Och på den dag då HERREN låter dig få ro från din vedermöda och ångest, och från den hårda träldom som har varit dig pålagd,
då skall du stämma upp denna visa över konungen i Babel, du skall säga: »Vilken ände har icke plågaren fått, vilken ände pinoorten!
HERREN har brutit sönder de ogudaktigas stav, tyrannernas ris,
det ris som i grymhet slog folken med slag på slag, och i vrede härskade över folkslagen med skoningslös förföljelse.
Hela jorden har nu fått vila och ro; man brister ut i jubel.
Själva cypresserna glädja sig över ditt fall, så ock Libanons cedrar: 'Sedan du nu ligger där, drager ingen hitupp för att hugga ned oss.'
Dödsriket därnere störes i sin ro för din skull, när det måste taga emot dig.
Skuggorna där väckas upp för din skull, jordens alla väldige; folkens alla konungar måste stå upp från sina troner.
De upphäva alla sin röst och säga till dig: 'Så har då också du blivit maktlös såsom vi, ja, blivit vår like.'
Ned till dödsriket har din härlighet måst fara, och dina harpors buller; förruttnelse är bädden under dig, och maskar äro ditt täcke.
Huru har du icke fallit ifrån himmelen, du strålande morgonstjärna!
Huru har du icke blivit fälld till jorden, du folkens förgörare!
Det var du som sade i ditt hjärta: 'Jag vill stiga upp till himmelen; högt ovanför Guds stjärnor vill jag ställa min tron; jag vill sätta mig på gudaförsamlingens berg längst uppe i norr.
Jag vill stiga upp över molnens höjder, göra mig lik den Högste.'
Nej, ned till dödsriket måste du fara, längst ned i graven.
De som se dig stirra på dig, de betrakta dig och säga: 'Är detta den man som kom jorden att darra och riken att bäva,
den som förvandlade jordkretsen till en öken och förstörde dess städer, den som aldrig frigav sina fångar, så att de fingo återvända hem?'
Folkens alla konungar ligga allasammans med ära var och en i sitt vilorum;
men du ligger obegraven och bortkastad, lik en föraktad gren; du ligger där överhöljd av dräpta, av svärdsslagna män, av döda som hava farit ned i gravkammaren, lik ett förtrampat as.
Du skulle icke såsom de få vila i en grav, ty du fördärvade ditt land och dräpte ditt folk.
Om ogärningsmännens avföda skall man aldrig mer tala.
Anställen ett blodbad på hans söner för deras fäders missgärning.
De få ej stå upp och besitta jorden och fylla jordkretsens yta med städer.»
Nej, jag skall stå upp emot dem, säger HERREN Sebaot; och jag skall utrota ur Babel både namn och kvarleva, både barn och efterkommande, säger HERREN.
Och jag skall göra det till ett tillhåll för rördrommar och fylla det med sumpsjöar; ja, jag skall bortsopa det med ödeläggelsens kvast, säger HERREN Sebaot.
HERREN Sebaot har svurit och sagt: Sannerligen, såsom jag har tänkt, så skall det ske, och vad jag har beslutit, det skall fullbordas.
Jag skall krossa Assur i mitt land, och på mina berg skall jag förtrampa honom.
Så skall hans ok bliva borttaget ifrån dem och hans börda tagas av deras skuldra.
Detta är det beslut som är fattat mot hela jorden; detta är den hand som är uträckt mot alla folk.
Ty HERREN Sebaot har beslutit det; vem kan då göra det om intet?
Hans hand är det som är uträckt; vem kan avvända den?
I det år då konung Ahas dog förkunnades följande utsaga:
Gläd dig icke, du filistéernas hela land, över att det ris som slog dig är sönderbrutet; ty från ormens rot skall en basilisk komma fram, och dennes avkomma bliver en flygande drake.
De utarmade skola sedan få bete och de fattiga få lägra sig i trygghet; men telningarna från din rot skall jag döda genom hunger, och vad som bliver kvar av dig skall dräpas.
Jämra dig, du port; ropa, du stad; försmält av ångest, du filistéernas hela land.
Ty norrifrån kommer en rök; i fiendeskarornas tåg bliver ingen efter.
Vad skall man då svara det främmande folkets sändebud?
Jo, att det är HERREN som har grundat Sion, och att de betryckta bland hans folk där hava sin tillflykt.
Utsaga om Moab.
Ja, med Ar-Moab är det ute den natt då det förstöres.
Ja, med Kir-Moab är det ute den natt då det förstöres.
Habbait och Dibon stiga upp på offerhöjderna för att gråta; uppe i Nebo och Medeba jämrar sig Moab; alla huvuden där äro skalliga, alla skägg avskurna.
På dess gator bär man sorgdräkt, så ock på dess tak; på dess torg jämra sig alla och flyta i tårar.
Hesbon och Eleale höja klagorop, så att det höres ända till Jahas.
Därför skria ock Moabs krigare; hans själ våndas i honom.
Mitt hjärta klagar över Moab, ty hans flyktingar fly ända till Soar, till Eglat-Selisia; uppför Halluhits höjd stiger man under gråt, och på vägen till Horonaim höjas klagorop över förstörelsen.
Nimrims vatten bliva torr ökenmark, gräset förtorkas, brodden vissnar, intet grönt lämnas kvar.
Återstoden av sitt förvärv, sitt sparda gods, bär man därför nu bort över Pilträdsbäcken.
Ja, klagoropen ljuda runtom i Moabs land; till Eglaim når dess jämmer och till Beer-Elim dess jämmer.
Dimons vatten äro fulla av blod.
Ja, ännu något mer skall jag låta komma över Dimon; ett lejon över Moabs räddade, över det som bliver kvar av landet.
»Sänden åstad de lamm som landets herre bör hava från Sela genom öknen till dottern Sions berg.»
Och såsom flyktande fåglar, lika skrämda fågelungar komma Moabs döttrar till Arnons vadställen.
De säga: »Giv oss råd, bliv medlare för oss.
Låt din skugga vara såsom natten, nu mitt i middagshettan.
Skydda de fördrivna; röj icke de flyktande.
Låt mina fördrivna finna härbärge hos dig, var för Moab ett beskärm mot fördärvaren, till dess att utpressaren ej mer är till och fördärvet får en ände och förtryckarna försvinna bort ur landet.
Så skall genom eder mildhet eder tron bliva befäst, och på den skall sitta trygg i Davids hydda en furste som far efter vad rätt är och främjar rättfärdighet.»
Vi hava hört om Moabs högmod, det övermåttan höga, om hans högfärd, högmod och övermod och opålitligheten i hans lösa tal.
Därför måste nu Moab jämra sig över Moab, hela landet måste jämra sig.
Över Kir-Haresets druvkakor måsten I sucka i djup bedrövelse.
Ty Hesbons fält äro förvissnade, så ock Sibmas vinträd, vilkas ädla druvor slogo folkens herrar till marken, vilkas rankor nådde till Jaeser och förirrade sig i öknen, vilkas skott bredde ut sig och gingo över havet.
Därför gråter jag över Sibmas vinträd, såsom Jaeser gråter; med mina tårar vattnar jag dig, Hesbon, och dig, Eleale.
Ty mitt i din sommar och din bärgningstid har ett skördeskri slagit ned.
Glädje och fröjd är nu avbärgad från de bördiga fälten, och i vingårdarna höjes intet glädjerop, höres intet jubel; ingen trampar vin i pressarna, på skördeskriet har jag gjort slut.
Därför klagar mitt hjärta såsom en harpa över Moab, ja, mitt innersta över Kir-Heres.
Ty huru än Moab ävlas att träda upp på offerhöjden och huru han än går in i sin helgedom och beder, så uträttar han intet därmed.
Detta är det ord, som HERREN tillförne talade till Moab.
Men nu har HERREN åter talat och sagt: Inom tre år, såsom dagakarlen räknar åren, skall Moab i sin härlighet, med alla sina stora skaror, varda aktad för intet; och vad som bliver kvar skall vara litet och ringa, icke mycket värt.
Utsaga om Damaskus.
Se, Damaskus skall upphöra att vara en stad; det skall falla och bliva en stenhop.
Aroers städer varda övergivna; de bliva tillhåll för hjordar, som lägra sig där ostörda.
Det är förbi med Efraims värn, med Damaskus' konungadöme och med kvarlevan av Aram.
Det skall gå med dem såsom med Israels barns härlighet, säger HERREN Sebaot.
Och det skall ske på den tiden att Jakobs härlighet vändes i armod, och att hans feta kropp bliver mager.
Det går, såsom när skördemannen samlar ihop säden och med sin arm skördar axen; det går, såsom när man plockar ax i Refaims-dalen:
en ringa efterskörd lämnas kvar där, såsom när man slår ned oliver, två eller tre bär lämnas kvar högst uppe i toppen, fyra eller fem på trädets kvistar, säger HERREN, Israels Gud.
På den tiden skola människorna blicka upp till sin Skapare och deras ögon se upp till Israels Helige.
Människorna skola ej vända sin blick till de altaren som deras händer hava gjort; på sina fingrars verk skola de icke se, icke på Aserorna eller på solstoderna.
På den tiden skola deras fasta städer bliva lika de övergivna fästen i skogarna och på bergstopparna, som övergåvos, när Israels barn drogo in; allt skall bliva ödelagt.
Ty du har förgätit din frälsnings Gud, och du tänker icke på din fasta klippa.
Därför planterar du ljuvliga planteringar och sätter i dem främmande vinträd.
Och väl får du dem att växa högt samma dag du planterar dem, och morgonen därefter får du dina plantor att blomma, men skörden försvinner på hemsökelsens dag, då plågan bliver olidlig.
Hör, det brusar av många folk, det brusar, såsom havet brusar.
Det dånar av folkslag, det dånar, såsom väldiga vatten dåna.
Ja, det dånar av folkslag, såsom stora vatten dåna.
Men han näpser dem, och de fly bort i fjärran; de jagas bort såsom agnar för vinden, uppe på bergen, och såsom virvlande löv för stormen.
När aftonen är inne, se, då kommer förskräckelsen, och förrän morgonen gryr, äro de sin kos.
Detta bliver våra skövlares del, våra plundrares lott.
Hör, du land där flygfän surra, du land bortom Etiopiens strömmar,
du som har sänt budbärare över havet, i rörskepp hän över vattnet!
Gån åstad, I snabba sändebud, till det resliga folket med glänsande hy, till folket som är så fruktat vida omkring, det starka och segerrika folket, vars land genomskäres av strömmar.
I jordkretsens alla inbyggare, I som bon på jorden: sen till, när man reser upp baner på bergen, och när man stöter i basun, så lyssnen därtill.
Ty så har HERREN sagt till mig: »I stillhet vill jag skåda ned från min boning, såsom solglans glöder från en klar himmel, såsom molnet utgjuter dagg under skördetidens hetta.»
Ty förrän skördetiden är inne, just när blomningen är slut och blomman förbytes i mognad druva, skall han avskära rankorna med vingårdskniv och hugga av rotskotten och skaffa dem bort.
Alltsammans skall lämnas till pris åt rovfåglarna på bergen och åt djuren på marken; rovfåglarna skola där hava sina nästen över sommaren och markens alla djur ligga där om vintern.
På den tiden skola skänker bäras fram till HERREN Sebaot från det resliga folket med glänsande hy, från folket som är så fruktat vida omkring, det starka och segerrika folket, vars land genomskäres av strömmar -- till den plats där HERREN Sebaots namn bor, till Sions berg.
Utsaga om Egypten.
Se, HERREN far fram på ett ilande moln och kommer till Egypten.
Egyptens avgudar bäva då för honom, och egyptiernas hjärtan förfäras i deras bröst.
Och jag skall uppegga egyptier mot egyptier, så att broder skall strida mot broder och vän mot vän, stad mot stad och rike mot rike.
Och egyptiernas förstånd skall försvinna ur deras hjärtan, och deras råd skall jag göra om intet; de skola då fråga sina avgudar och signare, sina andebesvärjare och spåmän.
Men jag skall giva egyptierna i en hård herres hand, och en grym konung skall få råda över dem, säger Herren, HERREN Sebaot.
Och vattnet skall försvinna ur havet, och floden skall sina bort och uttorka.
Strömmarna skola utbreda stank, Egyptens kanaler skola förminskas och sina bort; rör och vass skall förvissna.
Ängarna vid Nilfloden, längs flodens strand, och alla sädesfält vid floden, de skola förtorka, fördärvas och varda till intet.
Dess fiskare skola klaga, alla som kasta ut krok i floden skola sörja; och de som lägga ut nät i vattnet skola stå där modlösa.
De som arbeta i häcklat lin skola komma på skam, så ock de som väva fina tyger.
Landets stödjepelare skola bliva krossade och alla de som arbeta för lön gripas av ångest.
Såsom idel dårar stå då Soans furstar; Faraos visaste rådgivare giva blott oförnuftiga råd.
Huru kunnen I då säga till Farao: »Jag är en son av visa män, en son av forntidens konungar»?
Ja, var är dina vise?
Må de förkunna för dig -- ty de veta det ju -- vad HERREN Sebaot har beslutit över Egypten.
Nej, Soans furstar hava blivit dårar, Nofs furstar äro bedragna, Egypten föres vilse av dem som voro hörnstenar i dess stammar.
HERREN har där utgjutit en förvirringens ande, så att de komma Egypten att ragla, vadhelst det företager sig, såsom en drucken raglar i sina spyor.
Och Egypten skall icke hava framgång i vad någon där gör, evad han är huvud eller svans, evad han är palmtopp eller sävstrå.
På den tiden skola egyptierna vara såsom kvinnor: de skola bäva och förskräckas för HERREN Sebaots upplyfta hand, när han lyfter den mot dem.
Och Juda land skall bliva en skräck för egyptierna; så ofta man nämner det för dem, skola de förskräckas, för det besluts skull som HERREN Sebaot har fattat över dem.
På den tiden skola i Egyptens land finnas fem städer som tala Kanaans tungomål, och som svärja vid HERREN Sebaot; en av dem skall heta Ir-Haheres.
På den tiden skall ett altare vara rest åt HERREN mitt i Egyptens land, så ock en stod åt HERREN vid landets gräns.
Och de skola vara till tecken och vittnesbörd för HERREN Sebaot i egyptiernas land: när de ropa till HERREN om hjälp mot förtryckare, då skall han sända dem en frälsare och försvarare, och han skall rädda dem.
Och HERREN skall göra sig känd för egyptierna, ja, egyptierna skola lära känna HERREN på den tiden; och de skola tjäna honom med slaktoffer och spisoffer, de skola göra löften åt HERREN och få infria dem.
Så skall då HERREN slå Egypten -- slå, men ock hela; när de omvända sig till HERREN, skall han bönhöra dem och hela dem.
På den tiden skall en banad väg leda från Egypten till Assyrien, och assyrierna skola komma in i Egypten, och egyptierna in i Assyrien; och egyptierna skola hålla gudstjänst tillsammans med assyrierna.
På den tiden skall Israel, såsom den tredje i förbundet, stå vid sidan av Egypten och Assyrien, till en välsignelse på jorden.
Och HERREN Sebaot skall välsigna dem och säga: Välsignad vare du Egypten, mitt folk, och du Assyrien, mina händer verk, och du Israel, min arvedel!
I det år då Tartan kom till Asdod, utsänd av Sargon, konungen i Assyrien -- varefter han ock belägrade Asdod och intog det --
på den tiden talade HERREN genom Jesaja, Amos' son, och sade: »Upp, lös säcktygsklädnaden från dina länder, och drag dina skor av dina fötter.»
Och denne gjorde så och gick naken och barfota.
Sedan sade HERREN: »Likasom min tjänare Jesaja har gått naken och barfota och nu i tre år varit till tecken och förebild angående Egypten och Etiopien,
så skall konungen i Assyrien låta fångarna ifrån Egypten och de bortförda från Etiopien, både unga och gamla, vandra åstad nakna och barfota, med blottad bak, Egypten till blygd.
Då skola de häpna och blygas över Etiopien, som var deras hopp, och över Egypten, som var deras stolthet.
På den dagen skola inbyggarna här i kustlandet säga: 'Se, så gick det med dem som voro vårt hopp, med dem till vilka vi flydde, för att få hjälp och bliva räddade undan konungen i Assyrien; huru skola vi då själva kunna undkomma?'»
Utsaga om Öknen vid havet.
Likasom en storm som far fram i Sydlandet kommer det från öknen, från det fruktansvärda landet.
En gruvlig syn har blivit mig kungjord: »Härjare härja, rövare röva.
Drag upp, du Elam!
Träng på, du Mediens folk!
På all suckan vill jag göra slut.»
Fördenskull darra nu mina länder, ångest griper mig, lik en barnaföderskas ångest; förvirring kommer över mig, så att jag icke kan höra, förskräckelse fattar mig, så att jag icke kan se.
Mitt hjärta är utom sig, jag kväljes av förfäran; skymningen, som jag längtade efter, vållar mig nu skräck.
Man dukar bord, man breder ut täcken, man äter och dricker.
Nej, stån upp, I furstar; smörjen edra sköldar!
Ty så har Herren sagt till mig: »Gå och ställ ut en väktare; vad han får se, det må han förkunna.
Och om han ser ett tåg, ryttare par efter par, ett tåg av åsnor, ett tåg av kameler, då må han giva akt, noga giva akt.»
Och denne ropade, såsom ett lejon ryter: »Herre, här står jag på vakt beständigt, dagen igenom, och jag förbliver här på min post natt efter natt.
Och se, nu kommer här ett tåg av män, ryttare par efter par!»
Och åter talade han och sade: »Fallet, fallet är Babel!
Alla dess gudabeläten äro nedbrutna till jorden.»
O du mitt krossade, mitt söndertröskade folk, vad jag har hört av HERREN Sebaot, Israels Gud, det har jag förkunnat för eder.
Utsaga om Duma.
Man ropar till mig från Seir: »Väktare, vad lider natten?
Väktare, vad lider natten?»
Väktaren svarar: »Morgon har kommit, och likväl är det natt.
Viljen I fråga mer, så frågen; kommen tillbaka igen.»
Utsaga över Arabien.
Tagen natthärbärge i Arabiens vildmark, I karavaner från Dedan.
Må man komma emot de törstande och giva dem vatten.
Ja, inbyggarna i Temas land gå de flyktande till mötes med bröd.
Ty de fly undan svärd, undan draget svärd, och undan spänd båge och undan krigets tunga.
Ty så har Herren sagt till mig: Om ett år, såsom dagakarlen räknar året, skall all Kedars härlighet vara förgången,
och föga skall då vara kvar av Kedars hjältars bågar, så många de äro.
Ty så har HERREN, Israels Gud, talat.
Utsaga om Synernas dal.
Vad är då på färde, eftersom allt ditt folk stiger upp på taken?
Du larmuppfyllda, du bullrande stad, du glada stad!
Dina slagna hava icke blivit slagna med svärd, ej dödats i strid.
Alla dina furstar hava samfällt flytt undan, utan bågskott blevo de fångar.
Ja, så många som påträffades hos dig blevo allasammans fångar, huru långt bort de än flydde.
Därför säger jag: Vänden blicken ifrån mig, jag måste gråta bitterligen; trugen icke på mig tröst för att dottern mitt folk har blivit förstörd.
Ty en dag med förvirring, nedtrampning och bestörtning kommer från Herren, HERREN Sebaot, i Synernas dal, med nedbrutna murar och med rop upp mot berget.
Elam hade fattat kogret, vagnskämpar och ryttare följde honom; Kir hade blottat skölden.
Dina skönaste dalar voro fyllda med vagnar, och ryttarna hade fattat stånd vid porten.
Juda blev blottat och låg utan skydd.
Då skådade du bort efter vapnen i Skogshuset.
Och I sågen att Davids stad hade många rämnor, och I samladen upp vattnet i Nedre dammen.
Husen i Jerusalem räknaden I, och I bröten ned husen för att befästa muren.
Och mellan de båda murarna gjorden I en behållare för vattnet från Gamla dammen.
Men I skådaden icke upp till honom som hade verkat detta; till honom som för länge sedan hade bestämt det sågen I icke.
Herren, HERREN Sebaot kallade eder på den dagen till gråt och klagan, till att raka edra huvuden och hölja eder i sorgdräkt.
Men i stället hängåven I eder åt fröjd och glädje; I dödaden oxar och slaktaden får, I åten kött och drucken vin, I saden: »Låtom oss äta och dricka, ty i morgon måste vi dö.»
Därför ljuder från HERREN Sebaot denna uppenbarelse i mina öron: Sannerligen, denna eder missgärning skall icke bliva försonad, så länge I leven, säger Herren, HERREN Sebaot.
Så sade Herren, HERREN Sebaot: Gå bort till honom där, förvaltaren, överhovmästaren Sebna, och säg till honom:
Vad gör du här, och vem tänker du lägga här, eftersom du här hugger ut en grav åt dig?
Du som hugger ut din grav så högt uppe, du som i klippan urholkar en boning åt dig,
du må veta att HERREN skall slunga dig långt bort, en sådan man som du är.
Han skall rulla dig tillhopa till en klump,
han skall hopnysta dig såsom ett nystan, och kasta dig såsom en boll bort till ett land som har utrymme nog för dig; där skall du dö, och dit skola dina härliga vagnar komma, du skamfläck för din herres hus.
Ja, jag skall stöta dig bort ifrån din plats, och från din tjänst skall du bliva avsatt.
Och på den dagen skall jag kalla på min tjänare Eljakim, Hilkias son;
honom skall jag ikläda din livklädnad, och med ditt bälte skall jag omgjorda honom, och skall lägga ditt välde i hans hand, så att han bliver en fader för Jerusalems invånare och för Juda hus.
Och jag skall giva honom Davids hus' nyckel att bära; när han upplåter, skall ingen tillsluta, och när han tillsluter, skall ingen upplåta.
Och jag skall slå in honom till en stadig spik i en fast vägg, och han skall bliva ett äresäte för sin faders hus.
Men om då hans faders hus, så tungt det är, hänger sig på honom, med ättlingar och avkomlingar -- alla slags småkärl av vad slag som helst, skålar eller allahanda krukor --
då, på den dagen, säger HERREN Sebaot, skall spiken, som var inslagen i den fasta väggen lossna; den skall gå sönder och falla ned, och bördan som hängde därpå, skall krossas.
Ty så har HERREN talat.
Utsaga om Tyrus.
Jämren eder, I Tarsis-skepp!
Ty det är ödelagt, utan hus och utan gäster; från kittéernas land når dem budskapet härom.
Sitten stumma, I kustlandets invånare!
Köpmän från Sidon, sjöfarande män, uppfyllde dig;
av Sihors säd och Nilflodens skördar skaffade du dig vinning, i det du for över stora vatten och drev handel därmed bland folken.
Men stå där nu med skam, du Sidon; ty så säger havet, havets fäste: »Så är jag då utan avkomma och har icke fött några barn, icke uppfött ynglingar, icke fostrat jungfrur.»
När man får höra detta i Egypten, då bävar man vid ryktet om Tyrus.
Dragen bort till Tarsis och jämren eder, I kustlandets invånare.
Är detta eder glada stad, hon den urgamla, som av sina fötter bars till fjärran land, för att gästa där?
Vem beslöt detta över Tyrus, henne som delade ut kronor, vilkens köpmän voro furstar, vilkens krämare voro stormän på jorden?
HERREN Sebaot var den som beslöt det, för att slå ned all den stolta härligheten och ödmjuka alla stormän på jorden.
Bred nu ut dig över ditt land såsom Nilfloden, du dotter Tarsis; du bär ingen boja mer.
Han räckte ut sin hand över havet, han kom konungariken att darra; HERREN bjöd om Kanaans fästen att de skulle ödeläggas.
Han sade: »Du skall ej allt framgent få leva i fröjd, du kränkta jungfru, du dotter Sidon.
Stå upp och drag bort till kittéernas land; dock, ej heller där får du ro.
Se, kaldéernas land, folket som förr ej var till, de vilkas land Assyrien gjorde till boning åt öknens djur, de resa där sina belägringstorn och omstörta stadens platser och göra den till en grushög.
Jämren eder, I Tarsis-skepp, ty edert fäste är förstört.»
På den tiden skall Tyrus ligga förgätet i sjuttio år, såsom rådde där alltjämt en och samma konung; men efter sjuttio år skall det gå med Tyrus, såsom det heter i visan om skökan:
»Tag din harpa och gå omkring i staden, du förgätna sköka; spela vackert och sjung flitigt, så att man kommer ihåg dig.»
Ty efter sjuttio år skall HERREN se till Tyrus, och det skall åter få begynna att taga emot skökolön och bedriva otukt med jordens alla konungariken i den vida världen.
Men hennes handelsförvärv och vad hon får såsom skökolön skall vara helgat åt HERREN; det skall icke läggas upp och icke gömmas, utan de som bo inför HERRENS ansikte skola av hennes handelsförvärv hava mat till fyllest och präktiga kläder.
Se, HERREN ödelägger jorden och föröder den; han omvälver, vad därpå är, och förströr dess inbyggare.
Och det går prästen såsom folket, husbonden såsom tjänaren, husfrun såsom tjänarinnan, säljaren såsom köparen, låntagaren såsom långivaren, gäldenären såsom borgenären.
Jorden bliver i grund ödelagd och i grund utplundrad; ty HERREN har talat detta ord.
Jorden sörjer och tvinar bort, jordkretsen försmäktar och tvinar bort, vad högt är bland jordens folk försmäktar.
Ty jorden har blivit ohelgad under sina inbyggare; de hava överträtt lagarna, de hava förvandlat rätten, brutit det eviga förbundet.
Därför uppfräter förbannelse jorden, och de som bo där måste lida, vad de hava förskyllt; därför förtäras jordens inbyggare av hetta, så att ej många människor finnas kvar.
Vinmusten sörjer, vinträdet försmäktar; de som voro så hjärteglada sucka nu alla.
Det är förbi med fröjden vid pukornas ljud, de gladas larm ha tystnat; det är förbi med fröjden vid harpans klang.
Vin dricker man icke mer under sång, rusdrycken kännes bitter för dem som dricka den.
Nedbruten ligger den öde staden; vart hus är stängt, så att ingen kommer därin.
Därute höres klagorop över vinet; all glädje är såsom en nedgången sol, all jordens fröjd har flyktat.
Ödeläggelse allenast är kvar i staden, och porten är slagen i spillror.
Ty det måste så gå på jorden bland folken, såsom det går, när man slår ned oliver, såsom när man gör en efterskörd, sedan vinbärgningen är slut.
Dessa häva då upp sin röst och jubla; fröjderop över HERRENS höghet ljuda borta i väster:
»Ären därför HERREN i österns bygder, även i havsländerna HERRENS, Israels Guds, namn.»
Från jordens ända höra vi lovsånger: »En härlig lott får den rättfärdige!»
Men jag säger: Jag arme, jag arme, ve mig!
Härjare härja, ja härjande fara härjare fram.
Faror, fallgropar och fällor vänta eder, I jordens inbyggare.
Och om någon flyr undan farlighetsropen, så störtar han i fallgropen, och om han kommer upp ur fallgropen, så fångas han i fällan.
Ty fönstren i höjden äro öppnade, och jordens grundvalar bäva.
Jorden brister, ja, den brister; jorden rämnar, ja, den rämnar; jorden vacklar, ja, den vacklar;
jorden raglar, ja, den raglar såsom en drucken; den gungar såsom vaktskjulet i trädets topp.
Dess överträdelse vilar tung på den, och den faller och kan icke mer stå upp.
På den tiden skall HERREN hemsöka höjdens här uppe i höjden och jordens konungar nere på jorden.
Och de skola samlas tillhopa, såsom fångar hopsamlas i fånggropen, och skola inneslutas i fängelse; sent omsider når dem hemsökelsen.
Då skall månen blygas och solen skämmas; ty HERREN Sebaot skall då vara konung på Sions berg och i Jerusalem, och hans äldste skola skåda härlighet.
HERRE, du är min Gud; jag vill upphöja dig, jag vill prisa ditt namn, ty du gör underfulla ting, du utför rådslut ifrån fordom tid, fasta och beståndande.
Ja, du har gjort staden till en stenhop, den befästa staden till en grushög; främlingarnas palats står ej mer där såsom en stad, aldrig skall det byggas upp igen.
Därför måste nu det vilda folket ära dig, den grymma hednastaden frukta dig.
Ty du har varit ett värn för den arme, ett värn för den fattige i hans nöd, en tillflykt mot störtskurar, ett skygd under hettan.
Ty våldsverkarnas raseri är likasom en störtskur mot en vägg.
Och såsom du kuvar hettan, när det är som torrast, så kuvar du främlingarnas larm; ja, såsom hettan dämpas genom molnens skugga, så dämpas de grymmas segersång.
Och HERREN Sebaot skall på detta berg göra ett gästabud för alla folk, ett gästabud med feta rätter, ett gästabud med starkt vin, ja, med feta, märgfulla rätter, med starkt vin, väl klarat.
Och han skall på detta berg göra om intet det dok som höljer alla folk, och det täckelse som betäcker alla folkslag.
Han skall för alltid göra döden om intet; och Herren, HERREN skall avtorka tårarna från alla ansikten, och skall taga bort sitt folks smälek överallt på jorden.
Ty så har HERREN talat.
På den tiden skall man säga: Se, där är vår Gud, som vi förbidade och som skulle frälsa oss.
Ja, där är HERREN, som vi förbidade; låtom oss fröjdas och vara glada över hans frälsning.
Ty HERRENS hand skall vila över detta berg, men Moab skall bliva nedtrampad i sitt eget land, likasom strå trampas ned i gödselpölen.
Och huru han än där breder ut sina händer, lik simmaren, när han simmar, så skall dock hans högmod bliva nedbrutet, trots hans händers alla konster.
Ja, dina murars höga fäste störtar han omkull och ödmjukar, han slår det till jorden, ned i stoftet.
På den tiden skall man sjunga denna sång i Juda land: »Vår stad giver oss styrka; murar och värn bereda oss frälsning.
Låten upp portarna, så att ett rättfärdigt folk får draga därin, ett som håller tro.
Den som är fast i sitt sinne bevarar du i frid, i frid; ty på dig förtröstar han.
Förtrösten då på HERREN till evig tid; ty HERREN, HERREN är en evig klippa.
Ty dem som trona i höjden, dem störtar han ned, ja, den höga staden; han ödmjukar den, ödmjukar den till jorden, han slår den ned i stoftet.
Den trampas under fötterna, under de förtrycktas fötter, under de armas steg.»
Men den rättfärdiges väg är jämn; åt den rättfärdige bereder du en jämnad stig.
Ja, på dina domars väg, HERRE, förbida vi dig; till ditt namn och ditt pris står vår själs trängtan.
Min själ trängtar efter dig om natten, och anden i mig söker dig bittida; ty när dina domar drabbar jorden, lära sig jordkretsens inbyggare rättfärdighet.
Om nåd bevisas mot den ogudaktige, så lär han sig icke rättfärdighet; i det land, där rätt skulle övas, gör han då vad orätt är och ser icke HERRENS höghet.
HERRE, din hand är upplyft, men de se det icke; må de nu med blygsel se din nitälskan för folket; ja, må eld förtära dina ovänner.
HERRE, du skall skaffa frid åt oss, ty allt vad vi hava uträttat har du utfört åt oss.
HERREN, vår Gud, andra herrar än du hava härskat över oss, men allenast dig prisa vi, allenast ditt namn.
De döda få icke liv igen, skuggorna stå ej åter upp; därför hemsökte och förgjorde du dem och utrotade all deras åminnelse.
Du förökade en gång folket, HERRE; du förökade folket och bevisade dig härlig; du utvidgade landets alla gränser.
HERRE, i nöden hava de nu sökt dig, de hava utgjutit tysta böner, när din tuktan kom över dem.
Såsom en havande kvinna, då hon är nära att föda, våndas och ropar i sina kval, så var det med oss inför ditt ansikte, o HERRE.
Vi voro också havande och våndades; men när vi födde, var det vind.
Vi kunde icke bereda frälsning åt landet; inga människor födas mer till att bo på jordens krets.
Men dina döda må få liv igen; mina dödas kroppar må åter stå upp.
Vaknen upp och jublen, I som liggen i graven; ty din dagg är en ljusets dagg, och jorden skall giva igen de avsomnade.
Välan då, mitt folk, gå in i dina kamrar och stäng igen dörrarna om dig; göm dig ett litet ögonblick, till dess att vreden har gått förbi.
Ty se, HERREN träder ut ur sin boning, för att hemsöka jordens inbyggare för deras missgärning; och jorden skall låta komma i dagen allt blod som där har blivit utgjutet, och skall icke längre betäcka dem som där hava blivit dräpta.
På den tiden skall HERREN med sitt svärd, det hårda, det stora och starka, hemsöka Leviatan, den snabba ormen, och Leviatan, den ringlande ormen, och skall dräpa draken, som ligger i havet.
På den tiden skall finnas en vingård, rik på vin, och man skall sjunga om den:
Jag, HERREN, är dess vaktar, åter och åter vattnar jag den.
För att ingen skall skada den, vaktar jag den natt och dag.
Jag vredgas icke på den; nej, om tistel och törne ville begynna strid, så skulle jag gå löst därpå och bränna upp alltsammans.
Eller ock måste man söka skydd hos mig och göra fred med mig; ja, fred måste man göra med mig.
I tider som komma skall Jakob skjuta rötter och Israel grönska och blomstra; jordkretsen skola de uppfylla med sin frukt.
Har man väl plågat dem så, som han plågade deras plågare?
Eller dräptes de så, som deras dräpta fiender blevo dräpta?
Nej, väl näpste han folket, när han förkastade och försköt det, väl ryckte han bort det med sin hårda vind, på östanstormens dag;
men därför kan ock Jakobs missgärning då bliva försonad och deras synds borttagande då giva fullmogen frukt, när alla stenar i deras altaren äro förstörda -- såsom då man krossar sönder kalkstycken -- och när Aseror och solstoder ej mer resas upp.
Se, den fasta staden ligger öde, den har blivit en folktom plats, övergiven såsom en öken, kalvar gå där i bet och lägra sig där och avbita de kvistar där finnas.
Och när grenarna äro torra, bryter man av dem, och kvinnor komma och göra upp eld med dem.
Ty detta är icke ett folk med förstånd; därför visar deras skapare dem intet förbarmande, och deras danare dem ingen misskund.
Och det skall ske på den tiden att HERREN anställer en inbärgning, från den strida floden intill Egyptens bäck; och I skolen varda insamlade, en och en, I Israels barn.
Och det skall ske på den tiden att man stöter i en stor basun; och de som hava varit borttappade i Assyriens land och fördrivna till Egyptens land, de skola då komma; och de skola tillbedja HERREN på det heliga berget i Jerusalem.
Ve dig, du Efraims druckna mäns stolta krona, du hans strålande härlighets vissnande blomster på bergshjässan ovan de vinberusades bördiga dal!
Se, från Herren kommer en som är stark och väldig, lik en hagelskur, en förödande storm, lik en störtskur med väldiga, översvämmande vatten, som slår allt till jorden med mat.
Under fötterna bliver den då trampad, Efraims druckna mäns stolta krona.
Och det går med hans strålande härlighets vissnande blomma på bergshjässan ovan den bördiga dalen, såsom det går med ett fikon därnere, ett som har mognat före sommarskörden: så snart någon får syn därpå, slukar han det, medan han ännu har det i sin hand.
På den tiden skall HERREN Sebaot bliva en härlig krona och en strålande krans för kvarlevan av sitt folk;
och han skall bliva en rättens ande för den som skipar rätt, och en starkhetsmakt för dem som driva fienden på porten.
Men också här raglar man av vin, stapplar man av starka drycker; både präster och profeter ragla av starka drycker, de äro överlastade av vin, de stappla av starka drycker; de ragla, när de profetera, de vackla, när de skipa rätt.
Ja, alla bord äro fulla av vämjeliga spyor, ingen ren fläck finnes.
-- »Vem är det då han vill lära förstånd, och vem skall han få att giva akt på sin predikan?
Äro vi då nyss avvanda från modersmjölken, nyss tagna från modersbröstet?
Det är ju gnat på gnat, gnat på gnat, prat på prat, prat på prat, litet här, litet där!»
-- Ja väl, genom stammande läppar och på ett främmande tungomål skall han tala till detta folk,
han som en gång sade till dem: »Här är vilostaden, låten den trötte få vila; här är vederkvickelsens ort.»
Men sådant ville de icke höra.
Så skall då HERRENS ord bliva för dem »gnat på gnat, gnat på gnat, prat på prat, prat på prat, litet här, litet där».
Och så skola de, bäst de gå där, falla baklänges och krossas, varda snärjda och fångade.
Hören därför HERRENS ord, I bespottare, I som råden över folket här i Jerusalem.
Eftersom I sägen: »Vi hava slutit ett förbund med döden, med dödsriket hava vi ingått ett fördrag; om ock gisslet far fram likt en översvämmande flod, skall det icke nå oss, ty vi hava gjort lögnen till vår tillflykt och falskheten till vårt beskärm»,
därför säger Herren, HERREN så: Se, jag har lagt i Sion en grundsten, en beprövad sten, en dyrbar hörnsten, fast grundad; den som tror på den behöver icke fly.
Och jag skall låta rätten vara mätsnöret och rättfärdigheten sänklodet.
Och hagel skall slå ned eder lögntillflykt, och vatten skall skölja bort edert beskärm.
Och edert förbund med döden skall bliva utplånat, och edert fördrag med dödsriket skall icke bestå; när gisslet far fram likt en översvämmande flod, då solen I varda nedtrampade.
Så ofta det far fram, skall det träffa eder; ty morgon efter morgon skall det fara fram, ja, både dag och natt.
Idel förskräckelse bliver det, när I måsten akta på den predikan.
Ty sängen bliver då för kort att sträcka ut sig på och täcket för knappt att svepa in sig i.
Ty HERREN skall stå upp likasom på Perasims berg, och han skall låta se sin vrede likasom i Gibeons dal.
Han skall utföra sitt verk, ett sällsamt verk; han skall förrätta sitt arbete, ett förunderligt arbete.
Så hören nu upp med eder bespottelse, för att edra band ej må bliva än hårdare; ty om förstöring och oryggligt besluten straffdom över hela jorden har jag hört från Herren, HERREN Sebaot.
Lyssnen och hören min röst, akten härpå och hören mitt tal.
När åkermannen vill så, plöjer han då beständigt och hackar upp och harvar sin mark?
Nej, fastmer: sedan han har jämnat fältet, strör han ju där svartkummin och kastar dit kryddkummin och sår vete i rader och korn på dess särskilda plats och spält i kanten.
Ty hans Gud har undervisat honom och lärt honom det rätta sättet.
Man tröskar ju ej heller svartkummin med tröskvagn och låter ej vagnshjul gå över kryddkummin, utan klappar ut svartkummin med stav och kryddkummin med käpp.
Och brödsäden, tröskar man sönder den?
Nej, man plägar icke oavlåtligt tröska den och driva sina vagnshjul och hästar däröver; man vill ju icke tröska sönder den.
Också detta kommer från HERREN Sebaot; han är underbar i råd och stor i vishet.
Ve dig, Ariel, Ariel, du stad, där David slog upp sitt läger!
Läggen år till år och låten högtiderna fullborda sitt kretslopp,
så skall jag bringa Ariel i trångmål; jämmer skall följa på jämmer, och då bliver det för mig ett verkligt Ariel.
Jag skall slå läger runt omkring dig och omsluta dig med vallar och resa upp bålverk emot dig.
Då skall du tala djupt nedifrån jorden, och dina ord skola dämpade komma fram ur stoftet; din röst skall höras såsom en andes ur jorden, och ur stoftet skall du viska fram dina ord.
Men främlingshopen skall bliva såsom fint damm och våldsverkarhopen såsom bortflyende agnar; plötsligt och med hast skall detta ske.
Från HERREN Sebaot skall hemsökelsen komma, med tordön och jordbävning och stort dunder, med storm och oväder och med lågor av förtärande eld.
Och hela hopen av alla de folk som drogo i strid mot Ariel, de skola vara såsom en drömsyn om natten, alla som drogo i strid mot det och dess borg och bragte det i trångmål.
Såsom när den hungrige drömmer att han äter, men vaknar och känner sin buk vara tom, och såsom när den törstande drömmer att han dricker, men vaknar och känner sig törstig och försmäktande, så skall det gå med hela hopen av alla de folk som drogo i strid mot Sions berg.
Stån där med häpnad, ja, varen häpna; stirren eder blinda, ja, varen blinda, I som ären druckna, men icke av vin, I som raglen, men icke av starka drycker.
Ty HERREN har utgjutit över eder en tung sömns ande och har tillslutit edra ögon; han har höljt mörker över profeterna och över siarna, edra ledare.
Och så har profetsynen om allt detta blivit för eder lik orden i en förseglad bok: om man räcker en sådan åt någon som kan läsa och säger: »Läs detta», så svarar han: »Jag kan det icke, den är ju förseglad»,
och om man räcker den åt någon som icke kan läsa och säger: »Läs detta», så svarar han: »Jag kan icke läsa.»
Och HERREN har sagt: Eftersom detta folk nalkas mig med sin mun och ärar mig med sina läppar, men låter sitt hjärta vara långt ifrån mig, så att deras fruktan för mig består i inlärda människobud,
därför skall jag ännu en gång göra underbara ting mot detta folk, ja, underbara och förunderliga; de visas vishet skall förgås, och de förståndigas förstånd skall bliva förmörkat.
Ve eder, I som söken att dölja edra rådslag för HERREN i djupet, och som bedriven edra verk i mörkret, I som sägen: »Vem ser oss, och vem känner oss?»
Huru förvända ären I icke!
Skall då leret aktas lika med krukmakaren?
Skall verket säga om sin mästare: »Han har icke gjort mig»?
Eller skall bilden säga om honom som har format den: »Han förstår intet»?
Se, ännu allenast en liten tid, och Libanon skall förvandlas till ett bördigt fält och det bördiga fältet räknas såsom vildmark.
De döva skola på den tiden höra vad som läses för de, och de blindas ögon skola se och vara fria ifrån dunkel och mörker;
och de ödmjuka skola då känna allt större glädje i HERREN; och de fattigaste bland människor skola fröjda sig i Israels Helige.
Ty våldsverkarna äro då icke mer till, bespottarna hava fått en ände, och de som stodo efter fördärv äro alla utrotade,
de som genom sitt tal gjorde att oskyldiga blevo fällda och snärjde den som skulle skipa rätt i porten och genom lögn vrängde rätten för den rättfärdige.
Därför säger HERREN så till Jakobs hus, han som förlossade Abraham: Nu skall Jakob icke mer behöva blygas, nu skall hans ansikte ej vidare blekna;
ty när han -- hans barn -- få se mina händer verk ibland sig, då skola de hålla mitt namn heligt, de skola hålla Jakobs Helige helig och förskräckas för Israels Gud.
De förvillade skola då få förstånd, och de knorrande skola taga emot lärdom.
Ve eder, I vanartiga barn, säger HERREN, I som gören upp rådslag som icke komma från mig, och sluten förbund, utan att min Ande är med, så att I därigenom hopen synd på synd,
I som dragen ned till Egypten, utan att hava rådfrågat min mun, för att söka eder ett värn hos Farao och en tillflykt under Egyptens skugga!
Se, Faraos värn skall bliva eder till skam, och tillflykten under Egyptens skugga skall bliva eder till blygd.
Ty om ock hans furstar äro i Soan, och om än hans sändebud komma ända till Hanes,
så skall dock var man få blygas över detta folk, som icke kan hjälpa dem, icke vara till bistånd och hjälp, utan allenast till skam och smälek.
Utsaga om Söderlandets odjur.
Genom ett farornas och ångestens land, där lejoninnor och lejon hava sitt tillhåll, jämte huggormar och flygande drakar, där föra de på åsnors ryggar sina rikedomar och på kamelers pucklar sina skatter till ett folk som icke kan hjälpa dem.
Ty Egyptens bistånd är fåfänglighet och tomhet; därför kallar jag det landet »Rahab, som ingenting uträttar».
Så gå nu in och skriv detta på en tavla, som må förvaras bland dem, och teckna upp det i en bok, så att det bevaras för kommande dagar, alltid och evinnerligen.
Ty det är ett gensträvigt folk, trolösa barn, barn som icke vilja höra HERRENS lag,
utan säga till siarna: »Upphören med edra syner», och till profeterna: »Profeteren icke för oss vad sant är; talen till oss sådant som är oss välbehagligt, profeteren bedrägliga ting;
viken av ifrån vägen, gån åt sidan från stigen, skaffen bort ur vår åsyn Israel Helige.»
Därför säger Israels Helige så: »Eftersom I förakten detta ord och förtrösten på våld och vrånghet och stödjen eder på sådant,
därför skall denna missgärning bliva för eder såsom ett fallfärdigt stycke på en hög mur, vilket mer och mer giver sig ut, till dess att muren plötsligt och med hast störtar ned och krossas;
den krossa, såsom när man våldsamt slår en lerkruka i bitar, så våldsamt att man bland bitarna icke kan finna en skärva stor nog att därmed taga eld från eldstaden eller ösa upp vatten ur dammen.»
Ty så säger Herren, HERREN, Israels Helige: »Om i vänden om och ären stilla, skolen I bliva frälsta, genom stillhet och förtröstan varden I starka.»
Men i viljen icke.
I sägen: »Nej, på hästar vilja vi jaga fram» -- därför skolen I också bliva jagade; »på snabba springare vilja vi rida åstad» -- därför skola ock edra förföljare vara snabba.
Tusen av eder skola fly för en enda mans hot eller för fem mäns hot, till dess att vad som är kvar av eder bliver såsom en ensam stång på bergets topp, såsom ett baner på höjden.
Ja, därför väntar HERREN, till dess att han kan vara eder nådig; därför tronar han i höghet, till dess att han kan förbarma sig över eder.
Ty en domens Gud är HERREN; saliga äro alla de som vänta efter honom.
Ja, du folk som bor på Sion, i Jerusalem, ingalunda må du gråta.
Han skall förvisso vara dig nådig, när du ropar; så snart han hör din röst, skall han svara dig.
Ty väl skall Herren giva eder nödens bröd och fångenskapens dryck, men sedan skola dina lärare icke mer sättas å sido, utan dina ögon skola se upp till dina lärare.
Och om du viker av, vare sig åt höger eller åt vänster, så skola dina öron höra detta ord ljuda bakom dig; »Här är vägen, vandren på en.»
Då skolen I akta för orent silvret varmed edra skurna beläten äro överdragna, och guldet varmed edra gjutna beläten äro belagda; du skall kasta ut det såsom orenlighet och säga till det: »Bort härifrån!»
Och han skall giva regn åt säden som du har sått på din mark, och han skall av markens gröda giva dig bröd som är kraftigt och närande; och din boskap skall på den tiden gå i bet på vida ängar.
Och oxarna och åsnorna med vilka man brukar jorden, de skola äta saltad blandsäd om man har kastat med vanna och kastskovel.
Och på alla höga berg och alla stora höjder skola bäckar rinna upp med strömmande vatten -- när den stora slaktningens dag kommer, då torn skola falla.
Och månens ljus skall bliva såsom solens ljus, och solens ljus skall varda sju gånger klarare, såsom ett sjufaldigt dagsljus, när den tid kommer, då HERREN förbinder sitt folks skador och helar såren efter slagen som det har fått.
Se, HERRENS namn kommer fjärran ifrån, med brinnande vrede och med tunga rökmoln; hans läppar äro fulla av förgrymmelse, och hans tunga är såsom förtärande eld;
hans andedräkt är lik en ström som svämmar över, så att den når ändå upp till halsen.
Ty han vill sålla folken i förintelsens såll och lägga i folkslagens mun ett betsel, till att leda dem vilse.
Då skolen I sjunga såsom i en natt då man firar helig högtid, och edra hjärtan skola glädja sig, såsom när man under flöjters ljud tågar upp på HERRENS berg, upp till Israels klippa.
Och HERREN skall låta höra sin röst i majestät och visa huru hans arm drabbar, i vredesförgrymmelse och med förtärande eldslåga, med storm och störtskurar och hagelstenar.
Ty för HERRENS röst skall Assur bliva förfärad, när han slår honom med sitt ris.
Och så ofta staven far fram och HERREN efter sitt rådslut låter den falla på honom skola pukor och harpor ljuda.
Gång på gång skall han lyfta sin arm till att strida mot honom.
Ty en Tofetplats är längesedan tillredd, ja ock för konungen är den gjord redo, och djup och vid är den; dess rund är fylld av eld och av ved i myckenhet, och lik en svavelström skall HERRENS Ande sätta den i brand.
Ve dem som draga åstad ned till Egypten för att få hjälp, i det de förlita sig på hästar, dem som sätta sin förtröstan på vagnar, därför att där finnas så många, och på ryttare, därför att mängden är så stor, men som ej vända sin blick till Israels Helige och icke fråga efter HERREN!
Också han är ju vis; han låter olyckan komma, och han ryggar icke sina ord.
Han reser sig upp mot de ondas hus och mot den hjälp som ogärningsmännen sända.
Ty egyptierna äro människor och äro icke Gud, deras hästar äro kött och icke ande.
Och HERREN skall räcka ut sin hand, och då skall hjälparen vackla och den hjälpte falla, och båda skola tillhopa förgås.
Ty så har HERREN sagt till mig: Såsom ett lejon ryter, ett ungt lejon över sitt rov, och icke skrämmes bort av herdarnas rop eller rädes för deras larm, när de i mängd samlas dit, så skall HERREN Sebaot fara ned för att strida på Sions berg och uppe på dess höjd.
Såsom fågeln breder ut sina vingar, så skall HERREN Sebaot beskärma Jerusalem; han skall beskärma och hjälpa, han skall skona och rädda.
Så vänden nu om till honom, från vilken I haven avfallit genom ett så djupt fall, I Israels barn.
Ty på den tiden skall var och en av eder kasta bort de avgudar av silver och de avgudar av guld, som edra händer hava gjort åt eder till synd.
Och Assur skall falla, men icke för en mans svärd; ett svärd, som icke är en människas, skall förtära honom.
Han skall fly för svärd, och hans unga män skola bliva trälar.
Och hans klippa skall förgås av skräck, och hans furstar skola i förfäran fly ifrån baneret.
Så säger HERREN, han som har sin eld på Sion och sin ugn i Jerusalem.
En konung skall uppstå, som skall regera med rättfärdighet, och härskare, som skola härska med rättvisa.
Var och en av dem skall vara såsom en tillflykt i stormen, ett skydd mot störtskuren; de skola vara såsom vattenbäckar i en ödemark, såsom skuggan av en väldig klippa i ett törstigt land.
Då skola de seendes ögon icke vara förblindade, och de hörandes öron skola lyssna till.
Då skola de lättsinnigas hjärtan bliva förståndiga och vinna kunskap, och de stammandes tungor skola tala flytande och tydligt.
Dåren skall då icke mer heta ädling, ej heller bedragaren kallas herre.
Ty en dåre talar dårskap, och hans hjärta reder till fördärv; så övar han gudlöshet och talar, vad förvänt är, om HERREN, så låter han den hungrige svälta och nekar den törstige en dryck vatten.
Och bedragaren brukar onda vapen, han tänker ut skändliga anslag till att fördärva de betryckta genom lögnaktiga ord, fördärva en fattig, som har rätt i sin talan.
Men en ädling tänker ädla tankar och står fast vid det som ädelt är.
I kvinnor, som ären så säkra, stån upp och hören min röst; I sorglösa jungfrur, lyssnen till mitt tal.
När år och dagar hava gått, då skolen I darra, I som ären så sorglösa, ty då är det slut med all vinbärgning, och ingen fruktskörd kommer mer.
Bäven, I som ären så säkra, darren, I som ären så sorglösa, läggen av edra kläder och blotten eder, kläden edra länder med säcktyg.
Slån eder för bröstet och klagen över de sköna fälten, över de fruktsamma vinträden,
över mitt folks åkrar som fyllas av törne och tistel, ja, över alla glädjens boningar i den yra staden.
Ty palatsen äro övergivna, den folkrika staden ligger öde, Ofelhöjden med vakttornet är förvandlad till grotthålor för evig tid, till en plats, där vildåsnor hava sin fröjd och där hjordar beta --
detta intill dess att ande från höjden bliver utgjuten över oss.
Då skall öknen bliva ett bördigt fält och det bördiga fältet räknas såsom vildmark;
då skall rätten taga sin boning i öknen och rättfärdigheten bo på det bördiga fältet.
Och rättfärdighetens frukt skall vara frid och rättfärdighetens vinning vara ro med trygghet till evig tid.
Och mitt folk skall bo i fridshyddor, i trygga boningar och på säkra viloplatser.
Men under hagelskurar skall skogen fällas, och djupt skall staden bliva ödmjukad.
Sälla ären då I som fån så vid alla vatten, I som kunnen låta edra oxar och åsnor fritt ströva omkring.
Ve dig, du fördärvare, som själv har gått fri ifrån fördärvet!
Ve dig, du härjare, som själv har undgått förhärjning!
När du har fyllt ditt mått att fördärva, drabbas du själv av fördärvet; när du har fullbordat till härjande drabbas du själv av förhärjning.
HERRE, var oss nådig, dig förbida vi.
Var dessas arm var morgon; ja, var vår frälsning i nödens tid.
För ditt väldiga dån fly folken bort; när du reser dig upp, förskingras folkslagen.
Och man får skövla och taga byte efter eder, såsom gräsmaskar skövla; såsom gräshoppor störta fram, så störtar man över det.
HERREN är hög, ty han bor i höjden; han uppfyller Sion med rätt och rättfärdighet.
Ja, trygga tider skola komma för dig!
Vishet och kunskap bereda Sion frälsning i rikt mått, och HERRENS fruktan skall vara deras skatt.
Hör, deras hjältar klaga därute, fredsbudbärarna gråta bitterligen.
Vägarna äro öde, ingen går mer på stigarna.
Han bryter förbund, han aktar städer ringa, människor räknar han för intet.
Landet ligger sörjande och försmäktar, Libanon blyges och står förvissnat, Saron har blivit likt en hedmark, Basans och Karmels skogar fälla sina löv.
Men nu vill jag stå upp, säger HERREN, nu vill jag resa mig upp, nu vill jag upphäva mig.
Med halm gån I havande, och strå föden I; edert raseri är en eld, som skall förtära eder själva.
Folken skola förbrännas och bliva till aska, ja, likna avhugget törne, som brinner upp i eld.
Så hören nu, I som fjärran ärer, vad jag har gjort; förnimmen min makt, I som nära ären.
Syndarna i Sion bliva förskräckta, bävan griper de gudlösa. »Vem av oss kan härda ut vid en förtärande eld, vem av oss kan bo vid en evig glöd?»
Den som vandrar i rättfärdighet och talar, vad rätt är, den som föraktar, vad som vinnes genom orätt och våld, och den som avhåller sina händer från att taga mutor, den som tillstoppar sina öron för att icke höra om blodsgärningar och tillsluter sina ögon för att icke se, vad ont är,
han skall bo på höjderna, klippfästen skola vara hans värn, sitt bröd skall han få, och vatten skall han hava beständigt.
Ja, dina ögon skola skåda en konung i hans härlighet, de skola blicka ut över ett vidsträckt land.
Då skall ditt hjärta tänka tillbaka på förskräckelsens tid: »Var är nu skatteräknaren, var är nu skattevägaren, var är den som räknade tornen?»
Du slipper då att se det fräcka folket, folket, vars obegripliga språk man ej kunde förstå, vars stammande tungomål ingen kunde tyda.
Men skåda på Sion, våra högtiders stad, låt dina ögon betrakta Jerusalem: det är en säker boning, ett tält, som icke flyttas bort, ett vars pluggar aldrig ryckas upp och av vars streck intet enda brister sönder.
Ja, vi hava där HERREN, den väldige; han är för oss såsom floder och breda strömmar; ingen roddflotta kommer där fram, och det väldigaste skepp kan ej fara däröver.
Ty HERREN är vår domare, HERREN är vår härskare, HERREN är vår konung, han frälsar oss.
Dina tåg hänga slappa, de hålla ej masten stadig, ej seglet spänt.
Men då skall rövat gods utskiftas i myckenhet, ja, också de lama skola då taga byte.
Och ingen av invånarna skall säga: »Jag är svag», ty folket, som där bor, har fått sin missgärning förlåten.
Träden fram, I folk, och hören; I folkslag, akten härpå.
Jorden höre och allt vad på den är, jordens krets och vad som alstras därav.
Ty HERREN är förtörnad på alla folk och vred på all deras här; han giver dem till spillo, han överlämnar dem till att slaktas.
Deras slagna kämpar ligga bortkastade, och stank stiger upp från deras döda kroppar, och bergen flyta av deras blod.
Himmelens hela härskara förgås, och himmelen själv hoprullas såsom en bokrulle; hela dess härskara faller förvissnad ned, lik vissnade löv från vinrankan, lik vissnade blad ifrån fikonträdet.
Ty mitt svärd har druckit sig rusigt i himmelen; se, det far ned på Edom till dom, på det folk jag har givit till spillo.
Ja, ett svärd har HERREN, det dryper av blod och är dränkt i fett, i lamms och bockars blod, i fett ifrån vädurars njurar; ty HERREN anställer ett offer i Bosra, ett stort slaktande i Edoms land.
Vildoxar fällas ock därvid, tjurar, både små och stora.
Deras land dricker sig rusigt av blod, och deras jord bliver dränkt i fett.
Ty detta är en HERRENS hämndedag, ett vedergällningens år, då han utför Sions sak.
Då bliva Edoms bäckar förvandlade till tjära och dess jord till svavel; ja, dess land bliver förbytt i brinnande tjära.
Varken natt eller dag skall den branden slockna, evinnerligen skall röken därav stiga upp.
Från släkte till släkte skall landet ligga öde, aldrig i evighet skall någon gå där fram.
Pelikaner och rördrommar skola taga det i besittning, uvar och korpar skola bo däri; ty förödelsens mätsnöre och förstörelsens murlod skall han låta komma däröver.
Av dess ädlingar skola inga finnas kvar där, som kunna utropa någon till konung; och alla dess furstar få en ände.
Dess palatser fyllas av törne, nässlor och tistlar växa i dess fästen; och det bliver en boning för ökenhundar och ett tillhåll för strutsar.
Schakaler bo där tillsammans med andra ökendjur, och gastar ropa där till varandra; ja, där kan Lilit få ro, där kan hon finna en vilostad.
Där reder pilormen sitt bo och lägger sina ägg och kläcker så ut ynglet och samlar det i sitt skygd; ja, där komma gamarna tillhopa, den ene möter där den andre.
Söken efter i HERRENS bok och läsen däri; icke ett enda av de djuren skall utebliva, det ena skall icke fåfängt söka det andra.
Ty det är hans mun, som bjuder det, det är hans Ande, som samlar dem tillhopa.
Det är han, som kastar lott för dem, hans hand tillskiftar dem deras mark efter mätsnöre; till evig tid skola de hava den till besittning, från släkte till släkte bo därpå.
Öknen och ödemarken skola glädja sig, och hedmarken skall fröjdas och blomstra såsom en lilja.
Den skall blomstra skönt och fröjda sig, ja, fröjda sig och jubla; Libanons härlighet skall bliva den given, Karmels och Sarons prakt.
Ja, de skola få se HERRENS härlighet, vår Guds prakt.
Stärken maktlösa händer, given kraft åt vacklande knän.
Sägen till de försagda: »Varen frimodiga, frukten icke.»
Se, eder Gud kommer med hämnd; vedergällning kommer från Gud, ja, själv kommer han och frälsar eder.
Då skola de blindas ögon öppnas och de dövas öron upplåtas.
Då skall den lame hoppa såsom en hjort, och den stummes tunga skall jubla.
Ty vatten skola bryta fram i öknen och strömmar på hedmarken.
Av förbränt land skall bliva en sjö och av torr mark vattenkällor; på den plats, där ökenhundar lägrade sig, skall växa gräs jämte vass och rör.
Och en banad väg, en farväg, skall gå där fram, och den skall kallas »den heliga vägen»; ingen oren skall färdas därpå, den skall vara för dem själva.
Den som vandrar den vägen skall icke gå vilse, om han ock hör till de fåkunniga.
Där skall icke vara något lejon, ej heller skall något annat vilddjur komma dit.
Intet sådant skall finnas där, men ett frälsat folk skall vandra på den.
Ja, HERRENS förlossade skola vända tillbaka och komma till Sion med jubel; evig glädje skall kröna deras huvuden, fröjd och glädje skola de undfå, men sorg och suckan skola fly bort.
Och i konung Hiskias fjortonde regeringsår hände sig, att Sanherib, konungen i Assyrien, drog upp och angrep alla befästa städer i Juda och intog dem.
Och konungen i Assyrien sände från Lakis åstad Rab-Sake med en stor här till Jerusalem mot konung Hiskia; och han stannade vid Övre dammens vattenledning, på vägen till Valkarfältet.
Då gingo överhovmästaren Eljakim, Hilkias son, och sekreteraren Sebna och kansleren Joa, Asafs son, ut till honom.
Och Rab-Sake sade till dem: »Sägen till Hiskia: Så säger den store konungen, konungen i Assyrien: Vad är det för en förtröstan, som du nu har hängivit dig åt?
Jag säger: Det är allenast munväder, att du vet råd och har makt att föra kriget.
På vem förtröstar du då, eftersom du har satt dig upp mot mig?
Du förtröstar väl på den bräckta rörstaven Egypten, men se, när någon stöder sig på den, går den i i hans hand och genomborrar den.
Ty sådan är Farao, konungen i Egypten, för alla som förtrösta på honom.
Eller säger du kanhända till mig: 'Vi förtrösta på HERREN, vår Gud?'
Var det då icke hans offerhöjder och altaren Hiskia avskaffade, när han sade till Juda och Jerusalem: 'Inför detta altare skolen I tillbedja'?
Men ingå nu ett vad med min herre, konungen i Assyrien: jag vill giva dig två tusen hästar, om du kan skaffa dig ryttare till dem.
Huru skulle du då kunna slå tillbaka en enda ståthållare, en av min herres ringaste tjänare?
Och du sätter din förtröstan till Egypten i hopp om att så få vagnar och ryttare!
Menar du då att jag utan HERRENS vilja har dragit upp till detta land för att fördärva det?
Nej, det är HERREN, som har sagt till mig: Drag upp mot detta land och fördärva det.»
Då sade Eljakim och Sebna och Joa till Rab-Sake: »Tala till dina tjänare på arameiska, ty vi förstå det språket, och tala icke till oss på judiska inför folket som står på muren.»
Men Rab-Sake svarade: »Är det då till din herre och till dig, som min herre har sänt mig att tala dessa ord?
Är det icke fastmer till de män som sitta på muren och som jämte eder skola nödgas äta sin egen träck och dricka sitt eget vatten?»
Därefter trädde Rab-Sake närmare och ropade med hög röst på judiska och sade: »Hören den store konungens, den assyriske konungens, ord.
Så säger konungen: Låten icke Hiskia bedraga eder, ty han förmår icke rädda eder.
Och låten icke Hiskia förleda eder att förtrösta på HERREN, därmed att han säger: 'HERREN skall förvisso rädda oss; denna stad skall icke bliva given i den assyriske konungens hand.'
Hören icke på Hiskia.
Ty så säger konungen i Assyrien: Gören upp i godo med mig och given eder åt mig, så skolen I få äta var och en av sitt vinträd och av sitt fikonträd och dricka var och en ur sin brunn,
till dess jag kommer och hämtar eder till ett land som är likt edert eget land, ett land med säd och vin, ett land med bröd och vingårdar.
Låten icke Hiskia förleda eder, när han säger: 'HERREN skall rädda oss.'
Har väl någon av de andra folkens gudar räddat sitt land ur den assyriske konungens hand?
Var äro Hamats och Arpads gudar?
Var äro Sefarvaims gudar?
Eller hava de räddat Samaria ur min hand?
Vilken bland dessa länders alla gudar har väl räddat sitt land ur min hand, eftersom I menen, att HERREN skall rädda Jerusalem ur min hand?»
Men de tego och svarade honom icke ett ord, ty konungen hade så bjudit och sagt: »Svaren honom icke.»
Och överhovmästaren Eljakim, Hilkias son, och sekreteraren Sebna och kansleren Joa, Asafs son, kommo till Hiskia med sönderrivna kläder och berättade för honom, vad Rab-Sake hade sagt.
Då nu konung Hiskia hörde detta, rev han sönder sina kläder och höljde sig i sorgdräkt och gick in i HERRENS hus.
Och överhovmästaren Eljakim och sekreteraren Sebna och de äldste bland prästerna sände han, höljda i sorgdräkt, till profeten Jesaja, Amos' son.
Och de sade till denne: »Så säger Hiskia: En nödens, tuktans och smälekens dag är denne dag, ty fostren hava väl kommit fram till födseln, men kraft att föda finnes icke.
Kanhända skall HERREN, din Gud, höra Rab-Sakes ord, med vilka hans herre, konungen i Assyrien, har sänt honom till att smäda den levande Guden, så att han straffar honom för dessa ord som han, HERREN, din Gud, har hört.
Så bed nu en bön för den kvarleva som ännu finnes.»
När nu konung Hiskias tjänare kommo till Jesaja,
sade Jesaja till dem: »Så skolen I säga till eder herre: Så säger HERREN: Frukta icke för de ord som du har hört, dem, med vilka den assyriske konungens tjänare hava hädat mig.
Se, jag skall låta en sådan ande komma in i honom, att han på grund av ett rykte som han skall få höra vänder tillbaka till sitt land; och jag skall låta honom falla för svärd i hans eget land.»
Och Rab-Sake vände tillbaka och fann den assyriske konungen upptagen med att belägra Libna; ty han hade hört, att han hade brutit upp från Lakis.
Men när Sanherib fick höra sägas om Tirhaka, konungen i Etiopien, att denne hade dragit ut för att strida mot honom, skickade han, så snart han hörde detta, sändebud till Hiskia och sade:
»Så skolen I säga till Hiskia, Juda konung: Låt icke din Gud, som du förtröstar på, bedraga dig, i det att du tänker: 'Jerusalem skall icke bliva givet i den assyriske konungens hand.'
Du har ju hört, vad konungarna i Assyrien hava gjort med alla andra länder, huru de hava givit dem till spillo.
Och du skulle nu bliva räddad!
Hava väl de folk, som mina fäder fördärvade, Gosan, Haran, Resef och Edens barn i Telassar, blivit räddade av sina gudar?
Var är Hamats konung och Arpads konung och konungen över Sefarvaims stad, över Hena och Iva?»
När Hiskia hade mottagit brevet av sändebuden och läst det, gick han upp i HERRENS hus, och där bredde Hiskia ut det inför HERRENS ansikte.
Och Hiskia bad till HERREN och sade:
»HERRE Sebaot, Israels Gud, du som tronar på keruberna, du allena är Gud, den som råder över alla riken på jorden; du har gjort himmel och jord.
HERRE, böj ditt öra härtill och hör; HERRE, öppna dina ögon och se.
Ja, hör alla Sanheribs ord, det budskap, varmed han har smädat den levande Guden.
Det är sant, HERRE, att konungarna i Assyrien hava förött alla länder såsom ock sitt eget land.
Och de hava kastat deras gudar i elden; ty dessa voro inga gudar, utan verk av människohänder, trä och sten; därför kunde de förgöra dem.
Men fräls oss nu, HERRE, vår Gud, ur hans hand, så att alla riken på jorden förnimma, att du, HERRE, är den ende.»
Då sände Jesaja, Amos' son, bud till Hiskia och lät säga: »Så säger HERREN, Israels Gud, jag, till vilken du har bett angående Sanherib, konungen i Assyrien:
Detta är det ord, som HERREN har talat om honom: Hon föraktar dig och bespottar dig, jungfrun dottern Sion; hon skakar huvudet efter dig, dottern Jerusalem.
Vem har du smädat och hädat, och mot vem har du upphävt din röst?
Alltför högt har du upplyft dina ögon -- ja, mot Israels Helige.
Genom dina tjänare smädade du HERREN, när du sade: 'Med mina många vagnar drog jag upp på bergens höjder, längst upp på Libanon; jag högg ned dess höga cedrar och väldiga cypresser; jag trängde fram till dess översta höjder, dess frodigaste skog;
jag grävde brunnar och drack ut vatten, och med min fot uttorkade jag alla Egyptens strömmar.'
Har du icke hört, att jag för länge sedan beredde detta?
Av ålder bestämde jag ju så; och nu har jag fört det fram: du fick makt att ödelägga befästa städer till grusade stenhopar.
Deras invånare blevo maktlösa, de förfärades och stodo med skam.
Det gick dem såsom gräset på marken och gröna örter, såsom det som växer på taken, och säd, som förgås, förrän strået har vuxit upp.
Om du sitter eller går ut eller går in, så vet jag det, och huru du rasar mot mig.
Men då du nu så rasar mot mig och då ditt övermod har nått till mina öron, skall jag sätta min krok i din näsa och mitt betsel i din mun och föra dig tillbaka samma väg, som du har kommit på.
Och detta skall för dig vara tecknet: man skall detta år äta, vad som växer upp av spillsäd, och nästa år självvuxen säd, men det tredje året skolen I få så och skörda och plantera vingårdar och äta deras frukt.
Och den räddade skaran av Juda hus, som bliver kvar, skall åter skjuta rot nedtill och bära frukt upptill.
Ty från Jerusalem skall utgå en kvarleva, en räddad skara från Sions berg.
HERREN Sebaots nitälskan skall göra detta.
Därför säger HERREN så om konungen i Assyrien: Han skall icke komma in i denna stad och icke skjuta någon pil ditin; han skall icke mot den föra fram någon sköld eller kasta upp någon vall mot den.
Samma väg han kom skall han vända tillbaka, och in i denna stad skall han icke komma, säger HERREN.
Ty jag skall beskärma och frälsa denna stad för min tjänare Davids skull.»
Och HERRENS ängel gick ut och slog i assyriernas läger ett hundra åttiofem tusen man; och när man bittida följande morgon kom ut, fick man se döda kroppar ligga där överallt.
Då bröt Sanherib, konungen i Assyrien, upp och tågade tillbaka; och han stannade sedan i Nineve.
Men när han en gång tillbad i sin gud Nisroks tempel, blev han dräpt med svärd av sina söner Adrammelek och Sareser; därefter flydde dessa undan till Ararats land.
Och hans son Esarhaddon blev konung efter honom.
Vid den tiden blev Hiskia dödssjuk; och profeten Jesaja, Amos' son, kom till honom och sade till honom: »Så säger HERREN: Beställ om ditt hus; ty du måste dö och skall icke tillfriskna.»
Då vände Hiskia sitt ansikte mot väggen och bad till HERREN.
Och han sade: »Ack HERRE, tänk dock på huru jag har vandrat inför dig i trohet och med hängivet hjärta och gjort, vad gott är i dina ögon.»
Och Hiskia grät bitterligen.
Då kom HERRENS ord till Jesaja: han sade:
»Gå och säg till Hiskia: Så säger HERREN, din fader Davids Gud: Jag har hört din bön, jag har sett dina tårar.
Se, jag skall föröka din livstid med femton år;
jag skall ock rädda dig och denna stad ur den assyriske konungens hand.
Ja, jag skall beskärma denna stad.
Och detta skall för dig vara tecknet från HERREN därpå att HERREN skall göra, vad han nu har lovat:
se, solvisarskuggan, som nu på Ahas' solvisare har gått nedåt med solen, skall jag låta gå tio steg tillbaka.»
Så gick solen tillbaka på solvisaren de tio steg, som den reda hade lagt till rygga.
En sång, skriven av Hiskia, Juda konung, när han hade varit sjuk och tillfrisknat från sin sjukdom:
Jag tänkte: Jag går hädan i mina bästa dagar, in genom dödsrikets portar; jag varder berövad återstoden av mina år.
Jag tänkte: Jag får icke mer se HERREN, HERREN i de levandes land.
Hos dem som bo i förgängelsens rike får jag ej mer skåda människor.
Min hydda ryckes upp och flyttas bort ifrån mig såsom en herdes tält.
Jag har vävt mitt liv till slut såsom en vävare sin väv, och jag skäres nu ned från bommen; innan dagen har gått över till natt, är du färdig med mig.
Jag måste ryta såsom ett lejon intill morgonen; så krossas alla bin i min kropp.
Ja, innan dagen har gått över till natt, är du färdig med mig.
Jag klagade såsom en svala, såsom en trana, jag suckade såsom en duva; matta blickade mina ögon mot höjden: »HERRE, jag lider nöd; tag dig an min sak.»
Men vad skall jag väl säga, då han nu har talat till mig och själv utfört sitt verk?
I ro får jag nu leva alla mina år till slut efter all min själs bedrövelse.
Herre, sådant länder till liv, min ande har i allo sitt liv därav.
Och så helar du mig -- ja, giv mig liv!
Se till mitt bästa kom denna bittra bedrövelse över mig.
I din kärlek räddade du min själ ifrån förintelsens grop, i det du kastade alla mina synder bakom din rygg.
Ty dödsriket tackar dig icke, döden prisar dig icke, och de som hava farit ned i graven hoppas ej mer på din trofasthet.
De som leva, de som leva, de tacka dig, såsom ock jag nu gör; och fäderna göra din trofasthet kunnig för barnen.
HERREN skall frälsa mig, och mina sånger skola vi då spela i alla våra livsdagar däruppe i HERRENS hus.
Och Jesaja tillsade, att man skulle taga en fikonkaka och lägga den såsom plåster på bulnaden, så skulle han tillfriskna.
Men Hiskia sade: »Vad för ett tecken gives mig därpå att jag skall få gå upp i HERRENS hus?»
Vid samma tid sände Merodak-Baladan, Baladans son, konungen i Babel, brev och skänker till Hiskia; och han fick höra, att denne hade varit sjuk, men blivit återställd.
Och Hiskia gladde sig över deras ankomst och visade dem sitt förrådshus, sitt silver och guld, sina välluktande kryddor och sina dyrbara oljor och hela sitt tyghus och allt vad som fanns i hans skattkamrar.
Intet fanns i Hiskias hus eller eljest i hans ägo, som han icke visade dem.
Men profeten Jesaja kom till konung Hiskia och sade till honom: »Vad hava dessa män sagt, och varifrån hava de kommit till dig?»
Hiskia svarade: »De hava kommit till mig ifrån fjärran land, ifrån Babel.»
Han sade vidare: »Vad hava de sett i ditt hus?»
Hiskia svarade: »Allt som är i mitt hus hava de sett: intet finnes i mina skattkamrar, som jag icke har visat dem.»
Då sade Jesaja till Hiskia: »Hör HERREN Sebaots ord:
Se, dagar skola komma, då allt som finnes i ditt hus och som dina fäder hava samlat ända till denna dag skall föras bort till Babel; intet skall bliva kvar, säger HERREN.
Och söner till dig, de som skola utgå av dig och som du skall föda, dem skall man taga, och de skola bliva hovtjänare i den babyloniske konungens palats.»
Hiskia sade till Jesaja: »Gott är det HERRENS ord, som du har talat.»
Och han sade ytterligare: »Frid och trygghet skola ju få råda i min tid.»
Trösten, trösten mitt folk, säger eder Gud.
Talen ljuvligt till Jerusalem och prediken för det, att dess vedermöda är slut, att dess missgärning är försonad och att det har fått dubbelt igen av HERRENS hand för all sina synder.
Hör, man ropar; »Bereden väg för HERREN i öknen, banen på hedmarken en jämn väg för vår Gud.
Alla dalar skola höjas och alla berg och höjder sänkas; vad ojämnt är skall jämnas, och vad oländigt är skall bliva slät mark.
HERRENS härlighet skall varda uppenbarad, och allt kött skall tillsammans se den.
Ty så har HERRENS mun talat.»
Hör, någon talar: »Predika!», och en annan svarar: »Vad skall jag predika?» »Allt kött är gräs och all dess härlighet såsom ett blomster på marken.
Gräset torkar bort, blomstret förvissnar, när HERRENS andedräkt blåser därpå.
Gräset torkar bort, blomstret förvissnar, men vår Guds ord förbliver evinnerligen.»
Stig upp på ett högt berg, Sion, du glädjens budbärarinna; häv upp din röst med kraft, Jerusalem, du glädjens budbärarinna: häv upp den utan fruktan, säg till Juda stöder: »Se, där är eder Gud!»
Ja, Herren, HERREN kommer med väldighet, och hans arm visar sin makt.
Se, han har med sig sin lön, och hans segerbyte går framför honom.
Han för sin hjord i bet såsom en herde, han samlar lammen i sin famn och bär dem i sitt sköte och sakta för han moderfåren fram.
Vem är det, som mäter upp havens vatten i sin hand och märker ut himmelens vidd med sina utspända fingrar?
Vem mäter upp stoftet på jorden med ett tredingsmått?
Vem väger bergen på en våg och höjderna på en viktskål?
Vem kan utrannsaka HERRENS Ande, och vem kan giva honom råd och undervisa honom?
Går han till råds med någon, för att denne skall giva honom förstånd och lära honom den rätta stigen, lära honom kunskap och visa honom förståndets väg?
Nej, folken äro att akta såsom en droppe ur ämbaret och såsom ett grand på vågskålen; se, havsländerna lyfter han såsom ett stoftkorn.
Libanons skog vore icke nog till offerved och dess djur icke nog till brännoffer.
Folken äro allasammans såsom ett intet inför honom; såsom alls intet och idel tomhet aktas de av honom.
Vid vem viljen I då likna Gud, och vad finnes honom likt att ställa vid hans sida?
Månne ett avgudabeläte? -- det gjutes av någon konstnär, och guldsmeden överdrager det sedan med guld, och med silverkedjor pryder så guldsmeden det.
Den som icke har råd att offra så mycket, han väljer ut ett stycke trä, som icke ruttnar, och söker sig en förfaren konstnär, som kan förfärdiga ett beläte, som ej faller omkull.
Haven I då intet förstånd?
Hören I då intet?
Blev detta icke förkunnat för eder från begynnelsen?
Haven I icke förstått, vad jordens grundvalar säga?
Han är den som tronar över jordens rund, och dess inbyggare äro såsom gräshoppor; han är den som utbreder himmelen såsom ett flor och spänner ut den såsom ett tält att bo inunder.
Han är den som gör furstarna till intet, förvandlar domarna på jorden till idel tomhet.
Knappt äro de planterade, knappt äro de sådda, knappt har deras stam slagit rot i jorden, så blåser han på dem, och de förtorka, och en stormvind för dem bort såsom strå.
Vid vem viljen I då likna mig, så agg jag skulle vara såsom han? säger den Helige.
Lyften upp edra ögon mot höjden och sen: vem har skapat allt detta?
Det har han som för härskaran däruppe fram i räknade hopar; han nämner dem alla vid namn.
Så stor är hans makt, så väldig hans kraft, att icke en enda utebliver.
Huru kan du säga sådant, du Jakob, och tala så, du Israel: »Min väg är fördold för HERREN, och min rätt är försvunnen för min Gud»?
Vet du då icke, har du ej hört det, att HERREN är en evig Gud, han som har skapat jordens ändar?
Han bliver ej trött och uppgives icke, hans förstånd är outrannsakligt.
Han giver den trötte kraft och förökar den maktlöses styrka.
Ynglingar kunna bliva trötta och uppgivas, och unga män kunna falla;
men de som bida efter HERREN hämta ny kraft, de få nya vingfjädrar såsom örnarna.
Så hasta de åstad utan att uppgivas, de färdas framåt utan att bliva trötta.
Tigen, I havsländer, och lyssnen till mig, och må folken hämta ny kraft; må de så komma fram och tala, ja, låt oss med varandra träda inför rätta.
Vem har i öster låtit denne uppstå, som mötes av seger, var han går fram?
Vem giver folkslag i hans våld och gör honom till härskare över konungar?
Vem gör deras svärd till stoft och deras bågar till strå som föres bort av vinden?
Han förjagar dem, där han går lyckosam fram, vanliga vägar trampar icke hans fot.
Vem har verkat och utfört detta?
Det har han som från begynnelsen kallade människors släkten fram: jag, HERREN, som är den förste och som intill det sista är densamme.
Havsländerna se det och frukta, och jordens ändar förskräckas.
Man närmar sig till varandra och kommer tillhopa.
Den ene vill hjälpa den andre; han säger till den andre: »Fatta mod!»
Träsnidaren sätter mod i guldsmeden, bleckslagaren i den som hamrar på städ.
Han säger om lödningen: »Den är god» och fäster bilden med spikar, så att den ej faller omkull.
Men du Israel, min tjänare, du Jakob, som jag har utvalt, du ättling av Abraham, min vän,
du som jag har hämtat från jordens ändar och kallat hit från dess yttersta hörn och till vilken jag har sagt: »Du är min tjänare, dig har jag utvalt och icke försmått»,
frukta icke, ty jag är med dig; var ej försagd, ty jag är din Gud.
Jag styrker dig, jag hjälper dig ock, jag uppehåller dig med min rättfärdighets högra hand.
Se, alla som äro dig hätska skola komma på skam och blygas; dina motståndare skola bliva till intet och skola förgås.
Du skall söka efter dina vedersakare, men icke finna dem; ja, de som strida mot dig skola bliva till intet och få en ände.
Ty jag är HERREN, din Gud, som håller dig vid din högra hand och som säger till dig: Frukta icke, jag hjälper dig.
Så frukta nu icke, du mask Jakob, du Israels lilla hop.
Jag hjälper dig, säger HERREN; din förlossare är Israels Helige.
Se, jag gör dig till en tröskvagn, ny och med skarpa taggar, så att du skall söndertröska berg och krossa dem till stoft och göra höjder lika agnar.
Du skall kasta dem med kastskovel, och vinden skall föra dem bort och stormen förskingra dem; men du själv skall fröjda dig i HERREN och berömma dig av Israels Helige.
De betryckta och fattiga söka förgäves efter vatten, deras tunga försmäktar av törst; men jag, HERREN, skall bönhöra dem, jag, Israels Gud, skall icke övergiva dem.
Jag skall låta strömmar rinna upp på höjderna och källor i dalarna; jag skall göra öknen till en vattenrik sjö och torrt land till källsprång.
Och jag skall låta cedrar och akacieträd växa upp i öknen jämte myrten och olivträd och skall på hedmarken plantera cypress tillsammans med alm och buxbom,
för att man skall både se och veta och akta på och förstå, att HERRENS hand har gjort detta, att Israels Helige har skapat det.
Så träden nu fram med eder sak, säger HERREN; kommen med edra bevis, säger Jakobs konung.
Ja, må man komma med dem och förkunna för oss, vad som skall ske.
Var äro edra forna utsagor?
Läggen fram dem, för att vi må akta på dem och se till, huru de hava gått i fullbordan.
Eller låten oss höra, vad som nu skall komma,
förkunnen, vad framdeles skall hända, för att vi må se, att I ären gudar.
Ja, gören någonting, vad det nu vara må, så att vi alla häpna, när vi se det.
Men se, I ären ett intet, och edert verk är alls intet; den som utväljer eder är en styggelse.
Jag lät i norr en man uppstå, och han kom, ja, i öster en som skulle åkalla mitt namn; och han skulle gå fram över landsherrarna, såsom vore de lerjord, lik en krukmakare, som trampar lera.
Vem förkunnade detta förut, så att vi fingo veta det, eller i förväg, så att vi kunde säga: »Du hade rätt»?
Ingen fanns, som förkunnade det, ingen, som lät oss höra det, ingen, som hörde eder tala därom.
Jag är den förste, som säger till Sion: »Se, se där äro de», den förste, som bringar Jerusalem detta glädjens budskap.
Jag ser mig om, men här finnes ingen, ingen bland dessa, som kan giva besked; ingen som kan giva ett svar på min fråga.
Se, de äro allasammans fåfänglighet, deras verk äro ett intet, deras beläten vind och tomhet.
Se, över min tjänare som jag uppehåller, min utkorade, till vilken min själ har behag, över honom har jag låtit min Ande komma; han skall utbreda rätten bland folken.
Han skall icke skria eller ropa och icke låta höra sin röst på gatorna.
Ett brutet rör skall han icke sönderkrossa, och en tynande veke skall han icke utsläcka; han skall i trofasthet utbreda rätten.
Hans kraft skall icke förtyna eller brytas, intill dess att han har grundat rätten på jorden; havsländerna vänta efter hans lag.
Så säger Gud, HERREN, han som har skapat himmelen och utspänt den, han som har utbrett jorden med vad som alstras därav, han som har givit liv åt folket som är därpå och ande åt dem som vandra där:
Jag, HERREN, har kallat dig i rättfärdighet, och jag vill fatta dig vid handen och bevara dig och fullborda i dig förbundet med folket och sätta dig till ett ljus för folkslagen,
för att du må öppna blinda ögon och föra fångar ut ur fängelset, ja, ur fångenskapen dem som sitta i mörkret.
Jag, HERREN, det är mitt namn; och jag giver icke min ära åt någon annan eller mitt lov åt belätena.
Se, vad jag förut förkunnade, det har nu kommit.
Nu förkunnar jag nya ting; förrän de visa sig, låter jag eder höra om dem.
Sjungen till HERRENS ära en ny sång, hans lov från jordens ända, I som faren på havet, så ock allt vad däri är, I havsländer med edra inbyggare;
stämmen upp, du öken med dina städer och I byar, där Kedar bor; jublen, I klippornas invånare, ropen från bergens toppar.
Given HERREN ära och förkunnen hans lov i havsländerna.
HERREN drager ut såsom en hjälte, han eggar upp sig till iver såsom en krigare; han uppgiver härskri, han ropar högt och visar sin makt mot sina fiender.
I lång tid har jag tegat, jag höll mig stilla och betvang mig; men nu skall jag höja rop såsom en barnaföderska, jag vill skaffa mig luft och andas ut.
Jag skall föröda berg och höjder och låta allt gräs på dem förtorka; jag skall göra strömmar till land och låta allt gräs på dem förtorka; jag skall göra strömmar till land och låta sjöar torka ut.
Och de blinda skall jag leda på en väg som de icke känna; på stigar som de icke känna skall jag föra dem.
Jag skall göra mörkret framför dem till ljus och det som är ojämnt till jämn mark.
Detta är, vad jag skall göra, och jag skall ej rygga mitt ord.
Men de som förtrösta på skurna beläten och som säga till gjutna beläten: »I ären våra gudar», de skola vika tillbaka och stå där med skam.
Hören, I döve; I blinde, skåden och sen.
Vem är blind, om icke min tjänare, och så döv som den budbärare jag sänder åstad?
Du har fått se mycket, men du aktar icke därpå; fastän öronen hava blivit öppnade, lyssnar ingen till.
Det är HERRENS behag, för hans rättfärdighets skull, att han vill låta sin lag komma till makt och ära.
Men detta är ett plundrat och skövlat folk; dess ynglingar äro alla lagda i bojor, och i fängelser hållas de gömda, de hava blivit givna till plundring, och ingen finnes, som räddar, till skövling, och ingen säger: »Giv tillbaka.»
Ack att någon bland eder ville lyssna härtill, för framtiden giva akt och höra härpå!
Vem har lämnat Jakob till skövling och Israel i plundrares våld?
Har icke HERREN gjort det; han, mot vilken vi hava syndat, han, på vilkens vägar man icke ville vandra och på vilkens lag man icke ville höra?
Därför utgöt han över dem i sin vrede förtörnelse och krigets raseri.
Och de förbrändes därav runt omkring, men besinnade det icke; de förtärdes därav, men aktade icke därpå.
Men nu säger HERREN så, han som har skapat dig, Jakob, han som har danat dig, Israel: Frukta icke, ty jag har förlossat dig, jag har kallat dig vid ditt namn, du är min.
Om du ock måste gå genom vatten, så är jag med dig, eller genom strömmar, så skola de icke fördränka dig; måste du än gå genom eld, så skall du ej bliva svedd, och lågorna skola ej förtära dig.
Ty jag är HERREN, din Gud, Israels Helige, din frälsare; jag giver Egypten till lösepenning för dig, Etiopien och Seba i ditt ställe.
Eftersom du är så dyrbar i mina ögon, så högt aktad och så älskad av mig, därför giver jag människor till lösen för dig och folk till lösen för ditt liv.
Frukta då icke, ty jag är med dig.
Jag skall låta dina barn komma från öster, och från väster skall jag samla dig tillhopa.
Jag skall säga till Norden: »Giv hit» och till södern: »Förhåll mig dem icke; för hit mina söner ifrån fjärran och mina döttrar ifrån jordens ända,
envar som är uppkallad efter mitt namn och som jag har skapat till min ära, envar som jag har danat och gjort.»
För hitut det blinda folket, som dock har ögon, och de döva, som dock hava öron.
Alla folk hava kommit tillsammans, folkslagen samla sig tillhopa.
Vem bland dem finnes, som skulle kunna förutsäga sådant?
Må de låta oss höra sina forna utsagor.
Må de ställa fram sina vittnen och bevisa sin rätt, så att dessa, när de höra det, kunna säga: »Det är sant.»
Men I ären mina vittnen, säger HERREN, I ären min tjänare, den som jag har utvalt, på det att I mån veta och tro mig och förstå, att det är jag; före mig är ingen Gud danad, och efter mig skall ingen komma.
Jag, jag är HERREN, och förutom mig finnes ingen frälsare.
Jag har förkunnat det och skaffat frälsning, jag har kungjort det och ingen främmande gud bland eder.
I ären mina vittnen, säger HERREN; och jag är Gud.
Ja, allt framgent är jag densamme, och ingen kan rädda från min hand.
När jag vill göra något, vem kan då avvända det?
Så säger HERREN, eder förlossare, Israels Helige: För eder skull sänder jag mitt bud mot Babel, och jag skall driva dem allasammans på flykten, jag skall driva kaldéerna ned på skeppen som voro deras fröjd.
Jag är HERREN, eder Helige, Israels skapare, eder konung.
Så säger HERREN, han som gör en väg i havet, en stig i väldiga vatten,
han som för vagnar och hästar ditut, ja, härskara och och stridsmakt, sedan ligga de där tillhopa och kunna icke stå upp, de äro utsläckta, de hava slocknat såsom en veke:
Tänken icke på vad förr har varit, akten icke på vad fordom har skett.
Se, jag vill göra något nytt.
Redan nu visar det sig; märken I det icke?
Ja, jag skall göra en väg i öknen och strömmar i ödemarken,
så att markens djur skola ära mig, schakaler och strutsar, därför att jag låter vatten flyta i öknen, strömmar i ödemarken, så att mitt folk, min utkorade, kan få dricka.
Det folk, som jag har danat åt mig, skall förtälja mitt lov.
Men icke har du, Jakob, kallat mig hit, i det du har gjort dig möda för min skull, du Israel.
Icke har du framburit åt mig dina brännoffersfår eller ärat mig med dina slaktoffer; icke har jag vållat dig arbete med spisoffer, ej heller möda med rökelse.
Icke har du köpt kalmus åt mig för dina penningar eller mättat mig med dina slaktoffers fett.
Nej, du har vållat mig arbete genom dina synder och möda genom dina missgärningar.
Jag, jag är den som utplånar dina överträdelser för min egen skull, och dina synder kommer jag icke mer ihåg.
Låt mig höra, vad du har att säga, och låt oss gå till rätta med varandra; tala du, för att du må finnas rättfärdig.
Men se, redan din stamfader syndade, och de som förde din talan begingo överträdelser mot mig.
Därför har jag måst låta helgedomens furstar utstå vanära och har överlämnat Jakob åt tillspillogivning, Israel åt försmädelse.
Men hör nu, du Jakob, min tjänare, du Israel, som jag har utvalt.
Så säger HERREN, han som har skapat dig, han som danade dig redan i moderlivet och som hjälper dig: Frukta icke, du min tjänare Jakob, du Jesurun, som jag har utvalt.
Ty jag skall utgjuta vatten över de törstiga och strömmar över det torra; jag skall utgjuta min Ande över din barn och min välsignelse över dina telningar,
så att de växa upp mitt ibland gräset såsom pilträd vid vattenbäckar.
Då skall den ene säga: »HERREN tillhör jag», och den andre skall åberopa Jakobs namn, och en tredje skall skriva på sin hand: »HERRENS egen» och skall bruka Israel såsom ett ärenamn.
Så säger HERREN, Israels konung, och hans förlossare, HERREN Sebaot: Jag är den förste, och jag är den siste, och förutom mig finnes ingen Gud.
Och vem talar, såsom jag har gjort, alltsedan jag lät urtidsfolket framträda?
Må han förkunna det och lägga det fram för mig.
Ja, må de förkunna det tillkommande, vad som skall ske.
Frukten icke och varen icke förskräckta.
Har jag icke för länge sedan låtit dig höra om detta och förkunnat det?
I ären ju mina vittnen.
Finnes väl någon Gud förutom mig?
Nej, ingen annan klippa finnes, jag vet av ingen.
Avgudamakarna äro allasammans idel tomhet, och deras kära gudar kunna icke hjälpa.
Deras bekännare se själva intet och förstå intet; därför måste de ock komma på skam.
Om någon formar en gud och gjuter ett beläte, så är det honom till intet gagn.
Se, hela dess följe skall komma på skam; konstnärerna själva äro ju allenast människor.
Må de församlas, så många de äro, och träda fram; de skola då alla tillhopa med förskräckelse komma på skam.
Smeden tager sitt verktyg och bearbetar sitt smide i glöden, han formar det med hammare, han bearbetar det med kraftig arm; till äventyrs får han därvid svälta, så att han bliver vanmäktig, och försaka att dricka, så att han bliver matt.
Träsnidaren spänner ut sitt mätsnöre och gör märken på trästycket med sitt ritstift, han arbetar därpå med sina eggjärn och märker ut det med passaren; och han gör så därav en mansbild, en prydlig människogestalt, som får bo i ett hus.
Man fäller åt sig cedrar; man tager plantor av stenek och vanlig ek och uppdrager dem åt sig bland skogens träd; man planterar åt sig lärkträd, och regnet giver dem växt.
Detta hava människorna till bränsle; och man tager därav och värmer sig därmed, man tänder på det och bakar bröd därvid.
Men därjämte förfärdigar man en gud därav och tillbeder den, man gör därav ett beläte och faller ned för det.
En del av träet bränner man alltså upp i eld, över en annan del därav tillagar man kött till att äta, steker sin stek och äter sig mätt; när man så har värmt sig, säger man: »Gott, nu är jag varm, nu njuter jag av brasan.»
Men av det som är kvar gör man en gud, man gör sig ett beläte, och för det faller man ned och tillbeder, man bönfaller inför det och säger: »Rädda mig, ty du är min gud.» --
Ja, sådana veta intet och förstå intet, ty igentäppta äro deras ögon, så att de icke se, och deras hjärtan, så att de intet begripa.
Ingen har så mycken eftertanke, så mycket vett eller förstånd, att han säger: »En del därav har jag bränt upp i eld, och på kolen har jag bakat bröd och stekt kött och har så ätit; skulle jag då av återstoden göra en styggelse?
Skulle jag falla ned för ett stycke trä?»
Den som så håller sig till vad som blott är aska, han är förledd av ett dårat hjärta, så att han icke förstår att rädda sin själ, icke att tänka: »Blott fåfänglighet är, vad jag håller i min högra hand.»
Tänk härpå, du Jakob, du Israel, ty du är min tjänare; jag har danat dig, ja, du är min tjänare.
Israel, du varder icke förgäten av mig.
Jag utplånar dina överträdelser såsom ett moln och dina synder såsom en sky.
Vänd om till mig, ty jag förlossar dig.
Jublen, I himlar, ty HERREN utför sitt verk; höjen glädjerop, I jordens djup, bristen ut i jubel, I berg, du skog med alla dina träd; ty HERREN förlossar Jakob, han bevisar sig härlig i Israel.
Så säger HERREN, din förlossare, han som danade dig redan i moderlivet: »Jag, HERREN, är den som för allt, den som ensam utspänner himmelen och utan någons hjälp breder ut jorden.
Jag är den som gör lögnprofeternas tecken om intet och gör spåmännen till dårar, den som låter de vise komma till korta och gör deras klokhet till dårskap,
men som låter sin tjänares ord bliva beståndande och fullbordar sina sändebuds rådslag.
Jag är den som säger om Jerusalem: »Det skall bliva bebott» och om Juda städer: »De skola varda uppbyggda; jag skall upprätta ruinerna där.»
Jag är den som säger till havsdjupet: »Sina ut; dina strömmar vill jag låta uttorka.»
Jag är den som säger om Kores: »Han är min herde, han skall fullborda all min vilja, och han skall säga om Jerusalem: 'Det skall bliva uppbyggt' och till templet: 'Din grund skall åter varda lagd.'»
Så säger HERREN till sin smorde, till Kores som jag har fattat vid hans högra hand, då jag nu vill slå ned folken inför honom och lösa svärdet från konungarnas länd, då jag vill öppna dörrarna för honom så att inga portar mer äro stängda:
Själv skall jag gå framför dig, backarna skall jag jämna ut; kopparportarna skall jag krossa, och järnbommarna skall jag bryta sönder.
Och jag skall giva dig dolda skatter och bortgömda rikedomar, för att du må förnimma, att jag, HERREN, är den som har kallat dig vid ditt namn, jag, Israels Gud.
För min tjänare Jakobs skull, för Israels, min utkorades, skull kallade jag dig vid ditt namn och gav dig ärenamn, innan du kände mig.
Jag är HERREN och eljest ingen, utom mig finnes ingen Gud; innan du kände mig, omgjordade jag dig,
för att man skulle förnimma både i öster och i väster, att alls ingen finnes förutom mig, att jag är HERREN och eljest ingen,
jag som danar ljuset och skapar mörkret, jag som giver lyckan och skapar olyckan.
Jag, HERREN, är den som gör allt detta.
Drypen, I himlar därovan, och må skyarna låta rättfärdighet strömma ned.
Må jorden öppna sig, och må dess frukt bliva frälsning; rättfärdighet låte den ock växa upp.
Jag, HERREN, skapar detta.
Ve dig som vill gå till rätta med din Skapare, ja, ve dig, du skärva bland andra skärvor av jord!
Skall väl leret säga till krukmakaren: »Vad kan du göra?»
Och skall ditt verk säga om dig: »Han har inga händer»?
Ve dig som säger till din fader: »Icke kan du avla barn» och till hans hustru: »Icke kan du föda barn»!
Så säger HERREN, Israels Helige, som ock är hans skapare: Frågen mig om det tillkommande; lämnen åt mig omsorgen om mina söner, mina händer verk.
Det är jag, som har gjort jorden och skapat människorna därpå; det är mina händer, som hava utspänt himmelen, och hela dess härskara har jag bådat upp.
Det är ock jag, som har låtit denne uppstå i rättfärdighet, och alla hans vägar skall jag göra jämna.
Han skall bygga upp min stad och släppa mina fångar lösa, och det icke för betalning eller för gåvor, säger HERREN Sebaot.
Så säger HERREN: Vad egyptierna hava förvärvat med sitt arbete och etiopiernas och Sebas resliga folk med sin handel, det skall allt övergå i din hand och höra dig till.
De skola följa bakom dig, i kedjor skola de gå.
Och de skola falla ned inför dig och ställa sin bön till dig: »Allenast i dig är Gud, och eljest finnes ingen, alls ingen annan Gud.»
Ja, du är sannerligen en outgrundlig Gud, du Israels Gud, du frälsare
De komma alla på skam och varda till blygd, de måste allasammans gå där med blygd, alla avgudamakarna.
Men Israel bliver frälst genom HERREN med en evig frälsning; aldrig i evighet skolen I komma på skam och varda till blygd.
Ty så säger HERREN, han som har skapat himmelen, han som är Gud, han som har danat jorden och gjort den, han som har berett den och som icke har skapat den till att vara öde, utan danat den till att bebos: Jag är HERREN och eljest ingen.
Jag har icke talat i det fördolda, någonstädes i ett mörkt land; jag har icke sagt till Jakobs släkt: Förgäves skolen I söka mig.
Jag är HERREN, som talar sanning, som förkunnar, vad rätt är.
Så församlen eder nu och kommen hit, träden fram allasammans, I räddade, som ären kvar av folken.
Ty de hava intet förstånd, de som föra sina träbeläten omkring i högtidståg och bedja till en gud som icke kan frälsa.
Förkunnen något och läggen fram det; alla tillhopa må rådslå därom.
Vem har långt förut låtit eder höra detta och för länge sedan förkunnat det?
Har icke jag, HERREN, gjort det jag, förutom vilken ingen Gud mer finnes, ingen Gud, som är rättfärdig och som frälsar, nej, ingen finnes jämte mig.
Vänden eder till mig, så varden I frälsta, I jordens alla ändar; ty jag är Gud och eljest ingen.
Jag har svurit vid mig själv, från min mun har utgått ett sanningsord, ett ord, som icke skall ryggas: För mig skola alla knän böja sig, och mig skola alla tungor giva sin ed.
Så har man betygat om mig: Allenast hos HERREN finnes rättfärdighet och makt.
Till honom skola komma med blygd alla de som hava varit honom hätska.
Ja, genom HERREN får all Israels släkt sin rätt, och av honom skola de berömma sig.
Bel sjunker ned, Nebo måste böja sig, deras bilder lämnas åt djur och fänad; de som I förden omkring i högtidståg, de lastas nu på ök som bära sig trötta av bördan.
Ja, de måste båda böja sig och sjunka ned; de kunna icke rädda någon börda, själva vandra de bort i fångenskap.
Så hören nu på mig, I av Jakobs hus, I alla som ären kvar av Israels hus, I som haven varit lastade på mig allt ifrån moderlivet och burna av mig allt ifrån modersskötet.
Ända till eder ålderdom är jag densamme, och intill dess I varden grå, skall jag bära eder; så har jag hittills gjort, och jag skall också framgent hålla eder uppe, jag skall bära och rädda eder.
Med vem viljen I likna och jämföra mig, och med vem viljen I sammanställa mig, så att jag skulle vara honom lik?
Man skakar ut guld ur pungen och väger upp silver på vågen, och så lejer man en guldsmed att göra det till en gud, för vilken man kan falla ned och tillbedja.
Den lyfter man på axeln och bär den bort och sätter ned den på dess plats, för att den skall stå där och ej vika från stället.
Men ropar någon till den, så svarar den icke och frälsar honom icke ur hans nöd.
Tänken härpå och kommen till förnuft; besinnen eder, I överträdare.
Tänken på vad förr var, redan i forntiden; ty jag är Gud och eljest ingen, en Gud, vilkens like icke finnes;
jag som i förväg förkunnar, vad komma skall, och långt förut, vad ännu ej har skett; jag som säger: »Mitt rådslut skall gå i fullbordan, och allt vad jag vill, det gör jag»;
jag som kallar på örnen från öster och ifrån fjärran land på mitt rådsluts man.
Vad jag har bestämt, det sätter jag ock i verket.
Så hören nu på mig, I stormodige, I som menen, att hjälpen är långt borta.
Se, jag låter min hjälp nalkas, den är ej långt borta, och min frälsning dröjer icke; jag giver frälsning i Sion och min härlighet åt Israel.
Stig ned och sätt dig i stoftet, du jungfru dotter Babel, sätt dig på jorden utan tron, du kaldéernas dotter; ty man skall icke mer kalla dig »den bortklemade och yppiga».
Tag till kvarnen och mal mjöl, lägg av din slöja, lyft upp släpet, blotta benet, vada genom strömmarna.
Din blygd skall varda blottad, och din skam skall ses.
Hämnd skall jag utkräva och ej skona någon människa.
Vår förlossares namn är HERREN Sebaot, Israels Helige!
Sitt tyst och drag dig undan i mörkret, du kaldéernas dotter; ty du skall icke mer bliva kallad »konungarikenas drottning».
Jag förtörnades på mitt folk, jag ohelgade min arvedel och gav dem i din hand.
Och du visade dem intet förbarmande; på gamla män lät du ditt ok tynga hårt.
Du tänkte: »Jag skall evinnerligen förbliva en drottning» därför ville du ej akta på och tänkte ej på änden.
Så hör nu detta, du som lever i vällust, du som tronar så trygg, du som säger i ditt hjärta: »Jag och ingen annan; aldrig skall jag sitta såsom änka, aldrig veta av, vad barnlöshet är.»
Se, båda dessa olyckor skola komma över dig med hast, på en och samma dag: både barnlöshet och änkestånd skola komma över dig i fullaste mått, trots myckenheten av dina trolldomskonster, trots dina besvärjelsers starka kraft.
Du kände dig trygg i din ondska, du tänkte: »Ingen ser mig.»
Din vishet och din kunskap var det, som förförde dig, så att du så sade i ditt hjärta: »Jag och ingen annan.»
Därför skall en olycka komma över dig, som du ej förmår besvärja bort, och ett fördärv skall falla över dig, som du icke skall kunna avvända; ja, plötsligt skall ödeläggelse komma över dig, när du minst anar det.
Träd fram med de besvärjelser och många trolldomskonster som du har mödat dig med från din ungdom; se till, om du så kan skaffa hjälp, om du så kan skrämma bort faran.
Du har arbetat dig trött med dina många rådslag.
Må de nu träda fram, må de frälsa dig, dessa som avmäta himmelen och spana i stjärnorna och var nymånad kungöra, varifrån ditt öde skall komma över dig.
Men se, de äro att likna vid strå som brännes upp i eld, de kunna icke rädda sitt liv ur lågornas våld.
Detta är ju ingen koleld att värma sig framför, ingen brasa att sitta vid.
Ja, så går det för dig med dem som du mödade dig för.
Och dina handelsvänner från ungdomstiden draga bort, var och en åt sitt håll och ingen finnes, som frälsar dig.
Hören detta, I av Jakobs hus, I som ären uppkallade med Israels namn och flutna ur Juda källa, I som svärjen vid HERRENS namn och prisen Israels Gud -- dock icke i sanning och rättfärdighet,
allt medan I kallen eder efter den heliga staden och stödjen eder på Israels Gud, på honom vilkens namn är HERREN Sebaot.
Vad förut skedde, det hade jag för länge sedan förkunnat; av min mun var det förutsagt, och jag hade låtit eder höra därom.
Plötsligt satte jag det i verket, och det inträffade.
Eftersom jag visste, att du var så styvsint, ja, att din nacksena var av järn och din panna av koppar,
därför förkunnade jag det för länge sedan och lät dig höra därom, innan det skedde, på det att du icke skulle kunna säga: »Min gudastod har gjort det, min gudabild, den skurna eller den gjutna har skickat det så.»
Du hade hört det, nu kan du se alltsammans; viljen I då icke erkänna det?
Nu låter jag dig åter höra om nya ting, om fördolda ting som du ej har vetat av.
Först nu hava de blivit skapade, icke tidigare, och förrän i dag fick du icke höra om dem, på det att du ej skulle kunna säga: »Det visste jag ju förut.»
Du fick icke förr höra något därom eller veta något därav, ej heller kom det tidigare för dina öron, eftersom jag visste, huru trolös du var och att du hette »överträdare» allt ifrån moderlivet.
Men för mitt namns skull är jag långmodig, och för min äras skull håller jag tillbaka min vrede, så att du icke bliver utrotad.
Se, jag har smält dig, men silver har jag icke fått; jag har prövat dig i lidandets ugn.
För min egen skull, ja, för min egen skull gör jag så, ty huru skulle jag kunna låta mitt namn bliva ohelgat?
Jag giver icke min ära åt någon annan.
Hör på mig, du Jakob, du Israel, som jag har kallat.
Jag är det; jag är den förste, jag är ock den siste.
Min hand har lagt jordens grund, och min högra hand har utspänt himmelen; jag kallar på dem, då stå de där båda.
Församlen eder, I alla, och hören: Vem bland dessa andra har förutsagt detta, att den man, som HERREN älskar, skall utföra hans vilja mot Babel och vara hans arm mot kaldéerna?
Jag, jag har talat detta, jag har ock kallat honom, jag har fört honom fram, så att hans väg har blivit lyckosam.
Träden hit till mig och hören detta; Mina förutsägelser har jag icke talat i det fördolda; när tiden kom, att något skulle ske, då var jag där.
Och nu har Herren, HERREN sänt mig och sänt sin Ande.
Så säger HERREN, din förlossare, Israels Helige: Jag är HERREN, din Gud, den som lär dig, vad nyttigt är, den som leder dig på den väg du skall vandra.
O att du ville akta på mina bud!
Då skulle frid tillflyta dig såsom en ström och din rätt såsom havets böljor;
dina barn skulle då vara såsom sanden och din livsfrukt såsom sandkornen, dess namn skulle aldrig bliva utrotat eller utplånat ur min åsyn.
Dragen ut från Babel, flyn ifrån kaldéernas land; förkunnen det med fröjderop och låten det bliva känt, utbreden ryktet därom till jordens ända; sägen: »HERREN har förlossat sin tjänare Jakob.»
De ledo ingen törst, när han förde dem genom ödemarker, ty han lät vatten strömma fram ur klippan åt dem, han klöv sönder klippan, och vattnet flödade.
Men de ogudaktiga få ingen frid, säger HERREN.
Hören på mig, I havsländer, och akten härpå, I folk, som bon i fjärran.
HERREN kallade mig, när jag ännu var i moderlivet, han nämnde mitt namn, medan jag låg i min moders sköte.
Och han gjorde min mun lik ett skarpt svärd och gömde mig under sin hands skugga; han gjorde mig till en vass pil och dolde mig i sitt koger.
Och han sade till mig: »Du är min tjänare, Israel, genom vilken jag vill förhärliga mig.»
Men jag tänkte: »Förgäves har jag mödat mig, fruktlöst och fåfängt har jag förtärt min kraft; dock, min rätt är hos HERREN och min lön hos min Gud.»
Och nu säger HERREN, han som danade mig till sin tjänare, när jag ännu var i moderlivet, på det att jag måtte föra Jakob tillbaka till honom, så att Israel icke rycktes bort -- ty jag är ärad i HERRENS ögon, och min Gud har blivit min starkhet --
han säger: Det är för litet för dig, då du är min tjänare, att allenast upprätta Jakobs stammar och föra tillbaka de bevarade av Israel; jag vill sätta dig till ett ljus för hednafolken, för att min frälsning må nå till jordens ända.
Så säger HERREN, Israels förlossare, hans Helige, till den djupt föraktade som är en styggelse för människor, en träl under tyranner: Konungar skola se det och stå upp, furstar skola se det och buga sig för HERRENS skull, som har bevisat sig trofast, för Israels Heliges skull, som har utvalt dig.
Så säger HERREN: Jag bönhör dig i behaglig tid, och jag hjälper dig på frälsningens dag; jag skall bevara dig och fullborda i dig förbundet med folket, så att du skall upprätta landet och utskifta de förödda arvslotterna
och säga till de fångna: »Dragen ut», till dem som sitta i mörkret: »Kommen fram.»
De skola finna bete utmed vägarna, ja, betesplatser på alla kala höjder;
de skola varken hungra eller törsta, ökenhettan och solen skola icke skada dem, ty deras förbarmare skall leda dem och skall föra dem till vattenkällor.
Och jag skall göra alla mina berg till öppna vägar, och mina farvägar skola byggas höga.
Se, där komma de fjärran ifrån, ja, somliga från norr och andra från väster, somliga ock från sinéernas land.
Jublen, I himlar, och fröjda dig, du jord, och bristen ut i jubel, I berg; ty HERREN tröstar sitt folk och förbarmar sig över sina betryckta.
Men Sion säger: »HERREN har övergivit mig, Herren har förgätit mig.»
Kan då en moder förgäta sitt barn, så att hon icke har förbarmande med sin livsfrukt?
Och om hon än kunde förgäta sitt barn, så skulle dock jag icke förgäta dig.
Se, på mina händer har jag upptecknat dig; dina murar stå alltid inför mina ögon.
Redan hasta dina söner fram, under det dina förstörare och härjare draga bort ifrån dig.
Lyft upp dina ögon och se dig omkring: alla komma församlade till dig.
Så sant jag lever, säger HERREN, du skall få ikläda dig dem alla såsom en skrud och lik en brud omgjorda dig med dem.
Ty om du förut låg i ruiner och var ödelagd, ja, om ock ditt land var förhärjat, så skall du nu i stället bliva för trång för dina inbyggare, och dina fördärvare skola vara långt borta.
Den tid stundar, då du skall få höra sägas av barnen som föddes under din barnlöshet: »Platsen är mig för trång, giv rum, så att jag kan bo här.»
Då skall du säga i ditt hjärta: »Vem har fött dessa åt mig?
Jag var ju barnlös och ofruktsam, landsflyktig och fördriven; vem har då fostrat dessa?
Se, jag var lämnad ensam kvar; varifrån komma då dessa?»
Så säger Herren, HERREN: Se, jag skall upplyfta min hand till tecken åt folken och resa upp mitt baner till tecken åt folkslagen; då skola de bära dina söner hit i sin famn och föra dina döttrar fram på sina axlar.
Och konungar skola vara dina barns vårdare och furstinnor deras ammor, de skola falla ned inför dig med ansiktet mot jorden och slicka dina fötters stoft.
Och du skall förnimma, att jag är HERREN och att de som förbida mig icke komma på skam.
Kan man taga ifrån hjälten hans byte eller rycka fångarna ifrån den som har segerns rätt?
Och om än så vore, säger HERREN, om man än kunde taga ifrån hjälten hans fångar och rycka bytet ur den väldiges hand, så skulle jag dock själv stå emot dina motståndare, och själv skulle jag frälsa dina barn.
Ja, jag skall tvinga dina förtryckare att äta sitt eget kött, och av sitt eget blod skola de bliva druckna såsom av druvsaft.
Och allt kött skall då förnimma, att jag, HERREN, är din frälsare och att den Starke i Jakob är din förlossare.
Så säger HERREN: Var är eder moders skiljebrev, det, varmed jag skulle hava förskjutit henne?
Eller finnes bland mina borgenärer någon som jag har sålt eder åt?
Nej, genom edra missgärningar bleven I sålda, och för edra överträdelsers skull blev eder moder förskjuten.
Varför var ingen tillstädes, när jag kom?
Varför svarade ingen, när jag ropade?
Har då min arm blivit för kort, så att den ej kan förlossa, eller finnes hos mig ingen kraft till att hjälpa?
Med min näpst uttorkar jag ju havet, och strömmarna gör jag till torrt land, så att fiskarna ruttna och dö av törst, eftersom vattnet är borta;
själva himmelen kläder jag i mörker och giver den sorgdräkt att bära.
Herren, HERREN har givit mig en tunga med lärdom, så att jag förstår att genom mina ord hugsvala den trötte; han väcker var morgon mitt öra, han väcker det till att höra på lärjungesätt.
Ja, Herren, HERREN har öppnat mitt öra, och jag har ej varit gensträvig, jag har ej vikit tillbaka.
Jag höll fram min rygg åt dem som slogo mig och mina kinder åt dem som ryckte mig i skägget; jag skylde icke mitt ansikte mot smädelse och spott.
Men Herren, HERREN hjälper mig, därför kände jag ej smädelsen, därför gjorde jag min panna hård såsom sten; jag visste ju, att jag ej skulle komma på skam.
Den som dömer mig fri är nära, vem vill då gå till rätta med mig?
Må han träda fram jämte mig.
Vem vill vara min anklagare?
Må han komma hit till mig.
Se, Herren, HERREN hjälper mig; vem vill då döma mig skyldig?
Se, de skola allasammans falla sönder såsom en klädnad; mal skall förtära dem.
Vem bland eder, som fruktar HERREN och hör hans tjänares röst?
Om han än vandrar i mörkret och icke ser någon ljusning, så förtröste han dock på HERRENS namn och stödje sig vid sin Gud.
Men se, I alla som tänden upp en brand och väpnen eder med glödande pilar, I hemfallen själva åt lågorna från eder brand och åt pilarna som I haven antänt.
Av min hand skall detta vederfaras eder; i kval skolen I komma att ligga.
Hören på mig, I som faren efter rättfärdighet, I som söken HERREN.
Skåden på klippan, ur vilken I ären uthuggna, och på gruvan, ur vilken I haven framhämtats:
ja, skåden på Abraham, eder fader, och på Sara som födde eder.
Ty när han ännu var ensam, kallade jag honom och välsignade honom och förökade honom.
Ja, HERREN skall varkunna sig över Sion, han skall varkunna sig över alla dess ruiner; han gör dess öken lik ett Eden och dess hedmark lik en HERRENS lustgård.
Fröjd och glädje skall höras därinne, tacksägelse och lovsångs ljud.
Akta på mig, du mitt folk; lyssna till mig, du min menighet.
Ty från mig skall lag utgå, och min rätt skall jag sätta till ett ljus för folken.
Min rättfärdighet är nära, min frälsning går fram, och mina armar skola skaffa rätt bland folken; havsländerna bida efter mig och hoppas på min arm.
Lyften upp edra ögon till himmelen, skåden ock på jorden härnere: se, himmelen skall upplösa sig såsom rök och jorden nötas ut såsom en klädnad, och dess inbyggare skola dö såsom mygg; men min frälsning förbliver evinnerligen, och min rättfärdighet varder icke om intet.
Hören på mig, I som kännen rättfärdigheten, du folk, som bär min lag i ditt hjärta; Frukten icke för människors smädelser och varen ej förfärade för deras hån.
Ty mal skall förtära dem såsom en klädnad, och mott skall förtära dem såsom ull; men min rättfärdighet förbliver evinnerligen och min frälsning ifrån släkte till släkte.
Vakna upp, vakna upp, kläd dig i makt, du HERRENS arm; vakna upp såsom i forna dagar, i förgångna tider.
Var det icke du, som slog Rahab och genomborrade draken?
Var det icke du, som uttorkade havet, det stora djupets vatten, och som gjorde havsbottnen till en väg, där ett frälsat folk kunde gå fram?
Ja, HERRENS förlossade skola vända tillbaka och komma till Sion med jubel; evig glädje skall kröna deras huvuden, fröjd och glädje skola de undfå, sorg och suckan skola fly bort.
Jag, jag är den som tröstar eder.
Vem är då du, att du fruktar för dödliga människor, för människobarn som bliva såsom torrt gräs?
Och därvid förgäter du HERREN, som har skapat dig, honom som har utspänt himmelen och lagt jordens grund.
Ja, beständigt, dagen igenom, förskräckes du för förtryckarens vrede, såsom stode han just redo till att fördärva.
Men vad bliver väl av förtryckarens vrede?
Snart skall den fjättrade lösas ur sitt tvång; han skall icke dö och hemfalla åt graven, ej heller skall han lida brist på bröd.
ty jag är HERREN, din Gud, han som rör upp havet, så att dess böljor brusa, han vilkens namn är HERREN Sebaot;
och jag har lagt mina ord i din mun och övertäckt dig med min hands skugga för att plantera en himmel och grunda en jord och för att säga till Sion: Du är mitt folk.
Vakna upp, vakna upp, stå upp, Jerusalem, du som av HERRENS hand har fått att dricka hans vredes bägare, ja, du som har tömt berusningens kalk till sista droppen.
Bland alla de söner hon hade fött fanns ingen som ledde henne, bland alla de söner hon hade fostrat ingen som fattade henne vid handen.
Dubbel är den olycka som har drabbat dig, och vem visar dig medlidande?
Här är förödelse och förstöring, hunger och svärd.
Huru skall jag trösta dig?
Dina söner försmäktade, de lågo vid alla gathörn, lika antiloper i jägarens garn, drabbade i fullt mått av HERRENS vrede, av din Guds näpst.
Därför må du höra detta, du arma, som är drucken, fastän icke av vin:
Så säger HERREN, som är din Herre, och din Gud, som utför sitt folks sak: Se, jag tager bort ur din hand berusningens bägare; av min vredes kalk skall du ej vidare dricka.
Och jag sätter den i dina plågares hand, deras som sade till dig: »Fall ned, så att vi få gå fram över dig»; och så nödgades du göra din rygg likasom till en mark och till en gata för dem som gingo där fram.
Vakna upp, vakna upp, ikläd dig din makt, o Sion; ikläd dig din högtidsskrud, Jerusalem, du heliga stad; ty ingen oomskuren eller oren skall vidare komma in i dig.
Skaka stoftet av dig, stå upp och intag din plats, Jerusalem; lös banden från din hals, du fångna dotter Sion.
Ty så säger HERREN: I haven blivit sålda för intet; så skolen I ock utan penningar bliva lösköpta.
Ja, så säger Herren, HERREN: Mitt folk drog i forna dagar ned till Egypten och bodde där såsom främlingar; sedan förtryckte Assur dem utan all rätt.
Och vad skall jag nu göra här, säger HERREN, nu då man har fört bort mitt folk utan sak, nu då dess tyranner så skräna, säger HERREN, och mitt namn beständigt, dagen igenom, varder smädat?
Jo, just därför skall mitt folk få lära känna mitt namn, just därför skall det förnimma på den dagen, att jag är den som talar; ja, se här är jag.
Huru ljuvliga äro icke glädjebudbärarens fotsteg, när han kommer över bergen för att förkunna frid och frambära gott budskap och förkunna frälsning, i det han säger till Sion: »Din Gud är nu konung!»
Hör, huru dina väktare upphäva sin röst och jubla allasammans, ty de se för sina ögon, huru HERREN vänder tillbaka till Sion.
Ja, bristen ut i jubel tillsammans, I Jerusalems ruiner; ty HERREN tröstar sitt folk, han förlossar Israel.
HERREN blottar sin heliga arm inför alla hedningars ögon, och alla jordens ändar få se vår Guds frälsning.
Bort, bort, dragen ut därifrån, kommen icke vid det orent är; dragen ut ifrån henne, renen eder, I som bären HERRENS kärl.
Se, I behöven icke draga ut med hast, icke vandra bort såsom flyktingar, ty HERREN går framför eder, och Israels Gud slutar edert tåg.
Se, min tjänare skall hava framgång; han skall bliva upphöjd och stor och högt uppsatt.
Såsom många häpnade över honom, därför att hans utseende var vanställt mer än andra människors och hans gestalt oansenligare än andra människobarns,
så skall han ock väcka förundran hos många folk; ja, konungar skola förstummas i förundran över honom.
Ty vad aldrig har varit förtäljt för dem, det få de se, och vad de aldrig hava hört, det få de förnimma.
Men vem trodde, vad som predikades för oss, och för vem var HERRENS arm uppenbar?
Han sköt upp såsom en ringa telning inför honom, såsom ett rotskott ur förtorkad jord.
Han hade ingen gestalt eller fägring; när vi sågo på honom, kunde hans utseende ej behaga oss.
Föraktat var han och övergiven av människor, en smärtornas man och förtrogen med krankhet; han var såsom en, för vilken man skyler sitt ansikte, så föraktat, att vi höllo honom för intet.
Men det var våra krankheter han bar, våra smärtor, dem lade han på sig, medan vi höllo honom för att vara hemsökt, tuktad av Gud och pinad.
Ja, han var sargad för våra överträdelsers skull och slagen för våra missgärningars skull; näpsten var lagd på honom, för att vi skulle få frid, och genom hans sår bliva vi helade.
Vi gingo alla vilse såsom får, var och en av oss ville vandra sin egen väg, men HERREN lät allas vår missgärning drabba honom.
Han blev plågad, fastän han ödmjukade sig och icke öppnade sin mun, lik ett lamm, som föres bort att slaktas, och lik ett får, som är tyst inför dem som klippa det ja, han öppnade icke sin mun.
Undan våld och dom blev han borttagen, men vem i hans släkte betänker detta?
Ja, han rycktes bort ifrån de levandes land, och för mitt folks överträdelses skull kom plåga över honom.
Och bland de ogudaktiga fick hans in grav bland de rika kom han först, när han var död fastän han ingen orätt hade gjort och fastän svek icke fanns i hans mun.
Det behagade HERREN att slå honom med krankhet: om hans liv så bleve ett skuldoffer, då skulle han få se avkomlingar och länge leva, och HERRENS vilja skulle genom honom hava framgång.
Ja, av den vedermöda hans själ har utstått skall han se frukt och så bliva mättad; genom sin kunskap skall han göra många rättfärdiga, han, den rättfärdige, min tjänare, i det han bär deras missgärningar.
Därför skall jag tillskifta honom hans lott bland de många, och med talrika skaror skall han få utskifta byte, eftersom han utgav sitt liv i döden och blev räknad bland överträdare, han som bar mångas synder och bad för överträdarna.
Jubla, du ofruktsamma, du som icke har fött barn; brist ut i jubel och ropa av fröjd, du som icke har blivit moder.
Ty den ensamma skall hava många barn, flera än den som har man, säger HERREN.
Vidga ut platsen för ditt tjäll, låt spänna ut tältet, under vilket du bor, och spar icke; förläng dina tältstreck och gör dina tältpluggar fastare.
Ty du skall utbreda dig både åt höger och vänster, och dina avkomlingar skola taga hedningarnas länder i besittning och åter befolka ödelagda städer.
Frukta icke, ty du skall ej komma på skam; blygs icke, ty du skall ej varda utskämd.
Nej, du skall få förgäta din ungdoms skam, och ditt änkestånds smälek skall du icke mer komma ihåg.
Ty den som har skapat dig är din man, han vilkens namn är HERREN Sebaot; och Israels Helige är din förlossare, han som kallas hela jordens Gud.
Ty såsom en övergiven kvinna i hjärtesorg kallades du av HERREN.
Sin ungdomsbrud, vill någon förskjuta henne? säger din Gud.
Ett litet ögonblick övergav jag dig, men i stor barmhärtighet vill jag åter församla dig.
I min förtörnelses översvall dolde jag ett ögonblick mitt ansikte för dig, men med evig nåd vill jag nu förbarma mig över dig, säger HERREN, din förlossare.
Ty såsom jag gjorde vid Noas flod, så gör jag ock nu: såsom jag då svor, att Noas flod icke mer skulle komma över jorden, så svär jag ock nu, att jag icke mer skall förtörnas på dig eller näpsa dig.
Ja, om än bergen vika bort och höjderna vackla, så skall min nåd icke vika ifrån dig och mitt fridsförbund icke vackla, säger HERREN; din förbarmare.
Du arma, som har blivit så hemsökt av stormar utan att få någon tröst, se, med spetsglans vill jag nu mura dina stenar och giva dig grundvalar av safirer,
jag vill göra dina tinnar av rubiner och dina portar av kristall och hela din ringmur av ädla stenar.
Och dina barn skola alla bliva HERRENS lärjungar, och stor frid skola dina barn då hava.
Genom rättfärdighet skall du bliva befäst.
All tanke på förtryck vare fjärran ifrån dig, ty du skall intet hava att frukta, och all tanke på fördärv, ty sådant skall icke nalkas dig.
Om man då rotar sig samman till anfall, så kommer det ingalunda från mig; och vilka de än äro, som rota sig samman mot dig, så skola de falla för dig.
Se, jag är den som skapar smeden, vilken blåser upp kolelden och så frambringar ett vapen, sådant han vill göra det; men jag är ock den som skapar fördärvaren, vilken förstör det.
Och nu skall intet vapen, som smides mot dig, hava någon lycka; var tunga, som upphäver sig för att gå till rätta med dig, skall du få domfälld.
Detta är HERRENS tjänares arvedel, den rätt de skola undfå av mig, säger HERREN.
Upp, alla I som ären törstiga, kommen hit och fån vatten; och I som inga penningar haven, kommen hit och hämten säd och äten.
Ja, kommen hit och hämten säd utan penningar och för intet både vin och mjölk.
Varför given I ut penningar för det som ej är bröd och edert förvärv för det som icke kan mätta?
Hören på mig, så skolen I få äta det gott är och förnöja eder med feta rätter.
Böjen edra öron hit och kommen till mig; hören, så får eder själ leva.
Jag vill sluta med eder ett evigt förbund: att I skolen undfå all den trofasta nåd jag har lovat David.
Se, honom har jag satt till ett vittne för folken, till en furste och hövding för folken.
Ja, du skall kalla på folkslag som du icke känner, och folkslag, som icke känna dig, skola hasta till dig för HERRENS, din Guds, skull, för Israels Heliges skull, när han förhärligar dig.
Söken HERREN, medan han låter sig finnas; åkallen honom, medan han är nära.
Den ogudaktige övergive sin väg och den orättfärdige sina tankar och vände om till HERREN, så skall han förbarma sig över honom, och till vår Gud, ty han skall beskära mycken förlåtelse.
Se, mina tankar äro icke edra tankar, och edra vägar äro icke mina vägar, säger HERREN.
Nej, så mycket som himmelen är högre än jorden, så mycket äro ock mina vägar högre än edra vägar och mina tankar högre än edra tankar.
Ty likasom regnet och snön faller ifrån himmelen och icke vänder tillbaka dit igen, förrän det har vattnat jorden och gjort den fruktsam och bärande, så att den giver säd till att så och bröd till att äta,
så skall det ock vara med ordet som utgår ur min mun; det skall icke vända tillbaka till mig fåfängt utan att hava verkat, vad jag vill, och utfört det, vartill jag hade sänt ut det.
Ty med glädje skolen I draga ut, och i frid skolen I föras åstad.
Bergen och höjderna skola brista ut i jubel, där I gån fram, och alla träd på marken skola klappa i händerna.
Där törnsnår nu finnas skola cypresser växa upp, och där nässlor stå skall myrten uppväxa.
Och detta skall bliva HERREN till ära och ett evigt tecken, som ej skall plånas ut.
Så säger HERREN: Akten på vad rätt är och öven rättfärdighet, ty min frälsning kommer snart, och snart bliver min rättfärdighet uppenbarad.
Säll är den människa, som gör detta, den människoson, som står fast därvid, den som håller sabbaten, så att han icke ohelgar den, och den som avhåller sin hand från att göra något ont.
Främlingen, som har slutit sig till HERREN, må icke säga så: »Säkert skall HERREN avskilja mig från sitt folk.»
Ej heller må den snöpte säga: »Se, jag är ett förtorkat träd.»
Ty så säger HERREN: De snöpta, som hålla mina sabbater och utvälja det mig behagar och stå fast vid mitt förbund,
åt dem skall jag i mitt hus och inom mina murar giva en åminnelse och ett namn, en välsignelse, som är förmer än söner och döttrar; jag skall giva dem ett evigt namn, som icke skall varda utrotat.
Och främlingarna, som hava slutit sig till HERREN för att tjäna honom och för att älska HERRENS namn och så vara hans tjänare, alla som hålla sabbaten, så att de icke ohelga den, och som stå fast vid mitt förbund,
dem skall jag låta komma till mitt heliga berg och giva dem glädje i mitt bönehus, och deras brännoffer och slaktoffer skola vara mig välbehagliga på mitt altare; ty mitt hus skall kallas ett bönehus för alla folk.
Så säger Herren, HERREN, han som församlar de fördrivna av Israel: Jag skall församla ännu flera till honom, utöver dem som redan äro församlade till honom.
I alla djur på marken, kommen och äten, ja, I alla skogens djur.
Väktarna här äro allasammans blinda, de hava intet förstånd; de äro allasammans stumma hundar, som icke kunna skälla; de ligga och drömma och vilja gärna slumra.
Men de hundarna äro ock glupska och kunna ej bliva mätta.
Ja, sådana människor äro herdar, dessa som intet kunna förstå!
De vilja allasammans vandra sin egen väg; var och en söker sin egen vinning, alla, så många de äro.
»Kommen, jag skall hämta vin, och så skola vi dricka oss druckna av starka drycker.
Och morgondagen skall bliva denna dag lik, en övermåttan härlig dag!»
Den rättfärdige förgås, och ingen finnes, som tänker därpå; fromma människor ryckas bort, utan att någon lägger märke därtill.
Ja, genom ondskans makt ryckes den rättfärdige bort
och går då in i friden; de som hava vandrat sin väg rätt fram få ro i sina vilorum.
Men träden fram hit, I söner av teckentyderskor, I barn av äktenskapsbrytare och skökor.
Över vem gören I eder lustiga?
Mot vem spärren I upp munnen och räcken I ut tungan?
Sannerligen, I ären överträdelsens barn, en lögnens avföda,
I som upptändens av brånad vid terebinterna, ja, under alla gröna träd, I som slakten edra barn i dalarna, i bergsklyftornas djup.
Stenarna i din dal har du till din del, de, just de äro din lott; också åt dem utgjuter du drickoffer och frambär du spisoffer.
Skulle jag giva mig till freds vid sådant?
På höga och stora berg redde du dig läger; också upp på sådana begav du dig för att offra slaktoffer.
Och bakom dörren och dörrposten satte du ditt märke.
Du övergav mig; du klädde av dig och besteg ditt läger och beredde plats där.
Du gjorde upp med dem, gärna delade du läger med dem vid första vink du såg.
Du begav dig till Melek med olja och tog med dig dina många salvor; du sände dina budbärare till fjärran land, ja, ända ned till dödsriket.
Om du än blev trött av din långa färd, sade du dock icke: »Förgäves!»
Så länge du kunde röra din hand, mattades du icke.
För vem räddes och fruktade du då, eftersom du var så trolös och eftersom du icke tänkte på mig och ej ville akta på?
Är det icke så: eftersom jag har tegat, och det sedan länge, därför fruktar du mig icke?
Men jag skall visa, huru det är med din rättfärdighet och med dina verk, de skola icke hjälpa dig.
När du ropar, då må ditt avgudafölje rädda dig.
Nej, en vind skall taga dem med sig allasammans och en fläkt föra dem bort.
Men den som tager sin tillflykt till mig skall få landet till arvedel och få besitta mitt heliga berg.
Ja, det skall heta: »Banen väg, banen och bereden väg; skaffen bort stötestenarna från mitt folks väg.»
Ty så säger den höge och upphöjde, han som tronar till evig tid och heter »den Helige»: Jag bor i helighet uppe i höjden, men ock hos den som är förkrossad och har en ödmjuk ande; ty jag vill giva liv åt de ödmjukas ande och liv åt de förkrossades hjärtan.
Ja, jag vill icke evinnerligen gå till rätta och icke ständigt förtörnas; eljest skulle deras ande försmäkta inför mig, de själar, som jag själv har skapat.
För hans girighetssynd förtörnades jag; jag slog honom, och i min förtörnelse höll jag mig dold.
Men i sin avfällighet fortfor han att vandra på sitt hjärtas väg.
Hans vägar har jag sett, men nu vill jag hela honom och leda honom och giva honom och hans sörjande tröst.
Jag skall skapa frukt ifrån hans läppar.
Frid över dem som äro fjärran och frid över dem som äro nära! säger HERREN; jag skall hela honom.
Men de ogudaktiga äro såsom ett upprört hav, ett som icke kan vara stilla, ett hav, vars vågor röra upp dy och orenlighet.
De ogudaktiga hava ingen frid, säger min Gud.
Ropa med full hals utan återhåll, häv upp din röst såsom en basun och förkunna för mitt folk deras överträdelse, för Jakobs hus deras synder.
Väl söka de mig dag ut och dag in och vilja hava kunskap om mina vägar.
Såsom vore de ett folk, som övade rättfärdighet och icke övergåve sin Guds rätt, så fråga de mig om rättfärdighetens rätter och vilja, att Gud skall komma till dem:
»Vartill gagnar det, att vi fasta, när du icke ser det, vartill, att vi späka oss, när du icke märker det?»
Men se, på edra fastedagar sköten I edra sysslor, och alla edra arbetare driven I blott på.
Och se, I hållen eder fasta med kiv och split, med hugg och slag av gudlösa nävar.
I hållen icke mer fasta på sådant sätt, att I kunnen göra eder röst hörd i höjden.
Skulle detta vara en fasta, sådan som jag vill hava?
Skulle detta vara en rätt späkningsdag?
Att man hänger med huvudet såsom ett sävstrå och sätter sig i säck och aska, vill du kalla sådant att hålla fasta, att fira en dag till HERRENS behag?
Nej, detta är den fasta, som jag vill hava: att I lossen orättfärdiga bojor och lösen okets band, att I given de förtryckta fria och krossen sönder alla ok,
ja, att du bryter ditt bröd åt den hungrige och skaffar de fattiga och husvilla härbärge att du kläder den nakne, var du ser honom, och ej drager dig undan för den som är ditt kött och blod.
Då skall ljus bryta fram för dig såsom en morgonrodnad, och dina sår skola läkas med hast, och din rätt skall då gå framför dig och HERRENS härlighet följa dina spår.
Då skall HERREN svara, när du åkallar honom; när du ropar, skall han säga: »Se, här är jag.»
Om hos dig icke får finnas någon som pålägger ok och pekar finger och talar, vad fördärvligt är,
om du delar med dig av din nödtorft åt den hungrige och mättar den som är i betryck, då skall ljus gå upp för dig i mörkret, och din natt skall bliva lik middagens sken.
Och HERREN skall leda dig beständigt; han skall mätta dig mitt i ödemarken och giva styrka åt benen i din kropp.
Och du skall vara lik en vattenrik trädgård och likna ett källsprång, vars vatten aldrig tryter.
Och dina avkomlingar skola bygga upp de gamla ruinerna, du skall åter upprätta grundvalar ifrån forna släkten; och du skall kallas »han som murar igen revor», »han som återställer stigar, så att man kan bo i landet.»
Om du är varsam med din fot på sabbaten, så att du icke på min heliga dag utför dina sysslor; om du kallar sabbaten din lust och HERRENS helgdag en äredag, ja, om du ärar den, så att du icke går dina egna vägar eller sköter dina sysslor eller talar tomma ord,
då skall du finna din lust i HERREN, och jag skall föra dig fram över landets höjder och giva dig till näring din fader Jakobs arvedel.
Ja, så har HERRENS mun talat.
Se, HERRENS arm är icke för kort, så att han ej kan frälsa, och hans öra är icke tillslutet, så att han ej kan höra.
Nej, det är edra missgärningar, som skilja eder och eder Gud från varandra, och edra synder dölja hans ansikte för eder, så att han icke hör eder.
Ty edra händer äro fläckade av blod och edra fingrar av missgärning, edra läppar tala lögn, och eder tunga frambär orättfärdighet.
Ingen höjer sin röst i rättfärdighetens namn, och ingen visar redlighet i vad till rätten hör.
De förtrösta på idel tomhet, de tala falskhet, de gå havande med olycka och föda fördärv.
De kläcka ut basiliskägg och väva spindelnät.
Om någon äter av deras ägg, så dör han, och trampas ett sådant sönder, så kommer en huggorm ut.
Deras spindelnät duga icke till kläder, och de kunna ej skyla sig med vad de hava tillverkat; deras verk äro fördärvliga verk, och våldsgärningar öva deras händer.
Deras fötter hasta till vad ont är och äro snara, när det gäller att utgjuta oskyldigt blod; deras tankar äro fördärvliga tankar, förödelse och förstöring är på deras vägar.
Fridens väg känna de icke, och rätten följer ej i deras spår; de gå krokiga stigar, och ingen som vandrar så vet, vad frid är.
Därför är rätten fjärran ifrån oss, och rättfärdighet tillfaller oss icke; vi bida efter ljus, men se, mörker råder, efter solsken, men vi få vandra i djupaste natt.
Vi måste famla utefter väggen såsom blinda, famla, såsom hade vi inga ögon; vi stappla mitt på dagen, såsom vore det skymning, mitt i vår fulla kraft äro vi såsom döda.
Vi brumma allasammans såsom björnar och sucka alltjämt såsom duvor; vi bida efter rätten, men den kommer icke, efter frälsningen, men den är fjärran ifrån oss.
Ty många äro våra överträdelser inför dig, och våra synder vittna emot oss; ja, våra överträdelser hava vi för våra ögon, och våra missgärningar känna vi.
Genom överträdelse och förnekelse hava vi felat mot HERREN, vi hava vikit bort ifrån vår Gud; vi hava talat förtryck och avfällighet, lögnläror hava vi förkunnat och hämtat fram ur våra hjärtan.
Rätten tränges tillbaka, och rättfärdigheten står långt borta, ja, sanningen vacklar på torget, och vad rätt är kan ej komma fram.
Så måste sanningen hålla sig undan, och den som vände sig ifrån det onda blev plundrad.
Detta såg HERREN, och det misshagade honom, att det icke fanns någon rätt.
Och han såg, att ingen trädde fram; han förundrade sig över att ingen grep in.
Då hjälpte honom hans egen arm, och hans rättfärdighet understödde honom.
Och han klädde sig i rättfärdighet såsom i ett pansar och satte frälsningens hjälm på sitt huvud; han klädde sig i hämndens dräkt såsom i en livklädnad och höljde sig i nitälskan såsom i en mantel.
Efter deras gärningar skall han nu vedergälla dem; vrede skall han låta komma över sina ovänner och över sina fiender lönen för vad de hava gjort; ja, havsländerna skall han vedergälla, vad de hava gjort.
Så skall HERRENS namn bliva fruktat i väster och hans härlighet, där solen går upp.
När fienden bryter fram lik en ström, skall HERRENS andedräkt förjaga honom.
Men såsom en förlossare kommer HERREN för Sion och för dem i Jakob, som omvända sig från sin överträdelse, säger HERREN.
Och detta är det förbund, som jag å min sida gör med dem, säger HERREN: min Ande, som är över dig, och orden, som jag har lagt i din mun, de skola icke vika ur din mun, ej heller ur dina barns eller barnbarns mun från nu och till evig tid, säger HERREN.
Stå upp, var ljus, ty ditt ljus kommer, och HERRENS härlighet går upp över dig.
Se, mörker övertäcker jorden och töcken folken, men över dig uppgår HERREN, och hans härlighet uppenbaras över dig.
Och folken skola vandra i ditt ljus och konungarna i glansen som går upp över dig.
Lyft upp dina ögon och se dig omkring: alla komma församlade till dig; dina söner komma fjärran ifrån, och dina döttrar bäras fram på armen.
Då, vid den synen skall du stråla av fröjd, och ditt hjärta skall bäva och vidga sig; ty havets rikedomar skola föras till dig, och folkens skatter skola falla dig till.
Skaror av kameler skola övertäcka dig, kamelfålar från Midjan och Efa; från Saba skola de alla komma, guld och rökelse skola de bära och skola förkunna HERRENS lov.
Alla Kedars hjordar skola församlas till dig, Nebajots vädurar skola vara dig till tjänst.
Mig till välbehag skola de offras på mitt altare, och min härlighets hus skall jag så förhärliga.
Vilka äro dessa som komma farande lika moln, lika duvor, som flyga till sitt duvslag?
Se, havsländerna bida efter mig, och främst komma Tarsis' skepp; de vilja föra dina söner hem ifrån fjärran land, och de hava med sig silver och guld åt HERRENS, din Guds, namn, åt Israels Helige, ty han förhärligar dig.
Och främlingar skola bygga upp dina murar, och deras konungar skola betjäna dig.
Ty väl har jag slagit dig i min förtörnelse, men i min nåd förbarmar jag mig nu över dig.
Och dina portar skola hållas öppna beständigt, varken dag eller natt skola de stängas, så att folkens skatter kunna föras in i dig, med deras konungar i hyllningståget.
Ty det folk eller rike, som ej vill tjäna dig, skall förgås; ja, sådana folk skola i grund förgöras.
Libanons härlighet skall komma till dig, både cypress och alm och buxbom, för att pryda platsen, där min helgedom är; ty den plats, där mina fötter stå, vill jag göra ärad.
Och bugande skola dina förtryckares söner komma till dig, och dina föraktare skola allasammans falla ned för dina fötter.
Och man skall kalla dig »HERRENS stad», »Israels Heliges Sion».
I stället för att du var övergiven och hatad, så att ingen ville taga vägen genom dig, skall jag göra dig till en härlighetens boning evinnerligen och till en fröjdeort ifrån släkte till släkte.
Och du skall dia folkens mjölk, ja, konungabröst skall du dia; och du skall förnimma, att jag, HERREN, är din frälsare och att den Starke i Jakob är din förlossare.
Jag skall låta guld komma i stället för koppar och låta silver komma i stället för järn och koppar i stället för trä och järn i stället för sten.
Och jag vill sätta frid till din överhet och rättfärdighet till din behärskare.
Man skall icke mer höra talas om våld i ditt land, om ödeläggelse och förstöring inom dina gränser, utan du skall kalla dina murar för »frälsning» och dina portar för »lovsång».
Solen skall icke mer vara ditt ljus om dagen, och månen skall icke mer lysa dig med sitt sken, utan HERREN skall vara ditt eviga ljus, och din Gud skall vara din härlighet.
Din sol skall då icke mer gå ned och din måne icke mer taga av; ty HERREN skall vara ditt eviga ljus, och dina sorgedagar skola hava en ände.
Och i ditt folk skola alla vara rättfärdiga, evinnerligen skola de besitta landet; de äro ju en telning, som jag har planterat, ett verk av mina händer, som jag vill förhärliga mig med.
Av den minste skola komma tusen, och av den ringaste skall bliva ett talrikt folk.
Jag är HERREN; när tiden är inne, skall jag med hast fullborda detta.
Herrens, HERRENS Ande är över mig, ty HERREN har smort mig till att förkunna glädjens budskap för de ödmjuka; han har sänt mig till att läka dem som hava ett förkrossat hjärta, till att predika frihet för de fångna och förlossning för de bundna,
till att predika ett nådens år från HERREN och en hämndens dag från vår Gud, en dag, då han skall trösta alla sörjande,
då han skall låta de sörjande i Sion få huvudprydnad i stället för aska, glädjeolja i stället för sorg, högtidskläder i stället för en bedrövad ande; och de skola kallas »rättfärdighetens terebinter», »HERRENS plantering, som han vill förhärliga sig med».
Och de skola bygga upp de gamla ruinerna och upprätta förfädernas ödeplatser; de skola återställa de förödda städerna, de platser, som hava legat öde släkte efter släkte.
Främlingar skola stå redo att föra edra hjordar i bet, och utlänningar skola bruka åt eder åkrar och vingårdar.
Men I skolen heta HERRENS präster, och man skall kalla eder vår Guds tjänare; I skolen få njuta av folkens skatter, och deras härlighet skall övergå till eder.
För eder skam skolen I få dubbelt igen, och de som ledo smälek skola nu jubla över sin del.
Så skola de få dubbelt att besitta i sitt land; evig glädje skola de undfå.
Ty jag, HERREN, älskar, vad rätt är, och hatar orättfärdigt rov; och jag skall giva dem deras lön i trofasthet och sluta ett evigt förbund med dem.
Och deras släkte skall bliva känt bland folken och deras avkomma bland folkslagen; alla som se dem skola märka på dem, att de äro ett släkte, som HERREN har välsignat.
Jag gläder mig storligen i HERREN, och min själ fröjdar sig i min Gud, ty han har iklätt mig frälsningens klädnad och höljt mig i rättfärdighetens mantel, likasom när en brudgum sätter högtidsbindeln på sitt huvud eller likasom när en brud pryder sig med sina smycken.
Ty likasom jorden låter sina växter spira fram och en trädgård sin sådd växa upp, så skall Herren, HERREN låta rättfärdighet uppväxa och lovsång inför alla folk.
För Sions skull vill jag icke tiga, och för Jerusalems skull vill jag ej unna mig ro, förrän dess rätt går upp såsom solens sken och dess frälsning lyser såsom ett brinnande bloss.
Och folken skola se din rätt och alla konungar din härlighet; och du skall få ett nytt namn, som HERRENS mun skall bestämma.
Så skall du vara en härlig krona i HERRENS hand, en konungslig huvudbindel i din Guds hand.
Du skall icke mer kallas »den övergivna», ej heller skall ditt land mer kallas »ödemark», utan du skall få heta »hon som jag har min lust i», och ditt land skall få heta »äkta hustrun»; ty HERREN har sin lust i dig, och ditt land har fått sin äkta man.
Ty såsom när en ung man bliver en jungrus äkta herre, så skola dina barn bliva dina äkta herrar, och såsom en brudgum fröjdar sig över sin brud, så skall din Gud fröjda sig över dig.
På dina murar, Jerusalem, har jag ställt väktare; varken dag eller natt få de någonsin tystna.
I som skolen ropa till HERREN, given eder ingen ro.
Och given honom ingen ro förrän han åter har byggt upp Jerusalem och låtit det bliva ett ämne till lovsång på jorden.
HERREN har svurit vid sin högra hand och sin starka arm: Jag skall icke mer giva din säd till mat åt dina fiender, och främlingar skola icke dricka ditt vin, frukten av din möda.
Nej, de som insamla säden skola ock äta den och skola lova HERREN, och de som inbärga vinet skola dricka det i min helgedoms gårdar.
Dragen ut, dragen ut genom portarna, bereden väg för folket; banen, ja, banen en farväg rensen den från stenar, resen upp ett baner för folken.
Hör, HERREN höjer ett rop, och det når till jordens ända: Sägen till dottern Sion: Se, din frälsning kommer.
Se, han har med sig sin lön, och hans segerbyte går framför honom.
Och man skall kalla dem »det heliga folket», »HERRENS förlossade»; och dig själv skall man kalla »den mångbesökta staden», »staden, som ej varder övergiven».
Vem är han som kommer från Edom, från Bosra i högröda kläder, så präktig i sin dräkt, så stolt i sin stora kraft? »Det är jag, som talar i rättfärdighet, jag, som är en mästare till att frälsa.»
Varför är din dräkt så röd?
Varför likna dina kläder en vintrampares?
»Jo, en vinpress har jag trampat, jag själv allena, och ingen i folken bistod mig.
Jag trampade dem i min vrede, trampade sönder dem i min förtörnelse.
Då stänkte deras blod på mina kläder, och så fick jag hela min dräkt nedfläckad.
Ty en hämndedag hade jag beslutit, och mitt förlossningsår hade kommit.
Och jag skådade omkring mig, men ingen hjälpare fanns; jag stod där i förundran, men ingen fanns, som understödde mig.
Då hjälpte mig min egen arm, och min förtörnelse understödde mig.
Jag trampade ned folken i min vrede och gjorde dem druckna i min förtörnelse, och jag lät deras blod rinna ned på jorden.»
HERRENS nådegärningar vill jag förkunna, ja, HERRENS lov, efter allt vad HERREN har gjort mot oss, den nåderike mot Israels hus, vad han har gjort mot dem efter sin barmhärtighet och sin stora nåd.
Ty han sade: »De äro ju mitt folk, barn, som ej svika.»
Och så blev han deras frälsare.
I all deras nöd var ingen verklig nöd, ty hans ansiktes ängel frälste dem.
Därför att han älskade dem och ville skona dem, förlossade han dem.
Han lyfte dem upp och bar dem alltjämt, i forna tider.
Men de voro gensträviga, och de bedrövade hans heliga Ande; därför förvandlades han till deras fiende, han själv stridde mot dem.
Då tänkte hans folk på forna tider, de tänkte på Mose: Var är nu han som förde dem upp ur havet, jämte herdarna för hans hjord?
Var är han som lade i deras bröst sin helige Ande,
var är han som lät sin härliga arm gå fram vid Moses högra sida, han som klöv vattnet framför dem och så gjorde sig ett evigt namn,
han som lät dem färdas genom djupen, såsom hästar färdas genom öknen, utan att stappla?
Likasom när boskapen går ned i dalen så fördes de av HERRENS Ande till ro.
Ja, så ledde du ditt folk och gjorde dig ett härligt namn.
Skåda ned från himmelen och se härtill från din heliga och härliga boning.
Var äro nu din nitälskan och dina väldiga gärningar, var är ditt hjärtas varkunnsamhet och din barmhärtighet?
De hålla sig tillbaka från mig.
Du är ju dock vår fader; ty Abraham vet icke av oss, och Israel känner oss icke.
Men du, HERRE, är vår fader; »vår förlossare av evighet», det är ditt namn.
Varför, o HERRE, låter du oss då gå vilse från dina vägar och förhärdar våra hjärtan, så att vi ej frukta dig?
Vänd tillbaka för dina tjänares skull, för din arvedels stammars skull.
Allenast helt kort fick ditt heliga folk behålla sin besittning; våra ovänner trampade ned din helgedom.
Det är oss nu så, som om du aldrig hade varit herre över oss, om om vi ej hade blivit uppkallade efter ditt namn.
O att du läte himmelen rämna och fore hitned, så att bergen skälvde inför dig,
likasom när ris antändes av eld och vatten genom eld bliver sjudande, så att du gjorde ditt namn kunnigt bland dina ovänner och folken darrade för dig!
O att du fore hitned med underbara gärningar som vi icke kunde vänta, så att bergen skälvde inför dig!
Aldrig någonsin har man ju hört, aldrig har något öra förnummit, aldrig har något öga sett en annan Gud än dig handla så mot dem som vänta efter honom.
Du kom dem till mötes, som övade rättfärdighet med fröjd, dem som på dina vägar tänkte på dig.
Men se, du blev förtörnad, och vi stodo där såsom syndare.
Så hava vi länge stått; skola vi väl bliva frälsta?
Vi blevo allasammans lika orena människor, och all vår rättfärdighet var såsom en fläckad klädnad.
Vi vissnade allasammans såsom löv, och våra missgärningar förde oss bort såsom vinden.
Ingen fanns, som åkallade ditt namn, ingen, som vaknade upp för att hålla sig till dig; ty du dolde ditt ansikte för oss och lät oss försmäkta genom vår missgärning.
Men HERRE, du är ju vår fader; vi äro leret, och du är den som har danat oss, vi äro allasammans verk av din hand.
Var då ej så högeligen förtörnad, HERRE; och tänk icke evinnerligen på vår missgärning; nej, se därtill att vi allasammans äro ditt folk.
Dina heliga städer hava blivit en öken, Sion har blivit en öken, Jerusalem en ödemark.
Vårt heliga och härliga tempel, där våra fäder lovade dig, det har blivit uppbränt i eld; och allt vad dyrbart vi ägde har lämnats åt förödelsen.
Kan du vid allt detta hålla dig tillbaka, o HERRE?
Kan du tiga stilla och plåga oss så svårt?
Jag har låtit mig bliva uppenbar för dem som icke frågade efter mig, jag har låtit mig finnas av dem som icke sökte mig; till ett folk som icke var uppkallat efter mitt namn har jag sagt: Se, här är jag, här är jag.
Hela dagen har jag uträckt mina händer till ett gensträvigt folk som vandrar på den väg som icke är god, i det att de följa sina egna tankar --
ett folk, som beständigt förtörnar mig utan att hava någon försyn, som frambär offer i lustgårdar och tänder offereld på tegelaltaren,
som har sitt tillhåll bland gravar och tillbringar natten i undangömda nästen, som äter svinens kött och har vederstygglig spis i sina kärl,
som säger: »Bort med dig, kom icke vid mig, ty jag är helig för dig.»
De äro såsom rök i min näsa, en eld, som brinner beständigt.
Se, detta står upptecknat inför mina ögon; jag skall icke tiga, förrän jag har givit vedergällning, ja, vedergällning i deras sköte,
både för deras egna missgärningar och för deras fäders, säger HERREN, vedergällning för att de tände offereld på bergen och för att de smädade mig på höjderna; ja, först skall jag mäta upp lönen åt dem i deras sköte.
Så säger HERREN: Likasom man säger om en druvklase, när däri finnes saft: »Fördärva den icke, ty välsignelse är däri», så skall ock jag göra för mina tjänares skull: jag skall icke fördärva alltsammans.
Jag skall låta en avkomma utgå från Jakob, från Juda en arvinge till mina berg; ty mina utkorade skola besitta landet, och mina tjänare skola bo däri.
Saron skall bliva en betesmark för får och Akors dal en lägerplats för fäkreatur, och de skola givas åt mitt folk, när det söker mig.
Men I som övergiven HERREN och förgäten mitt heliga berg, I som duken bord åt Gad och iskänken vindryck åt Meni,
eder har jag bestämt åt svärdet, och I skolen alla få böja eder ned till att slaktas, därför att I icke svaraden, när jag kallade, och icke hörden, när jag talade, utan gjorden, vad ont var i mina ögon, och utvalden det som var mig misshagligt.
Därför säger Herren, HERREN så: Se, mina tjänare skola äta, men I skolen hungra; se, mina tjänare skola dricka, men I skolen törsta; se, mina tjänare skola glädjas, men I skolen få blygas.
Ja, mina tjänare skola jubla i sitt hjärtas fröjd, men I skolen ropa i edert hjärtas plåga och jämra eder i förtvivlan.
Och I skolen lämna edert namn till ett förbannelsens ord, så att mina utkorade skola säga: »Sådan död give dig Herren, HERREN.»
Men åt sina tjänare skall han giva ett annat namn:
den som då välsignar sig i landet skall välsigna sig i »den sannfärdige Guden», och den som svär i landet, han skall svärja vid »den sannfärdige Guden».
Ty de förra bedrövelserna äro då förgätna och dolda för mina ögon.
Ty se, jag vill skapa nya himlar och en ny jord; och man skall ej mer komma ihåg det förgångna eller tänka därpå.
Nej, I skolen fröjdas och jubla till evig tid över det som jag skapar; ty se, jag vill skapa Jerusalem till jubel och dess folk till fröjd.
Och jag skall jubla över Jerusalem och fröjda mig över mitt folk, och där skall icke mer höras gråt eller klagorop.
Där skola icke mer finnas barn som leva allenast några dagar, ej heller gamla män, som icke fylla sina dagars mått; nej, den som dör ung skall dö först vid hundra års ålder, och först vid hundra års ålder skall syndaren drabbas av förbannelsen.
När de bygga hus, skola de ock få bo i dem; när de plantera vingårdar, skola de ock få äta deras frukt.
När de bygga hus, skall det ej bliva andra, som få bo i dem; när de plantera något, skall det ej bliva andra, som få äta därav.
Ty samma ålder, som ett träd uppnår, skall man uppnå i mitt folk, och mina utkorade skola själva njuta av sina händers verk.
De skola icke möda sig förgäves, och barnen, som de föda, drabbas ej av plötslig död; ty de äro ett släkte av HERRENS välsignade, och deras avkomlingar få leva kvar bland dem.
Och det skall ske, att förrän de ropa, skall jag svara, och medan de ännu tala, skall jag höra.
Då skola vargar gå i bet tillsammans med lamm, och lejon skola äta halm likasom oxar, och stoft skall vara ormens föda.
Ingenstädes på mitt heliga berg skall man då göra, vad ont och fördärvligt är, säger HERREN.
Så säger HERREN: Himmelen är min tron, och jorden är min fotapall; vad för ett hus skullen I då kunna bygga åt mig, och vad för en plats skulle tjäna mig till vilostad?
Min hand har ju gjort allt detta, och så har allt detta blivit till, säger HERREN.
Men till den skådar jag ned, som är betryckt och har en förkrossad ande, och till den som fruktar för mitt ord.
Den däremot, som slaktar sin offertjur, men ock är en mandråpare, den som offrar sitt lamm, men tillika krossar nacken på en hund, den som frambär ett spisoffer, men därvid frambär svinblod, den som offrar rökelse, men därunder hyllar en fåfänglig avgud -- likasom det lyster dessa att gå sina egna vägar och likasom deras själ har behag till deras styggelser,
så lyster det ock mig att fara illa fram med dem och att låta förskräckelse komma över dem, eftersom ingen svarade, när jag kallade, och eftersom de icke hörde, när jag talade, utan gjorde, vad ont var i mina ögon, och hade sin lust i att göra, vad mig misshagligt var.
Hören HERRENS ord, I som frukten för hans ord.
Edra bröder, som hata eder och stöta eder bort för mitt namns skull, de säga: »Må HERREN förhärliga sig, så att vi få se eder glädje.»
Men de skola komma på skam.
Hör, huru det larmar i staden, hör dånet i templet!
Hör dånet, när HERREN vedergäller sina fiender, vad de hava gjort!
Innan Sion har känt någon födslovånda, föder hon barnet; innan kval har kommit över henne, bliver hon förlöst med ett gossebarn.
Vem har hört något sådant, vem har sett något dylikt?
Kan då ett land komma till liv på en enda dag, eller kan ett folk födas i ett ögonblick, eftersom Sion födde fram sina barn, just då våndan begynte?
Ja, ty skulle jag väl låta fostret bliva fullgånget, men icke giva kraft att föda fram det? säger HERREN.
Eller skulle jag giva kraft att föda, men sedan hålla fostret tillbaka? säger din Gud.
Glädjens med Jerusalem och fröjden eder över henne, alla I som haven henne kär; jublen högt med henne, alla I som haven sörjt över henne.
Så skolen I få dia eder mätta vid hennes hugsvalelses bröst; så skolen I få suga med lust av hennes rika barm.
Ty så säger HERREN: Se, jag vill låta frid komma över henne såsom en ström och folkens rikedomar såsom en översvämmande flod, och I skolen så få dia, I skolen bliva burna på armen och skolen få sitta i knäet och bliva smekta.
Såsom en moder tröstar sin son, så skall jag trösta eder; ja, i Jerusalem skolen I få tröst.
Och edra hjärtan skola glädja sig, när I fån se detta, och benen i edra kroppar skola hava livskraft såsom spirande gräs; och man skall förnimma, att HERRENS hand är med hans tjänare och att ogunst kommer över hans fiender.
Ty se, HERREN skall komma i eld, och hans vagnar skola vara såsom en stormvind; och han skall låta sin vrede drabba med hetta och sin näpst med eldslågor.
Ty HERREN skall hålla dom med eld, och med sitt svärd skall han slå allt kött, och många skola de vara, som bliva slagna av HERREN.
De som låta inviga sig och rena sig till gudstjänst i lustgårdar, anförda av en som står där i mitten, de som äta svinkött och annan styggelse, ja, också möss, de skola allasammans förgås, säger HERREN.
Jag känner deras gärningar och tankar.
Den tid kommer, då jag skall församla alla folk och tungomål; och de skola komma och se min härlighet.
Och jag skall göra ett tecken bland dem; och några av dem som bliva räddade skall jag sända såsom budbärare till hednafolken, till Tarsis, till Pul och Lud, bågskyttfolken, till Tubal och Javan, till havsländerna i fjärran, som icke hava hört något om mig eller sett min härlighet; och de skola förkunna min härlighet bland folken.
Och på hästar och i vagnar och bärstolar och på mulåsnor och dromedarer skola de från alla folk föra alla edra bröder fram till mitt heliga berg i Jerusalem såsom ett spisoffer åt HERREN, säger HERREN, likasom Israels barn i rena kärl föra fram spisoffer till HERRENS hus.
Och jämväl sådana skall jag taga till mina präster, till mina leviter, säger HERREN.
Ty likasom de nya himlar och den nya jord, som jag vill göra, bliva beståndande inför mig, säger HERREN, så skall det ock vara med edra barn och med edert namn.
Och nymånadsdag efter nymånadsdag och sabbatsdag efter sabbatsdag skall det ske, att allt kött kommer och tillbeder inför mig, säger HERREN.
Och man skall gå ut och se med lust, huru de människor, som avföllo från mig, nu ligga där döda; ty deras mask skall icke dö, och deras eld skall icke utsläckas, och de skola vara till vämjelse för allt kött.
Detta är vad som talades av Jeremia, Hilkias son, en av prästerna i Anatot i Benjamins land.
Till honom kom HERRENS ord i Josias, Amons sons, Juda konungs, tid, i hans trettonde regeringsår,
Och sedan i Jojakims, Josias sons, Juda konungs, tid, intill slutet av Sidkias, Josias sons, Juda konungs, elfte regeringsår, då Jerusalems invånare i femte månaden fördes bort i fångenskap.
HERRENS ord kom till mig; han sade:
»Förrän jag danade dig i moderlivet, utvalde jag dig, och förrän du utgick ur modersskötet, helgade jag dig; jag satte dig till en profet för folken.»
Men jag svarade: »Ack Herre HERRE!
Se, jag förstår icke att tala, ty jag är för ung.
Då sade HERREN till mig: »Säg icke: 'Jag är för ung', utan gå åstad vart jag än sänder dig, och tala vad jag än bjuder dig.
Frukta icke för dem; ty jag är med dig och vill hjälpa dig, säger HERREN.»
Och HERREN räckte ut sin hand och rörde vid min mun; och HERREN sade till mig: »Se, jag lägger mina ord i din mun.
Ja, jag sätter dig i dag över folk och riken, för att du skall upprycka och nedbryta, förgöra och fördärva, uppbygga och plantera.»
Och HERRENS ord kom till mig; han sade: »Vad ser du, Jeremia?»
Tag svarade: »Jag ser en gren av ett mandelträd.»
Och HERREN sade till mig: »Du har sett rätt, ty jag skall vaka över mitt ord och låta det gå i fullbordan.»
Och HERRENS ord kom till mig för andra gången; han sade: »Vad ser du?»
Jag svarade: »Jag ser en sjudande gryta; den synes åt norr till.»
Och HERREN sade till mig: »Ja, från norr skall olyckan bryta in över alla landets inbyggare.
Ty se, jag skall kalla på alla folkstammar i rikena norrut, säger HERREN; och de skola komma och resa upp var och en sitt säte vid ingången till Jerusalems portar och mot alla dess murar, runt omkring, och mot alla Juda städer.
Och jag skall gå till rätta med dem för all deras ondska, därför att de hava övergivit mig och tänt offereld åt andra gudar och tillbett sina händers verk.
Så omgjorda nu du dina länder, och stå upp och tala till dem allt vad Jag bjuder dig.
Var icke förfärad för dem, på det att jag icke må låta vad förfärligt är komma över dig inför dem.
Ty se, jag själv gör dig i dag till en fast stad och till en järnpelare och en kopparmur mot hela landet, mot Juda konungar, mot dess furstar, mot dess präster och mot det meniga folket,
så att de icke skola bliva dig övermäktiga, om de vilja strida mot dig; ty jag är med dig, säger HERREN, och jag vill hjälpa dig.»
Och HERRENS ord kom till mig; han sade:
Gå åstad och predika för Jerusalem och säg: Så säger HERREN: Jag kommer ihåg, dig till godo, din ungdoms kärlek, huru du älskade mig under din brudtid, huru du följde mig i öknen, i landet där man intet sår.
Ja, en HERRENS heliga egendom är Israel, förstlingen av hans skörd; alla som vilja äta därav ådraga sig skuld, olycka kommer över dem, säger HERREN.
Hören HERRENS ord, I av Jakobs hus, I alla släkter av Israels hus.
Så säger HERREN: Vad orätt funno edra fäder hos mig, eftersom de gingo bort ifrån mig och följde efter fåfängliga avgudar och bedrevo fåfänglighet?
De frågade icke: »Var är HERREN, han som förde oss upp ur Egyptens land, han som ledde oss i öknen, det öde och oländiga landet, torrhetens och dödsskuggans land, det land där ingen vägfarande färdades, och där ingen människa bodde?»
Och jag förde eder in i det bördiga landet, och I fingen äta av dess frukt och dess goda.
Men när I haden kommit ditin, orenaden I mitt land och gjorden min arvedel till en styggelse.
Prästerna frågade icke: »Var är HERREN?»
De som hade lagen om händer ville icke veta av mig, och herdarna avföllo från mig; profeterna profeterade i Baals namn och följde efter sådana som icke kunde hjälpa.
Därför skall jag än vidare gå till rätta med eder, säger HERREN, ja, ännu med edra barnbarn skall jag gå till rätta.
Dragen bort till kittéernas öländer och sen efter, sänden bud till Kedar och forsken noga efter; sen till, om något sådant där har skett.
Har väl något hednafolk bytt bort sina gudar?
Och dock äro dessa inga gudar.
Men mitt folk har bytt bort sin ära mot en avgud som icke kan hjälpa.
Häpnen häröver, I himlar; förskräckens och bäven storligen, säger HERREN.
Ty mitt folk har begått en dubbel synd: mig hava de övergivit, en källa med friskt vatten, och de hava gjort sig brunnar, usla brunnar, som icke hålla vatten.
Är väl Israel en träl eller en hemfödd slav, eftersom han så har lämnats till plundring?
Lejon ryta mot honom, de låta höra sitt skri.
De göra hans land till en ödemark, hans städer brännas upp, så att ingen kan bo i dem.
Till och med Nofs och Tapanhes' barn avbeta dina berg.
Men är det ej du själv som vållar dig detta, därmed att du övergiver HERREN din Gud, när han vill leda dig på den rätta vägen?
Varför vill du nu gå till Egypten och dricka av Sihors vatten?
Och varför vill du gå till Assyrien och dricka av flodens vatten?
Det är din ondska som bereder dig tuktan, det är din avfällighet som ådrager dig straff.
Märk därför och besinna vilken olycka och sorg det har med sig att du övergiver HERREN, din Gud, och icke vill frukta mig, säger Herren, HERREN Sebaot.
Ty för länge sedan bröt du sönder ditt ok och slet av dina band och sade: »Jag vill ej tjäna.»
Och på alla höga kullar och under alla gröna träd lade du dig ned för att öva otukt.
Jag hade ju planterat dig såsom ett ädelt vinträd av alltigenom äkta art; huru har du då kunnat förvandlas för mig till vilda rankor av ett främmande vinträd?
Ja, om du ock tvår dig med lutsalt och tager än så mycken såpa, så förbliver dock din missgärning oren inför mig, säger Herren, HERREN.
Huru kan du säga: »Jag har ej orenat mig, jag har icke följt efter Baalerna»?
Besinna vad du har bedrivit i dalen, ja, betänk vad du har gjort.
Du är lik ett ystert kamelsto, som löper hit och dit.
Du är lik en vildåsna, fostrad i öknen, en som flåsar i sin brunst, och vars brånad ingen kan stävja; om någon vill till henne, behöver han ej löpa sig trött; när hennes månad kommer, träffar man henne.
Akta din fot, så att den icke tappar skon, och din strupe, så att den ej bliver torr av törst.
Men du svarar: »Du mödar dig förgäves.
Nej, jag älskar de främmande, och efter dem vill jag följa.»
Såsom tjuven står där med skam, när han ertappas, så skall Israels hus komma på skam, med sina konungar, och furstar, med sina präster och profeter,
dessa som säga till trästycket: »Du är min fader», och säga till stenen: »Du har fött mig.»
Ty de vända ryggen till mig och icke ansiktet; men när olycka är på färde, ropa de: »Upp och fräls oss!»
Var äro då dina gudar, de som du gjorde åt dig?
Må de stå upp.
Kunna de frälsa dig i din olyckas tid?
Ty så många som dina städer äro, så många hava dina gudar blivit, du Juda.
Huru kunnen I gå till rätta med mig?
I haven ju alla avfallit från mig, säger HERREN.
Förgäves har jag slagit edra barn; de hava icke velat taga emot tuktan.
Edert svärd har förtärt edra profeter, såsom vore det ett förhärjande lejon.
Du onda släkte, giv akt på HERRENS ord.
Har jag då för Israel varit en öken eller ett mörkrets land, eftersom mitt folk säger: »Vi hava gjort oss fria, vi vilja ej mer komma till dig»?
Icke förgäter en jungfru sina smycken eller en brud sin gördel?
Men mitt folk har förgätit mig sedan urminnes tid.
Huru skickligt går du icke till väga, när du söker älskog!
Därför har du ock blivit förfaren på det ondas vägar.
Ja, på dina mantelflikar finner man blod av arma och oskyldiga, som du har dödat, icke därför att de ertappades vid inbrott, nej, därför att din håg står till allt sådant.
Och dock säger du: »Jag går fri ifrån straff; hans vrede mot mig har förvisso upphört.»
Nej, jag vill gå till rätta med dig, om du än säger: »Jag har icke syndat.»
Varför har du nu så brått att vandra åstad på en annan väg?
Också med Egypten skall du komma på skam, likasom du kom på skam med Assyrien.
Också därifrån skall du få gå din väg, med händerna på huvudet.
Ty HERREN förkastar dem som du förlitar dig på, och du skall icke bliva lyckosam med dem.
Det är sagt: Om en man skiljer sig från sin hustru, och hon så går bort ifrån honom och bliver en annan mans hustru, icke får han då åter komma tillbaka till henne?
Bleve icke då det landet ohelgat?
Och du, som har bedrivit otukt med så många älskare, du vill ändå få komma tillbaka till mig! säger HERREN.
Lyft upp dina ögon till höjderna och se: var lät du icke skända dig?
Vid vägarna satt du och spejade efter dem, såsom en arab i öknen, och ohelgade landet genom din otukt och genom din ondska.
Väl blevo regnskurarna förhållna, och intet vårregn föll; men du hade en äktenskapsbryterskas panna, du ville icke blygas.
Och ändå har du nyss ropat till mig: »Min fader!», Min ungdoms vän är du!»
»Skulle han kunna behålla vrede evinnerligen, skulle han framhärda så för alltid?»
Så talar du och gör dock vad ont är, ja, fullbordar det ock.
Och HERREN sade till mig i konung Josias tid: Har du sett vad Israel, den avfälliga kvinnan, har gjort?
Hon gick upp på alla höga berg och bort under alla gröna träd och bedrev där otukt.
Och jag tänkte att sedan hon hade gjort allt detta, skulle hon vända tillbaka till mig.
Men hon vände icke tillbaka.
Och hennes syster Juda, den trolösa kvinnan, såg det.
Och jag såg, att fastän jag hade skilt mig från Israel, den avfälliga, och givit henne skiljebrev just för hennes äktenskapsbrotts skull, så skrämdes dock hennes syster Juda den trolösa, icke därav, utan gick likaledes åstad och bedrev otukt
och ohelgade så landet genom sin lättfärdiga otukt, i det hon begick äktenskapsbrott med sten och trä.
Ja, oaktat allt detta vände hennes syster Juda, den trolösa, icke tillbaka till mig av fullt hjärta, utan allenast med skrymteri, säger HERREN.
Och HERREN sade till mig: Israel, den avfälliga, har bevisat sig rättfärdigare än Juda, den trolösa.
Gå bort och predika så norrut och säg: Vänd om, Israel, du avfälliga, säger HERREN, så vill jag icke längre med ogunst se på eder; ty jag är nådig, säger HERREN, jag behåller icke vrede evinnerligen.
Allenast må du besinna din missgärning, att du har varit avfällig från HERREN, din Gud, och lupit hit och dit till främmande gudar under alla gröna träd; ja, I haven icke velat höra min röst, säger HERREN.
Vänden om, I avfälliga barn, säger HERREN, ty jag är eder rätte herre; så vill jag hämta eder, en från var stad och två från var släkt, och föra eder till Sion.
Och jag vill giva eder herdar efter mitt hjärta, och de skola föra eder i bet med förstånd och insikt.
Och det skall ske, att när I på den tiden föröken eder och bliven fruktsamma i landet, säger HERREN, då skall man icke mer tala om HERRENS förbundsark eller tänka på den; man skall icke komma ihåg den eller sakna den, och man skall icke göra någon ny sådan.
Utan på den tiden skall man kalla Jerusalem »HERRENS tron»; och dit skola församla sig alla hednafolk, till HERRENS namn i Jerusalem.
Och de skola icke mer vandra efter sina onda hjärtans hårdhet.
På den tiden skall Juda hus gå till Israels hus, och tillsammans skola de komma från nordlandet in i det land som jag gav edra fäder till arvedel.
Jag tänkte: »Vilken plats skall jag ej förläna dig bland barnen, och vilket ljuvligt land skall jag icke giva dig, den allra härligaste arvedel bland folken!»
Och jag tänkte: »Då skolen I kalla mig fader och icke mer vika bort ifrån mig.»
Men såsom när en hustru är trolös mot sin make, så haven I av Israels hus varit trolösa mot mig, säger HERREN.
Därför höras rop på höjderna, gråt och böner av Israels barn; ty de hava gått på förvända vägar och förgätit HERREN, sin Gud.
Så vänden nu om, I avfälliga barn, så vill jag hela eder från edert avfall.
Ja se, vi komma till dig, ty du är HERREN, vår Gud.
Sannerligen, bedrägligt var vårt hopp till höjderna, blott tomt larm gåvo oss bergen.
Sannerligen, det är hos HERREN, vår Gud, som frälsning finnes för Israel.
Men skändlighetsguden har förtärt frukten av våra fäders arbete, allt ifrån vår ungdom, deras får och fäkreatur, deras söner och döttrar.
Så vilja vi nu ligga här i vår skam, och blygd må hölja oss.
Ty mot HERREN, vår Gud, hava vi syndat, vi och våra fäder, ifrån vår ungdom ända till denna dag; vi hava icke velat höra HERRENS, vår Guds, röst.
om du omvänder dig, Israel, säger HERREN, skall du få vända tillbaka till mig; och om du skaffar bort dina styggelser från min åsyn, skall du slippa vandra flyktig omkring.
Då skall du svärja i sanning, rätt och rättfärdighet: »Så sant HERREN lever», och hednafolken skola välsigna sig i honom och berömma sig av honom.
Ja, så säger HERREN till Juda män och till Jerusalem: Bryten eder ny mark, och sån ej bland törnen.
Omskären eder åt HERREN; skaffen bort edert hjärtas förhud, I Juda män och I Jerusalems invånare.
Eljest skall min vrede bryta fram såsom en eld och brinna så, att ingen kan utsläcka den, för edert onda väsendes skull.
Förkunnen i Juda, kungören i Jerusalem och påbjuden, ja, stöten i basun i landet, ropen ut med hög röst och sägen: »Församlen eder och låt oss fly in i de befästa städerna.»
Resen upp ett baner som visar åt Sion, bärgen edert gods och dröjen icke ty jag skall låta olycka komma från norr, med stor förstöring.
Ett lejon drager fram ur sitt snår och en folkfördärvare bryter upp, han går ut ur sin boning, för att göra ditt land till en ödemark; då bliva dina städer förstörda, så att ingen kan bo i dem.
Så höljen eder nu i sorgdräkt, klagen och jämren eder, ty HERRENS vredes glöd upphör icke över oss.
På den tiden, säger HERREN, skall det vara förbi med konungens och furstarnas mod, och prästerna skola bliva förfärade och profeterna stå häpna.
Men jag sade: »Ack Herre, HERRE, svårt bedrog du sannerligen detta folk och Jerusalem, då du sade: »Det skall gå eder väl.»
Svärdet är ju nära att taga vårt liv.
På den tiden skall det sägas om detta folk och om Jerusalem: En brännande vind från höjderna i öknen kommer emot dottern mitt folk, icke en sådan vind som passar, när man kastar säd eller rensar korn;
nej, en våldsammare vind än som så låter jag komma.
Ja, nu vill jag gå till rätta med dem!
Se, såsom ett moln kommer han upp och såsom en stormvind äro hans vagnar; hans hästar äro snabbare än örnar, ve oss, vi äro förlorade!
Så två nu ditt hjärta rent från ondska, Jerusalem, för att du må bliva frälst.
Huru länge skola fördärvets tankar bo i ditt bröst?
Från Dan höres ju en budbärare ropa, och från Efraims bergsbygd en som bådar fördärv.
Förkunnen för folken, ja, kungören över Jerusalem att en belägringshär kommer ifrån fjärran land och häver upp sitt rop mot Juda städer.
Såsom väktare kring ett åkerfält samla de sig runt omkring henne, därför att hon har varit gensträvig mot mig, säger HERREN.
Ja, ditt eget leverne och dina egna varningar vålla dig detta; det är din ondskas frukt att det bliver dig så bittert, och att plågan träffar dig ända in i hjärtat.
I mitt innersta våndas jag, i mitt hjärtas djup.
Mitt hjärta klagar i mig, jag kan icke tiga, ty basunljud hör du, min själ, och krigiskt härskri.
Olycka efter olycka ropas ut, ja, hela landet bliver förött; plötsligt bliva mina hyddor förödda, i ett ögonblick mina tält.
Huru länge skall jag se stridsbaneret och höra basunljud?
Ja, mitt folk är oförnuftigt, de vilja ej veta av mig.
De äro dåraktiga barn och hava intet förstånd.
Visa äro de till att göra vad ont är, men att göra vad gott är förstå de ej.
Jag såg på jorden, och se, den var öde och tom, och upp mot himmelen, och där lyste intet ljus.
Jag såg på bergen, och se, de bävade, och alla höjder vacklade.
Jag såg mig om, och då fanns där ingen människa, och alla himmelens fåglar hade flytt bort.
Jag såg mig om, och då var det bördiga landet en öken, och alla dess städer voro nedbrutna, för HERRENS ansikte, för hans vredes glöd,
Ty så säger HERREN: Hela landet skall bliva en ödemark, om jag än ej alldeles vill göra ände därpå.
Därför sörjer jorden, och himmelen därovan kläder sig i sorgdräkt, därför att jag så har talat och beslutit och ej kan ångra det eller taga det tillbaka.
För larmet av ryttare och bågskyttar tager hela staden till flykten.
Man giver sig in i skogssnåren och upp bland klipporna.
Alla städer äro övergivna, ingen människa bor mer i dem.
Vad vill du göra i din förödelse?
Om du än kläder dig i scharlakan, om du än pryder dig med gyllene smycken om du än söker förstora dina ögon genom smink, så gör du dig dock skön förgäves.
Dina älskare förakta dig, ja, de stå efter ditt liv.
Ty jag hör rop såsom av en barnaföderska, nödrop såsom av en förstföderska.
Det är dottern Sion som ropar; hon flämtar, hon räcker ut sina händer: »Ack, ve mig!
I mördares våld försmäktar min själ.»
Gån omkring på gatorna i Jerusalem, och sen till och given akt; söken på dess torg om I finnen någon, om där är någon som gör rätt och beflitar sig om sanning; då vill jag förlåta staden.
Men säga de än: »Så sant HERREN lever», så svärja de dock falskt.
HERRE, är det ej sanning dina ögon söka?
Du slog dem, men de kände ingen sveda.
Du förgjorde dem, men de ville ej taga emot tuktan.
De gjorde sina pannor hårdare än sten, de ville icke omvända sig.
Då tänkte jag: »Detta är allenast de ringa i folket; de äro dåraktiga, ty de känna icke HERRENS väg, sin Guds rätt.
Jag vill nu gå till de stora och tala med dem; de måste ju känna HERRENS väg, sin Guds rätt.»
Men ock dessa hade alla brutit sönder oket och slitit av banden.
Därför bliva de slagna av lejonet från skogen och fördärvade av vargen från hedmarken; pantern lurar vid deras städer, och envar som vågar sig ut därifrån bliver ihjälriven.
Ty många äro deras överträdelser och talrika deras avfällighetssynder.
Huru skulle jag då kunna förlåta dig?
Dina barn hava ju övergivit mig och svurit vid gudar som icke äro gudar.
Jag gav dem allt till fyllest, men de blevo mig otrogna och samlade sig i skaror till skökohuset.
De likna välfödda, ystra hästar; de vrenskas var och en efter sin nästas hustru.
Skulle jag icke för sådant hemsöka dem? säger HERREN.
Och skulle icke min själ hämnas på ett sådant folk som detta är?
Stormen då hennes murar och för stören dem, dock utan att alldeles göra ände på henne.
Riven bort hennes vinrankor, de äro ju icke HERRENS.
Ty både Israels hus och Juda hus hava varit mycket trolösa mot mig, säger HERREN.
De hava förnekat HERREN och sagt: »Han betyder intet.
Olycka skall icke komma över oss, svärd och hunger skola vi icke se.
Men profeterna skola försvinna såsom en vind, och han som säges tala är icke i dem; dem själva skall det så gå.»
Därför säger HERREN, härskarornas Gud: Eftersom I fören ett sådant tal, se, därför skall jag göra mina ord i din mun till en eld, och detta folk till ved, och elden skall förtära dem.
Se, jag skall låta komma över eder, I av Israels hus, ett folk ifrån fjärran land, säger HERREN, ett starkt folk, ett urgammalt folk, ett folk vars tungomål du icke känner, och vars tal du icke förstår.
Deras koger är en öppen grav; de äro allasammans hjältar.
De skola förtära din skörd och ditt bröd, de skola förtära dina söner och döttrar, de skola förtära dina får och fäkreatur, de skola förtära dina vinträd och fikonträd.
Dina befästa städer, som du förlitar dig på, dem skola de förstöra med svärd.
Dock vill jag på den tiden, säger HERREN, icke alldeles göra ände på eder.
Och om I då frågen: »Varför har HERREN, vår Gud, gjort oss allt detta?», så skall du svara dem: »Såsom I haven övergivit mig och tjänat främmande gudar i edert eget land, så skolen I nu få tjäna främlingar i ett land som icke är edert.»
Förkunnen detta i Jakobs hus, kungören det i Juda och sägen:
Hör detta, du dåraktiga och oförståndiga folk, I som haven ögon, men icke sen, I som haven öron, men icke hören.
Skullen I icke frukta mig, säger HERREN, skullen I icke bäva för mig, for mig som har satt stranden till en damm for havet, till en evärdlig gräns, som det icke kan överskrida, så att dess böljor, huru de än svalla, ändå intet förmå, och huru de än brusa, likväl icke kunna överskrida den?
Men detta folk har ett gensträvigt och upproriskt hjärta; de hava avfallit och gått sin väg.
De sade icke i sina hjärtan: »Låtom oss frukta HERREN, vår Gud, honom som giver regn i rätt tid, både höst och vår, och som ständigt beskär oss de bestämda skördeveckorna.»
Edra missgärningar hava nu fört dessa i olag, och edra synder hava förhållit för eder detta goda.
Ty bland mitt folk finnas ogudaktiga människor: de ligga i försåt, likasom fågelfängaren ligger på lur, de sätta ut giller till att fånga människor.
Såsom när en bur är full av fåglar, så äro deras hus fulla av svek.
Därigenom hava de blivit så stora och rika; de hava blivit feta och skinande.
För sina ogärningar veta de icke av någon gräns, de hålla icke rätten vid makt, icke den faderlöses rätt, till att främja den; och i den fattiges sak fälla de icke rätt dom.
Skulle jag icke för sådant hemsöka dem? säger HERREN.
Skulle icke min själ hämnas på ett sådant folk som detta är?
Förfärliga och gruvliga ting ske i landet.
Profeterna profetera lögn, och prästerna styra efter deras råd; och mitt folk vill så hava det.
Men vad skolen I göra, när änden på detta kommer?
Bärgen edert gods ut ur Jerusalem, I Benjamins barn, stöten i basun i Tekoa, och resen upp ett högt baner ovanför Bet-Hackerem; ty en olycka hotar från norr, med stor förstöring.
Hon som är så fager och förklemad, dottern Sion, henne skall jag förgöra.
Herdar skola komma över henne med sina hjordar; de skola slå upp sina tält runt omkring henne, avbeta var och en sitt stycke.
Ja, invigen eder till strid mot henne. »Upp, låt oss draga åstad, medan middagsljuset varar!
Ack att dagen redan lider till ända!
Ack att aftonens skuggor förlängas!
Välan, så låt oss draga ditupp om natten och förstöra hennes palatser.»
Ty så säger HERREN Sebaot: Fällen träd och kasten upp vallar emot Jerusalem.
Hon är staden som skall hemsökas, hon som i sig har idel förtryck
Likasom en brunn låter vatten välla fram, så låter hon ondska framvälla.
Våld och förödelse hör man där, sår och slag äro beständigt inför min åsyn.
Låt varna dig, Jerusalem, så att min själ ej vänder sig ifrån dig, så att jag icke gör dig till en ödemark, till ett obebott land.
Så säger HERREN Sebaot: En efterskörd, likasom på ett vinträd, skall man hålla på kvarlevan av Israel.
Räck ut din hand åter och åter, såsom när man plockar av druvor från rankorna.
Men inför vem skall jag tala och betyga för att bliva hörd?
Se, deras öron äro oomskurna, så att de icke kunna höra.
Ja, HERRENS ord har blivit till smälek bland dem; de hava intet behag därtill.
Därför är jag uppfylld av HERRENS vrede, jag förmår icke hålla den inne.
Utgjut den över barnen på gatan och över alla de unga männens samkväm; ja, både man och kvinna skola drabbas därav, jämväl den gamle och den som har fyllt sina dagars mått.
Och deras hus skola gå över i främmandes ägo så ock deras åkrar och deras hustrur, ty jag vill uträcka min hand mot landets inbyggare, säger HERREN.
Ty alla, både små och stora, söka där orätt vinning, och både profeter och präster fara allasammans med lögn,
de taga det lätt med helandet av mitt folks skada; de säga: »Allt står väl till, allt står väl till», och dock står icke allt väl till.
De skola komma på skam, ty de övade styggelse.
Likväl känna de alls icke någon skam och veta icke av någon blygsel.
Därför skola de falla bland de andra; när min hemsökelse träffar dem, skola de komma på fall, säger HERREN,
Så sade HERREN: »Ställen eder vid vägarna och sen till, och frågen efter forntidens stigar, frågen vilken väg som är den goda vägen, och vandren på den, så skolen I finna ro för edra själar.»
Men de svarade: »Vi vilja icke vandra på den.»
Och när jag då satte väktare över eder och sade: »Akten på basunens ljud», svarade de: »Vi vilja icke akta därpå.»
Hören därför, I hednafolk, och märk, du menighet, vad som sker bland dem.
Ja hör, du jord: Se, jag skall låta olycka komma över detta folk, såsom en frukt av deras anslag, eftersom de icke akta på mina ord, utan förkasta min lag.
Vad frågar jag efter rökelse, komme den ock från Saba, eller efter bästa kalmus ifrån fjärran land?
Edra brännoffer täckas mig icke, och edra slaktoffer behaga mig icke.
Därför säger HERREN så: Se, jag skall lägga stötestenar för detta folk; och genom dem skola både fader och söner komma på fall, den ene borgaren skall förgås med den andre.
Så säger HERREN: Se, ett folk kommer från nordlandet, ett stort folk reser sig vid jordens yttersta ända.
De föra båge och lans, de äro grymma och utan förbarmande.
Dånet av dem är såsom havets brus, och på sina hästar rida de fram, rustade såsom kämpar till strid, mot dig, du dotter Sion.
När vi höra ryktet om dem, sjunka våra händer ned, ängslan griper oss, ångest lik en barnaföderskas.
Gå icke ut på marken, och vandra ej på vägen, ty fienden bär svärd; skräck från alla sidor!
Du dotter mitt folk, höll dig i sorgdräkt, vältra dig i aska, höj sorgelåt likasom efter ende sonen, och håll bitter dödsklagan; ty plötsligt kommer förhärjaren över oss.
Jag har satt dig till en proberare i mitt folk -- såväl som till ett fäste -- på det att du må lära känna och pröva deras väg.
De äro allasammans avfälliga och gensträviga, de gå med förtal, de äro koppar och järn, allasammans äro de fördärvliga människor.
Blåsbälgen pustar, men ur elden kommer allenast bly fram; allt luttrande är förgäves, slagget bliver ändå icke frånskilt.
»Ett silver som må kastas bort», så kan man kalla dem, ty HERREN har förkastat dem.
Detta är det ord som kom till Jeremia från HERREN; han sade:
Ställ dig i porten till HERRENS hus, och predika där detta ord och säg: Hören HERRENS ord, I alla av Juda, som gån in genom dessa portar för att tillbedja HERREN.
Så säger HERREN Sebaot, Israels Gud: Bättren edert leverne och edert väsende, så vill jag låta eder bo kvar på denna plats.
Förliten eder icke på lögnaktigt tal, när man säger: »Här är HERRENS tempel, HERRENS tempel, HERRENS tempel!»
Nej, om I bättren edert leverne och edert väsende, om I dömen rätt mellan man och man,
om I upphören att förtrycka främlingen, den faderlöse och änkan, att utgjuta oskyldigt blod på denna plats och att följa efter andra gudar, eder själva till olycka,
då vill jag för evärdliga tider låta eder bo på denna plats, i det land som jag har givit åt edra fäder.
Men se, I förliten eder på lögnaktigt tal, som icke kan hjälpa.
Huru är det?
I stjälen, mörden och begån äktenskapsbrott, I svärjen falskt, I tänden offereld åt Baal och följen efter andra gudar, som I icke kännen;
sedan kommen I hit och träden fram inför mitt ansikte i detta hus, som är uppkallat efter mitt namn, och sägen: »Med oss är ingen nöd» -- för att därefter fortfara med alla dessa styggelser.
Hållen I det då för en rövarkula, detta hus, som är uppkallat efter mitt namn?
Ja, sannerligen, också jag anser det så, säger HERREN.
Gån bort till den plats i Silo, där jag först lät mitt namn bo, och sen huru jag har gjort med den, för mitt folk Israels ondskas skull.
Och eftersom I haven gjort alla dessa gärningar, säger HERREN, och icke haven velat höra, fastän jag titt och ofta har talat till eder, och icke haven velat svara, fastän jag har ropat på eder,
därför vill jag nu med detta hus, som är uppkallat efter mitt namn, och som I förliten eder på, och med denna plats, som jag har givit åt eder och edra fäder, göra såsom jag gjorde med Silo.
Och jag skall kasta eder bort ifrån mitt ansikte, såsom jag har bortkastat alla edra bröder all Efraims släkt.
Så må du nu icke bedja för detta folk eller frambära någon klagan och förbön för dem eller lägga dig ut för dem hos mig, ty jag vill icke höra dig.
Ser du icke vad de göra i Juda städer och på Jerusalems gator?
Barnen samla tillhopa ved, fäderna tända upp eld och kvinnorna knåda deg, allt för att baka offerkakor åt himmelens drottning; och drickoffer utgjuta de åt andra gudar, mig till sorg.
Men är det då mig som de bereda sorg därmed, säger HERREN, och icke fastmer sig själva, så att de komma på skam?
Därför säger Herren, HERREN så: Se, min vrede och förtörnelse skall utgjuta sig över denna plats, över både människor och djur, över både träden på marken och frukten på jorden; och den skall brinna och icke bliva utsläckt.
Så säger HERREN Sebaot, Israels Gud: Läggen edra brännoffer tillhopa med edra slaktoffer och äten så kött.
Ty på den tid då jag förde edra fäder ut ur Egyptens land gav jag dem icke någon befallning eller något bud angående brännoffer och slaktoffer;
utan detta var det bud jag gav dem: »Hören min röst, så vill jag vara eder Gud, och I skolen vara mitt folk; och vandren i allt på den väg som jag bjuder eder, på det att det må gå eder väl.»
Men de ville icke höra eller böja sitt öra till mig, utan vandrade efter sina egna rådslag, i sina onda hjärtans hårdhet, och veko tillbaka i stället för att gå framåt.
Allt ifrån den dag då edra fäder drogo ut ur Egyptens land ända till nu har jag dag efter dag, titt och ofta, sänt till eder alla mina tjänare profeterna.
Men man ville icke höra mig eller böja sitt öra till mig; de voro hårdnackade och gjorde ännu mer ont än deras fäder.
Och om du än säger dem allt detta, så skola de dock icke höra dig; och om du än ropar till dem, så skola de dock icke svara dig.
Säg därför till dem: »Detta är det folk som icke vill höra HERRENS, sin Guds, röst eller taga emot tuktan.
Sanningen är försvunnen och utrotad ur deras mun.»
Skär av dig ditt huvudhår och kasta det bort, och stäm upp en klagosång på höjderna.
Ty HERREN har förkastat och förskjutit detta släkte, som har uppväckt hans vrede.
Juda barn hava ju gjort vad ont är i mina ögon, säger HERREN; de hava satt upp sina styggelser i det hus som är uppkallat efter mitt namn, och de hava så orenat det.
Och Tofethöjderna i Hinnoms sons dal hava de byggt upp, för att där uppbränna sina söner och döttrar i eld, fastän jag aldrig har bjudit eller ens tänkt mig något sådant.
Se, därför skola dagar komma, säger HERREN, då man icke mer skall säga »Tofet» eller »Hinnoms sons dal», utan »Dråpdalen», och då man skall begrava i Tofet, därför att ingen annan plats finnes.
Ja, detta folks döda kroppar skola bliva mat åt himmelens fåglar och markens djur, och ingen skall skrämma bort dem.
Och i Juda städer och på Jerusalems gator skall jag göra slut på fröjderop och glädjerop, på rop för brudgum och rop för brud, ty landet skall bliva ödelagt.
på den tiden, säger HERREN, skall man kasta Juda konungars och furstars ben, och prästernas och profeternas ben, och Jerusalems invånares ben ut ur deras gravar
och kringströ dem inför solen och månen och himmelens hela härskara, som de hava älskat, tjänat och efterföljt, sökt och tillbett; man skall icke sedan samla dem tillhopa eller begrava dem, utan de skola bliva gödsel på marken.
Och alla kvarblivna, de som lämnas kvar av detta onda släkte, skola hellre vilja dö än leva, vilka än de orter må vara, dit dessa kvarlämnade bliva fördrivna av mig, säger HERREN Sebaot.
Du skall ock säga till dem: Så säger HERREN: Om någon faller, står han ju upp igen; om någon går bort, vänder han ju tillbaka.
Varför går det då bort i beständig avfällighet, detta folk i Jerusalem?
Varför hålla de fast vid sitt svek och vilja icke vända tillbaka?
Jag har givit akt och hört huru de tala vad orätt är; ingen enda finnes, som ångrar sin ondska, ingen säger: »Vad har jag gjort!»
Alla löpa de bort, lika hästar som rusa åstad i striden.
Till och med hägern under himmelen känner ju sin bestämda tid, och turturduvan, svalan och tranan taga i akt tiden för sin återkomst; mitt folk däremot känner ej HERRENS rätter.
Huru kunnen I då säga: »Vi äro visa och hava HERRENS lag ibland oss»?
Icke så, de skriftlärdes lögnpenna har förvandlat den i lögn.
Sådana visa skola komma på skam, komma till korta och bliva snärjda.
De hava ju förkastat HERRENS ord, vari äro de då visa?
Så skall jag nu giva deras hustrur åt andra och deras åkrar åt erövrare Ty alla, både små och stora, söka orätt vinning; både profeter och präster fara allasammans med lögn,
de taga det lätt med helandet av dottern mitt folks skada; de säga: »Allt står väl till, allt står väl till», och dock står icke allt väl
De skola komma på skam, övade styggelse.
Likväl känna de alls icke skam och veta icke av att blygas.
Därför skola de falla bland de andra; när hemsökelsen träffar dem, skola de komma på fall, säger HERREN.
Jag skall bortrycka och förgöra dem, säger HERREN.
Inga druvor växa på vinträden, och inga fikon på fikonträden, utan till och med löven äro vissnade: De bud jag gav dem överträda de.
Varför sitta vi här stilla?
Församlen eder och låt oss fly in i de befästa städerna och förgås där; ty HERREN, vår Gud, vill förgöra oss, han giver oss gift att dricka därför att vi syndade mot HERREN.
V bida efter frid, men intet gott kommer, efter en tid då vi skulle bliva helade, men se, förskräckelse kommer.
Från Dan hör man frustandet av hans hästar; för hans hingstars gnäggande bävar hela landet.
De komma och förtära landet med allt vad däri är, staden med dem som bo däri.
Ty se, jag sänder emot eder ormar, basilisker, mot vilka ingen besvärjelse hjälper, och de skola stinga eder, säger HERREN.
Var skall jag finna vederkvickelse i min sorg?
Mitt hjärta är sjukt i mig.
Hör, dottern mitt folk ropar i fjärran land: »Finnes då icke HERREN i Sion?
Är dennes konung icke mer där?»
Ja, varför hava de förtörnat mig med sina beläten, med sina främmande avgudar?
Skördetiden är förbi, sommaren är till ända, och ingen frälsning har kommit oss till del.
Jag är förkrossad, därför att dottern mitt folk så krossas, jag går sörjande, häpnad har gripit mig.
Finnes då ingen balsam i Gilead, finnes ingen läkare där?
Eller varför bliver dottern mitt folk icke helad från sina sår?
Ack att mitt huvud vore en vattenbrunn och mina ögon en tårekälla, så att jag kunde gråta dag och natt över de slagna hos dottern mitt folk!
Ack att jag hade ett härbärge i öknen, så att jag kunde övergiva mitt folk och draga bort ifrån dem!
Ty de äro allasammans äktenskapsbrytare, en församling av trolösa.
Sin tungas båge spänna de till att avskjuta lögner, och till sanning bruka de icke sin makt i landet.
Nej, de gå från ogärning till ogärning, men mig vilja de ej veta av, säger HERREN.
Var och en tage sig till vara för sin vän, och ingen förlite sig på någon sin broder; ty den ene brodern gör allt för att bedraga den andre, och den ene vännen går omkring och förtalar den andre.
Var och en handlar svikligt mot sin vän, och ingen talar vad sant är; de öva sina tungor i att tala lögn de arbeta sig trötta med att göra illa.
Du bor mitt ibland falskhet; i sin falskhet vilja de ej veta av mig, säger HERREN.
Därför säger HERREN Sebaot så.
Se, jag måste luttra och pröva dem; ty vad annat kan jag göra, då nu dottern mitt folk är sådan?
Deras tunga är en mördande pil; vad den talar är svek.
Med munnen tala de vänligt till sin nästa, men i hjärtat lägga de försåt för honom.
Skulle jag icke för sådant hemsöka dem? säger HERREN.
Skulle icke min själ hämnas på ett sådant folk som detta är?
Över bergen vill jag gråta och sjunga sorgesång; jag vill höja klagosång över betesmarkerna i öknen.
Ty de äro förbrända, så att ingen går där fram och inga läten av boskap där höras; både himmelens fåglar och fyrfotadjuren hava flytt och äro borta.
Jag skall göra Jerusalem till en stenhop, till en boning för schakaler, och Juda städer till en ödemark, där ingen bor.
Vem är en vis man, så att han förstår detta?
Och till vem har HERRENS mun talat, så att han kan förklara detta: varför landet har blivit så fördärvat, förbränt såsom en öken, där ingen går fram?
Och HERREN svarade: Jo, därför att de hava övergivit min lag, den som jag förelade dem, och icke hava hört min röst och vandrat efter den
utan vandrat efter sina egna hjärtans hårdhet och efterföljt Baalerna, såsom deras fader lärde dem.
Därför säger HERREN Sebaot, Israels Gud, så: Se, jag skall giva detta folk malört att äta och gift att dricka.
Och jag skall förströ dem bland folk som varken de eller deras fäder hava känt, och skall sända svärdet efter dem, till dess att jag har gjort ände på dem.
Så säger HERREN Sebaot: Given akt; tillkallen gråterskor, för att de må komma, och sänden efter förfarna kvinnor, och låten dem komma.
Låten dem med hast stämma upp sorgesång över oss, så att våra ögon flyta i tårar och vatten strömmar från våra ögonlock.
Ty sorgesång höres ljuda från Sion: Huru har ej förstörelse drabbat oss!
Vi hava kommit illa på skam, vi måste ju övergiva landet, ty våra boningar hava de slagit ned.
Ja, hören, I kvinnor, HERRENS ord, och edert öra fatte hans muns tal.
Lären edra döttrar sorgesång; ja, lären varandra klagosång.
Ty döden stiger in genom vara fönster, han kommer in i våra palats; han utrotar barnen från gatan och ynglingarna från torgen.
Ja, tala: Så säger HERREN: Och människornas döda kroppar ligga såsom gödsel på marken och såsom kärvar efter skördemannen, vilka ingen samlar upp.
Så säger HERREN: Den vise berömme sig icke av sin vishet, den starke berömme sig icke av sin styrka, den rike berömme sig icke av sin rikedom.
Nej, den som vill berömma sig, han berömme sig därav att han har förstånd till att känna mig: att jag är HERREN, som gör nåd, rätt och rättfärdighet på jorden.
Ty till sådana har jag behag, säger HERREN.
Se, dagar skola komma, säger HERREN, då jag skall hemsöka alla omskurna som dock äro oomskurna:
Egypten, Juda, Edom, Ammons barn, Moab och alla ökenbor med kantklippt hår.
Ty hednafolken äro alla oomskurna, och hela Israels hus har ett oomskuret hjärta.
Hören det ord som HERREN talar till eder, I av Israels hus.
Så säger HERREN:
I skolen icke vänja eder vid hedningarnas sätt och icke förfäras för himmelens tecken, därför att hedningarna förfäras för dem.
Ty vad folken predika är fåfängliga avgudar.
Se, av ett stycke trä från skogen hugger man ut dem, och konstnärens händer tillyxa dem;
med silver och guld pryder man dem och fäster dem med spikar och hammare, för att de icke skola falla omkull.
Lika fågelskrämmor på ett gurkfält stå de där och kunna ej tala; man måste bära dem, ty de kunna ej gå.
Frukten då icke för dem, ty de kunna ej göra något ont; och att göra något gott, det förmå de ej heller.
Men dig, HERRE, är ingen lik; du är stor, ditt namn är stort i makt.
Vem skulle icke frukta dig, du folkens konung?
Sådant tillkommer ju dig.
Ty bland folkens alla vise och i alla deras riken finnes ingen som är dig lik.
Nej, allasammans äro de oförnuftiga och dårar.
Avgudadyrkan är att dyrka trä,
silverplåt, hämtad från Tarsis, guld, fört ifrån Ufas, arbetat av en konstnär, av en guldsmeds händer.
I blått och rött purpurtyg stå de klädda, allasammans blott verk av konstförfarna män.
Men HERREN är en sann Gud, han är en levande Gud och en evig konung; för hans förtörnelse bävar jorden, och folken kunna icke uthärda hans vrede.
Så skolen I säga till dem: De gudar som icke hava gjort himmel och jord, de skola utrotas från jorden och ej få finnas under himmelen.
Han har gjort jorden genom sin kraft, han har berett jordens krets genom sin vishet, och genom sitt förstånd har han utspänt himmelen.
När han vill låta höra sin röst, då brusa himmelens vatten, då låter han regnskyar stiga upp från jordens ända; han låter ljungeldar komma med regn och för vinden ut ur dess förvaringsrum.
Såsom dårar stå då alla människor där och begripa intet; guldsmederna komma då alla på skam med sina beläten, ty deras gjutna beläten äro lögn, och ingen ande är i dem.
De äro fåfänglighet, en tillverkning att le åt; när hemsökelsen kommer över dem, måste de förgås.
Men sådan är icke han som är Jakobs del; nej, det är han som har skapat allt, och Israel är hans arvedels stam.
HERREN Sebaot är hans namn.
Samlen edert gods och fören det bort ur landet, I som sitten under belägring.
Ty så säger HERREN: Se, denna gång skall jag slunga bort landets inbyggare; jag skall bereda dem ångest, så att de förnimma det.
Ve mig, jag är sönderkrossad!
Oläkligt är mitt sår.
Men jag säger: Ja, detta är min plåga, jag måste bära den!
Mitt tält är förstört, och mina tältstreck äro alla avslitna.
Mina barn äro borta, de finnas icke mer; ingen är kvar, som kan slå upp mitt tält och sätta upp mina tältdukar.
Ty herdarna voro oförnuftiga, de frågade icke efter HERREN; därför hade de ingen framgång, och hela deras hjord blev förskingrad.
Lyssna, något höres!
Se, det nalkas!
Ett stort dån kommer från nordlandet för att göra Juda städer till en ödemark, till en boning för schakaler.
Jag vet det, HERRE: människans väg beror ej av henne, det står icke i vandrarens makt att rätt styra sina steg.
Så tukta mig, HERRE likväl med måtta; icke i din vrede, på det att du ej må göra mig till intet.
Utgjut din förtörnelse över hedningarna, som icke känna dig, och över de släkter som ej åkalla ditt namn. ty de hava uppätit Jakob, ja, uppätit och gjort ände på honom, och hans boning hava de förött.
Detta är det ord som kom till Jeremia från HERREN; han sade:
»Hören detta förbunds ord, och talen till Juda män och till Jerusalems invånare;
säg till dem: Så säger HERREN, Israels Gud: Förbannad vare den man som icke hör detta förbunds ord,
det som jag bjöd edra fader på den tid då jag förde dem ut ur Egyptens land, den smältugnen, i det jag sade: Hören min röst och gören detta, alldeles såsom jag bjuder eder, så skolen I vara mitt folk, och jag skall vara eder Gud,
på det att jag må hålla den ed som jag har svurit edra fäder: att giva dem ett land som flyter av mjölk och honung, såsom ock nu har skett.»
Och jag svarade och sade: »Ja, amen, HERRE.»
Och HERREN sade till mig: Predika allt detta i Juda städer och på gatorna i Jerusalem och säg: Hören detta förbunds ord och gören efter dem.
Ty både på den dag då jag förde edra fäder ut ur Egyptens land och sedan ända till denna dag har jag varnat dem, ja, titt och ofta har jag varnat dem och sagt: »Hören min röst»;
men de ville icke höra eller böja sitt öra därtill, utan vandrade var och en i sitt onda hjärtas hårdhet.
Därför lät jag ock komma över dem allt vad jag hade sagt i det förbund som jag bjöd dem hålla, men som de dock icke höllo.
Och HERREN sade till mig: Jag vet huru Juda män och Jerusalems invånare hava sammansvurit sig.
De hava vänt tillbaka till sina förfäders missgärningar, deras som icke ville höra mina ord.
Själva hava de så följt efter andra gudar och tjänat dem.
Ja, Israels hus och Juda hus hava brutit det förbund som jag slöt med deras fäder.
Därför säger HERREN så: Se, jag skall låta en olycka komma över dem, som de icke skola kunna undkomma; och när de då ropa till mig, skall jag icke höra dem.
Och om så Juda städer och Jerusalems invånare gå bort och ropa till de gudar åt vilka de pläga tända offereld, så skola dessa alls icke kunna frälsa dem i deras olyckas tid.
Ty så många som dina städer äro, så många hava dina gudar blivit, du Juda; och så många som gatorna äro i Jerusalem, så många altaren haven I satt upp åt skändlighetsguden: altaren till att tända offereld åt Baal.
Så må du nu icke bedja för detta folk eller frambära någon klagan och förbön för dem; ty jag vill icke höra, när de ropa till mig för sin olyckas skull.
Vad har min älskade att göra i mitt hus, då hon, ja, hela hopen, övar sådan skändlighet?
Kan heligt kött komma såsom offer från dig?
När du får bedriva din ondska, då fröjdar du dig ju.
»Ett grönskande olivträd, prytt med sköna frukter», så kallade HERREN dig; men nu har han med stort och väldigt dån tänt upp en eld omkring det trädet, så att dess grenar fördärvas.
Ja, HERREN Sebaot, han som planterade dig, har beslutit olycka över dig, för den ondskas skull som Israels och Juda hus hava bedrivit till att förtörna mig, i det att de hava tänt offereld åt Baal.
HERREN kungjorde det för mig, så att jag fick veta det; ja, du lät mig se vad de förehade.
Själv var jag såsom ett menlöst lamm som föres bort till att slaktas; jag visste ej att de förehade anslag mot mig: »Låt oss fördärva trädet med dess frukt, låt oss utrota honom ur de levandes land, så att man icke mer kommer ihåg hans namn.»
Men HERREN Sebaot är en rättfärdig domare, som prövar njurar och hjärta.
Så låt mig då få se din hämnd på dem, ty för dig har jag lagt fram min sak.
Därför säger HERREN så om Anatots män, dem som stå efter ditt liv och säga: »Profetera icke i HERRENS namn, om du icke vill dö för vår hand»
ja, därför säger HERREN Sebaot så: Se, jag skall hemsöka dem; deras unga män skola dö genom svärd, deras söner och döttrar skola dö genom hunger.
Och intet skall bliva kvar av dem; ty jag skall låta olycka drabba Anatots män, när deras hemsökelses år kommer.
HERRE, om jag vill gå till rätta med dig, så behåller du dock rätten.
Likväl måste jag tala med dig om vad rätt är.
Varför går det de ogudaktiga så väl?
Varför hava alla trolösa så god lycka?
Du planterar dem, och de slå rot; de växa och bära frukt.
Nära är du i deras mun, men fjärran är du från deras innersta.
Men du, HERRE, känner mig; du ser mig och prövar huru mitt hjärta är mot dig.
Ryck dem bort såsom får till att slaktas, och invig dem till en dödens dag.
Huru länge skall landet ligga sörjande och gräset på marken allestädes förtorka, så att både fyrfotadjur och fåglar förgås för inbyggarnas ondskas skull, under det att dessa säga: »Han skall icke se vår undergång»
Om du icke orkar löpa i kapp med fotgängare, huru vill du då taga upp tävlan med hästar?
Och om du nu känner dig trygg i ett fredligt land, huru skall det gå dig bland Jordanbygdens snår?
Se, till och med dina bröder och din faders hus äro ju trolösa mot dig; till och med dessa ropa med full hals bakom din rygg.
Du må icke tro på dem, om de ock tala vänligt till dig.
Jag har övergivit mitt hus, förskjutit min arvedel; det som var kärast för min själ lämnade jag i fiendehand.
Hon som är min arvedel blev mot mig såsom ett lejon i skogen; hon har höjt sin röst mot mig, därför har jag fattat hat till henne.
Skall min arvedel vara mot mig såsom en brokig rovfågel -- då må ock rovfåglar komma emot henne från alla sidor.
Upp, samlen tillhopa alla markens djur, och låten dem komma för att äta!
Herdar i mängd fördärva min vingård och förtrampa min åker; de göra min sköna åker till en öde öken.
Man gör den till en ödemark;
sörjande och öde ligger den framför mig.
Hela landet ödelägges, ty ingen finnes, som vill akta på.
Över alla höjder i öknen rycka förhärjare fram, ja, HERRENS svärd förtär allt, från den ena ändan av landet till den andra; intet kött kan finna räddning.
De hava sått vete, men skördat tistel; de hava mödat sig fåfängt.
Ja, I skolen komma på skam med eder gröda för HERRENS glödande vredes skull.
Så säger HERREN om alla de onda grannar som förgripa sig på den arvedel jag har givit åt mitt folk Israel: Se, jag skall rycka dem bort ur deras land, och Juda hus skall jag rycka undan ifrån dem.
Men därefter, sedan jag har ryckt dem bort, skall jag åter förbarma mig över dem och låta dem komma tillbaka, var och en till sin arvedel och var och en till sitt land.
Om de då rätt lära sig mitt folks vägar, så att de svärja vid mitt namn: »Så sant HERREN lever», likasom de förut lärde mitt folk att svärja vid Baal, då skola de bliva upprättade mitt ibland mitt folk.
Men om de icke vilja höra, så skall jag alldeles bortrycka och förgöra det folket, säger HERREN.
Så sade HERREN till mig: »Gå bort och köp dig en linnegördel, och sätt den omkring dina länder, men låt den icke komma i vatten.»
Och jag köpte en gördel, såsom HERREN hade befallt, och satte den omkring mina länder.
Då kom HERRENS ord till mig för andra gången; han sade:
»Tag gördeln som du har köpt, och som du bär omkring dina länder, och stå upp och gå bort till Frat, och göm den där i en stenklyfta.»
Och jag gick bort och gömde den vid Frat, såsom HERREN hade bjudit mig.
Sedan, en lång tid därefter, sade HERREN till mig: »Stå upp och gå bort till Frat, och hämta därifrån den gördel som jag bjöd dig gömma där.»
Och jag gick bort till Frat och grävde upp gördeln och hämtade fram den från det ställe där jag hade gömt den.
Och se, gördeln var fördärvad, så att den icke mer dugde till något.
Då kom HERRENS ord till mig; han sade:
Så säger HERREN: På samma sätt skall jag sända fördärv över Judas och Jerusalems stora högmod.
Detta onda folk, som icke vill höra mitt ord, utan vandrar i sitt hjärtas hårdhet och följer efter andra gudar och tjänar och tillbeder dem, det skall bliva såsom denna gördel vilken icke duger till något.
Ty likasom en mans gördel sluter sig tätt omkring hans länder, så lät jag hela Israels hus och hela Juda hus sluta sig till mig, säger HERREN, på det att de skulle vara mitt folk och bliva mig till berömmelse, lov och ära; men de ville icke höra.
Säg därför till dem detta ord: Så säger HERREN, Israels Gud: Alla vinkärl äro till för att fyllas med vin.
Och när de då säga till dig: »Skulle vi icke veta att alla vinkärl äro till för att fyllas med vin?»,
så svara dem: Så säger HERREN: Se, jag skall fylla detta lands alla inbyggare, konungarna som sitta på Davids tron, och prästerna och profeterna, ja, alla Jerusalems invånare, så att de bliva druckna.
Och jag skall krossa dem, den ene mot den andre, både fäder och barn, säger HERREN.
Jag skall icke hava någon misskund, icke skona och icke förbarma mig, så att jag avstår från att fördärva dem.
Hören och lyssnen härtill, varen icke övermodiga; ty HERREN har talat.
Given HERREN, eder Gud, ära, förrän han låter mörkret komma, och förrän edra fötter snubbla på bergen, när det skymmer; ty det ljus I förbiden skall han byta i dödsskugga och göra till töcken.
Men om I icke hören härpå, så måste min själ i lönndom sörja över sådant övermod, och mitt öga måste bitterligen gråta och flyta i tårar, därför att HERRENS hjord då bliver bortförd i fångenskap.
Säg till konungen och konungamodern: Sätten eder lågt ned, ty den härlighetens krona som prydde edert huvud har fallit av eder.
Städerna i Sydlandet äro tillslutna, och ingen finnes, som öppnar dem; hela Juda är bortfört i fångenskap, ja, bortfört helt och hållet.
Lyften upp edra ögon och sen huru de komma norrifrån.
Var är nu hjorden som var dig given, den hjord som var din ära?
Vad vill du säga, när han sätter till herrar över dig män som du själv har lärt att komma till dig såsom älskare?
Skulle du då icke gripas av vånda såsom en kvinna i barnsnöd?
Men om du säger i ditt hjärta: »Varför har det gått mig så?», så vet: for din stora missgärnings skull blev ditt mantelsläp upplyft och dina fötter nesligt blottade.
Kan väl en etiopier förvandla sin hud eller en panter sina fläckar?
Då skullen också I kunna göra något gott, I som ären så övade i ondska.
Välan, jag vill förskingra dem såsom strå som far bort för öknens vind.
Detta skall vara din lott och din beskärda del från mig, säger HERREN, därför att du har förgätit mig och förlitat dig på lögn.
Därför skall jag ock draga upp ditt mantelsläp över ditt ansikte, så att man får se din skam.
Din otukt, ditt vrenskande, ditt skändliga otuktsväsen -- på höjderna, på fältet har jag sett dina styggelser.
Ve dig, Jerusalem!
Du kommer icke att bliva ren -- på huru lång tid ännu?
Detta är det HERRENS ord som kom till Jeremia angående torkan.
Juda ligger sörjande, dess portar äro förfallna, likasom i sorgdräkt luta de mot jorden, och ett klagorop stiger upp från Jerusalem.
Stormännen där sända de små efter vatten, men när de komma till dammarna, finna de intet vatten; de måste vända tillbaka med tomma kärl.
De stå där med skam och blygd och måste hölja över sina huvuden.
För markens skull, som ligger vanmäktig, därför att intet regn faller på jorden, stå åkermännen med skam och måste hölja över sina huvuden.
Ja, också hinden på fältet övergiver sin nyfödda kalv, därför att intet grönt finnes
Och vildåsnorna stå på höjderna och flämta såsom schakaler; deras ögon försmäkta, därför att gräset är borta.
Om än våra missgärningar vittna emot oss, så hjälp dock, HERRE, för ditt namns skull.
Ty vår avfällighet är stor; mot dig hava vi syndat.
Du Israels hopp dess frälsare i nödens tid, varför är du såsom en främling i landet, lik en vägfarande som slår upp sitt tält allenast för en natt?
Varför är du lik en rådlös man, lik en hjälte som icke kan hjälpa?
Du bor ju dock mitt ibland oss, HERRE, och vi äro uppkallade efter ditt namn; så övergiv oss då icke.
Så säger HERREN om detta folk: På detta sätt driva de gärna omkring, de hålla icke sina fötter i styr.
Därför har HERREN intet behag till dem; nej, han kommer nu ihåg deras missgärning och hemsöker deras synder.
Och HERREN sade till mig: Du må icke bedja om något gott för detta folk.
Ty om de än fasta, så vill jag dock icke höra deras rop, och om de än offra brännoffer och spisoffer så har jag intet behag till dem, utan vill förgöra dem med svärd, hungersnöd och pest.
Då sade jag: »Ack Herre, HERRE!
Profeterna säga ju till dem: I skolen icke se något svärd, ej heller skall hungersnöd träffa eder, nej, en varaktig frid skall jag giva eder på denna plats.»
Men HERREN sade till mig: Profeterna profetera lögn i mitt namn; jag har icke sänt dem eller givit dem någon befallning eller talat till dem.
Lögnsyner och tomma spådomar och fåfängligt tal och sina egna hjärtans svek är det de profetera för eder.
Därför säger HERREN så om de profeter som profetera i mitt namn, fastän jag icke har sänt dem, och som säga att svärd och hungersnöd icke skola komma i detta land: Jo, genom svärd och hunger skola dessa profeter förgås.
Och folket som de profetera för, både män och hustrur, både söner och döttrar, skola komma att ligga på Jerusalems gator, slagna av hunger och svärd, och ingen skall begrava dem; och jag skall utgjuta deras ondska över dem.
Men du skall säga till dem detta ord: Mina ögon flyta i tårar natt och dag och få ingen ro, ty jungfrun, dottern mitt folk har drabbats av stor förstöring, av ett svårt och oläkligt sår.
Om jag går ut på marken, se, då ligga där svärdsslagna män; och kommer jag in i staden, så mötes jag där av hungerns plågor.
Ja, både profeter och präster nödgas draga från ort till ort, till ett land som de icke känna.
Har du då alldeles förkastat Juda?
Har din själ begynt försmå Sion?
Eller varför har du slagit oss så, att ingen kan hela oss?
Vi bida efter frid, men intet gott kommer, efter en tid då vi skulle bliva helade, men se, förskräckelse kommer.
HERRE, vi känna vår ogudaktighet, våra fäders missgärning, ty vi hava syndat mot dig.
För ditt namns skull, förkasta oss icke, låt din härlighets tron ej bliva föraktad; kom ihåg ditt förbund med oss, och bryt det icke.
Finnas väl bland hedningarnas fåfängliga avgudar sådana som kunna giva regn?
Eller kan himmelen av sig själv låta regnskurar falla?
Är det icke dig, HERRE, vår Gud, som vi måste förbida?
Det är ju du som har gjort allt detta.
Men HERREN sade till mig; Om än Mose och Samuel trädde inför mig, så skulle min själ dock icke vända sig till detta folk.
Driv dem bort ifrån mitt ansikte och låt dem gå.
Och om de fråga dig: »Vart skola vi gå?», så skall du svara dem: Så säger HERREN: I pestens våld den som hör pesten till, i svärdets våld den som hör svärdet till, i hungerns våld den som hör hungern till, i fångenskapens våld den som hör fångenskapen till.
Fyra slags hemsökelser skall jag låta komma över dem, säger HERREN: svärdet, som skall dräpa dem, hundarna, som skola släpa bort dem, himmelens fåglar och vilddjuren på marken, som skola äta upp och fördärva dem.
Och jag skall göra dem till en varnagel för alla riken på jorden, till straff för det som Manasse, Hiskias son, Juda konung, har gjort i Jerusalem.
Ty vem kan hava misskund med dig, Jerusalem, och vem kan ömka dig, och vem kan vilja komma för att fråga om det står väl till med dig?
Du själv försköt mig, säger HERREN; du gick din väg bort.
Därför uträckte jag mot dig min hand och fördärvade dig; jag hade tröttnat att förbarma mig.
Ja, jag kastade dem med kastskovel vid landets portar, jag gjorde föräldrarna barnlösa, jag förgjorde mitt folk, då de ej ville vända om från sina vägar.
Deras änkor blevo genom mig talrikare än sanden i havet; över mödrarna till deras unga lät jag förhärjare komma mitt på ljusa dagen; plötsligt lät jag ångest och förskräckelse falla över dem.
Om en moder än hade sju söner, måste hon dock giva upp andan i sorg; hennes sol gick ned, medan det ännu var dag, hon måste bliva till skam och blygd.
Och vad som är kvar av dem skall jag giva till pris åt deras fienders svärd, säger HERREN
»Ve mig, min moder, att du har fött mig, mig som är till kiv och träta för hela landet!
Jag har icke drivit ocker, ej heller har någon behövt ockra på mig; likväl förbanna de mig alla.»
Men HERREN svarade: »Sannerligen, jag skall styrka dig och låta det gå dig väl.
Sannerligen, jag skall så göra, att dina fiender komma och bönfalla inför dig i olyckans och nödens tid.
Kan man bryta sönder järn, järn från norden, eller koppar?» --
Ditt gods och dina skatter skall jag lämna till plundring, och det utan betalning, till straff för allt vad du har syndat i hela ditt land.
Och jag skall låta dina fiender föra dig in i ett land som du icke känner.
Ty min vredes eld är upptänd; mot eder skall det brinna.
HERRE, du vet det.
Tänk på mig och låt dig vårda om mig, och skaffa mig hämnd på mina förföljare; tag mig icke bort, du som är långmodig.
Betänk huru jag bär smälek för din skull
När jag fick dina ord, blevo de min spis, ja, dina ord blevo för mig mitt hjärtas fröjd och glädje; ty jag är uppkallad efter ditt namn, HERRE, härskarornas Gud.
Jag har icke suttit i gycklares samkväm och förlustat mig där; för din hands skull har jag måst sitta ensam, ty du har uppfyllt mig med förgrymmelse.
Varför skall jag då plågas så oavlåtligt, och varför är mitt sår så ohelbart?
Det vill ju icke läkas.
Ja, du bliver för mig såsom en försinande bäck, så som ett vatten som ingen kan lita på.
Därför säger HERREN så: Om du vänder åter, så vill jag låta dig komma åter och bliva min tjänare.
Och om du frambär ädel metall utan slagg, så skall du få tjäna mig såsom mun.
Dessa skola då vända åter till dig, men du skall icke vända åter till dem.
Och jag skall göra dig inför detta folk till en fast kopparmur, så att de icke skola bliva dig övermäktiga, om de vilja strida mot dig; ty jag är med dig och vill frälsa dig och vill hjälpa dig, säger HERREN.
Jag skall hjälpa dig ut ur de ondas våld och skall förlossa dig ur våldsverkarnas hand.
Och HERRENS ord kom till mig; han sade:
Du skall icke taga dig någon hustru eller skaffa dig några söner och döttrar på denna plats.
Ty så säger HERREN om de söner och döttrar som bliva I födda på denna plats, och om mödrarna som hava fött dem, och om fäderna som hava avlat dem i detta land:
Av svåra sjukdomar skola de dö; man skall icke hålla dödsklagan efter dem eller begrava dem, utan de skola bliva gödsel på marken.
Och genom svärd och hunger skola de förgås, och deras döda kroppar skola bliva mat åt himmelens fåglar och markens djur.
I
Ty så säger HERREN: Du skall icke gå in i något sorgehus och icke begiva dig åstad för att hålla dödsklagan, ej heller ömka dem; ty jag har tagit bort min frid ifrån detta folk, säger HERREN, ja, min nåd och barmhärtighet.
Och både stora och små skola dö i detta land, utan att bliva begravna; och man skall icke hålla dödsklagan efter dem, och ingen skall för deras skull rista märken på sig eller raka sitt huvud.
Man skall icke bryta bröd åt någon, för att trösta honom i sorgen efter en död, och icke giva någon tröstebägaren att dricka, när han har förlorat fader eller moder.
Och i gästabudshus skall du icke heller gå in för att sitta med dem och äta och dricka.
Ty så säger HERREN Sebaot, Israels Gud: Se, inför edra ögon, och medan I ännu leven, skall jag på denna plats göra slut på fröjderop och glädjerop, på rop för brudgum och rop för brud.
I
När du nu förkunnar alla dessa ord för detta folk och de då fråga dig: »Varför har HERREN uttalat över oss all denna stora olycka?
Och vari består den missgärning och synd som vi hava begått mot HERREN, vår Gud?»,
då skall du svara dem: »Jo, edra fäder övergåvo mig, säger HERREN, och följde efter andra gudar och tjänade och tillbådo dem; ja, mig övergåvo de och höllo icke min lag.
Och I själva haven gjort ännu mer ont, än edra fäder gjorde; ty se, I vandren var och en efter sitt onda hjärtas hårdhet, och I viljen icke höra mig.
Därför skall jag ock slunga eder bort ur detta land, till ett land son varken I eller edra fäder haven känt, och där Skolen I få tjäna andra gudar både dag och natt; ty jag skall icke hava någon misskund med eder.»
Se, därför skola dagar komma, säger HERREN, då man icke mer skall säga: »Så sant HERREN lever, han som har fört Israels barn upp ur Egyptens land»,
utan: »Så sant HERREN lever, han som har fört Israels barn upp ur nordlandet, och ur alla andra länder till vilka han hade drivit dem bort.»
Ty jag skall föra dem tillbaka till deras land, det som jag gav åt deras fäder.
Se, jag skall sända bud efter många fiskare, säger HERREN, och de skola fiska upp dem; och sedan skall jag sända bud efter många jägare, och de skola jaga dem ned från alla berg och alla höjder och ut ur stenklyftorna.
Ty mina ögon äro riktade på alla deras vägar; de kunna icke gömma sig för mitt ansikte och deras missgärning är icke fördold för mina ögon.
Och först skall jag i dubbelt mått vedergälla dem för deras missgärning och synd, för att de hava oskärat mitt land, i det att de hava uppfyllt min arvedel med sina styggeliga och skändliga avgudars döda kroppar.
HERRE, du min starkhet och mitt värn, du min tillflykt på nödens dag, till dig skola hedningarna komma från jordens ändar och skola säga: »Allenast lögn hava våra fäder fått i arv. fåfängliga avgudar, av vilka ingen kan hjälpa.
Kan väl en människa göra sig gudar?
Nej, de gudarna äro inga gudar.
Därför vill jag nu denna gång låta dem förnimma det, jag vill låta dem känna min hand och min makt, för att de må veta att mitt namn är HERREN.
Juda synd är uppskriven med järnstift, med diamantgriffel; den är inristad på deras hjärtas tavla och på edra altarens horn,
så visst som deras barn vid gröna träd och på höga kullar komma ihåg sina altaren och Aseror.
Du mitt berg på fältet, ditt gods, ja, alla dina skatter skall jag lämna till plundring, så ock dina offerhöjder, till straff för vad du har syndat i hela ditt land.
Och du skall nödgas avstå -- och detta genom din egen förskyllan -- från den arvedel som jag har givit dig; och jag skall låta dig tjäna dina fiender i ett land som du icke känner.
Ty I haven upptänt min vredes eld, och den skall brinna till evig tid.
Så säger HERREN: Förbannad är den man som förtröstar på människor och sätter kött sig till arm och med sitt hjärta viker av ifrån HERREN.
Han skall bliva såsom en torr buske på hedmarken och skall icke få se något gott komma, utan skall bo på förbrända platser i öknen, i ett land med salthedar, där ingen bor.
Men välsignad är den man som förtröstar på HERREN, den som har HERREN till sin förtröstan.
Han är lik ett träd som är planterat vid vatten, och som sträcker ut sina rötter till bäcken; ty om än hetta kommer, så förskräckes det icke, utan bevarar sina löv grönskande; och om ett torrt år kommer, så sörjer det icke och upphör ej heller att bara frukt.
Ett illfundigt och fördärvat ting är hjärtat framför allt annat; vem kan förstå det?
Dock, Jag, HERREN, utrannsakar hjärtat och prövar njurarna, och giver så åt var och en efter hans vägar, efter hans gärningars frukt.
Lik en rapphöna som ruvar på ägg, vilka hon ej själv har lagt, är den som samlar rikedom med orätt; i sina halva dagar måste han lämna den och vid sitt slut skall han stå såsom en dåre.
En härlighetens tron, en urgammal höjd är vår helgedoms plats.
HERREN är Israels hopp; alla som övergiva dig komma på skam. de som vika av ifrån mig likna en skrift i sanden; ty de hava övergivit HERREN, källan med det friska vattnet.
Hela du mig, HERRE, så varde jag helad; fräls mig du, så varder jag frälst.
Ty du är mitt lov.
Se, dessa säga till mig: »Vad bliver av HERRENS ord?
Må det fullbordas!»
Det är ju så, att jag ej har undandragit mig herdekallet i din efterföljd, och fördärvets dag har jag icke åstundat; du vet det själv.
Vad mina läppar hava uttalat, det har talats inför ditt ansikte.
Så bliv då icke till skräck för mig; du som är min tillflykt på olyckans dag.
Låt dem som förfölja mig komma på skam, men låt icke mig komma på skam; låt dem bliva förfärade, men låt ej mig bliva förfärad.
Låt en olycksdag komma över dem, och krossa dem i dubbelt mått.
Så sade HERREN till mig: Gå åstad och ställ dig i Menighetsporten, där Juda konungar gå in och gå ut, och sedan i Jerusalems alla andra portar;
och säg till dem: Hören HERRENS ord, I Juda konungar med hela Juda, och I alla Jerusalems invånare som gån in genom dessa portar.
Så säger HERREN: Tagen eder val till vara för att på sabbatsdagen bära någon börda eller föra in någon sådan genom Jerusalems portar.
Och fören icke på sabbatsdagen någon börda ut ur edra hus, och gören ej heller något annat arbete, utan helgen sabbatsdagen, såsom jag bjöd edra fäder,
fastän de icke ville höra eller böja sitt öra därtill, utan voro hårdnackade, så att de icke hörde eller togo emot tuktan.
Men om I viljen höra mig, säger HERREN, så att I på sabbatsdagen icke fören någon börda in genom denna stads portar, utan helgen sabbatsdagen, så att I på den icke gören något arbete,
då skola konungar och furstar som komma att sitta på Davids tron få draga in genom denna stads portar, på vagnar och hästar, följda av sina furstar, av Juda man och Jerusalems invånare; och denna stad skall då förbliva bebodd evinnerligen.
Och från Juda städer, från Jerusalems omnejd och från Benjamins land, från Låglandet, Bergsbygden och Sydlandet skall man komma och frambära brännoffer, slaktoffer, spisoffer och rökelse och frambära lovoffer till HERRENS hus.
Men om I icke hören mitt bud att helga sabbaten och att icke bära någon börda in genom Jerusalems portar på sabbatsdagen, då skall jag tända eld på dess portar, och elden skall förtära Jerusalems palatser och skall icke kunna utsläckas.
Detta är det ord som kom till Jeremia från HERREN; han sade
»Stå upp och gå ned till krukmakarens hus; där vill jag låta dig höra mina ord.»
Då gick jag ned till krukmakarens hus och fann honom upptagen med arbete på krukmakarskivan.
Och när kärlet som krukmakare höll på att göra av leret misslyckades i hans hand, begynte han omigen, och gjorde därav ett annat kärl så, som han ville hava det gjort.
Och HERRENS ord kom till mig han sade:
Skulle jag icke kunna göra med eder, I är Israels hus, såsom denne krukmakare gör? säger HERREN Jo, såsom leret är i krukmakarens hand, så ären ock I i min hand, I av Israels hus.
Den ena gången hotar jag ett folk och ett rike att jag vill upprycka, nedbryta och förgöra det;
men om då det folket omvänder sig från det onda väsende mot vilket jag vände mitt hot, så ångrar jag det onda som jag hade tänkt att göra dem.
En annan gång lovar jag ett folk och ett rike att jag vill uppbygga och plantera det;
men om det då gör vad ont är i mina ögon och icke hör min röst, så ångrar jag det goda som jag hade sagt att jag ville göra dem.
Så säg du nu till Juda man och Jerusalems invånare: Så säger HERREN: Se, jag bereder åt eder en olycka, och jag har i sinnet ett anslag mot eder.
Vänden därför om, var och en från sin onda väg, och bättren edert leverne och edert väsende.
Men de skola svara: »Du mödar dig förgäves.
Vi vilja följa vara egna tankar och göra var och er efter sitt onda hjärtas hårdhet.
Därför säger HERREN så: Frågen efter bland hednafolken om någon har hört något sådant.
Alltför gruvliga ting har jungfrun Israel bedrivit.
Övergiver då Libanons snö sin upphöjda klippa, eller sina de friska vatten ut, som strömma ifrån fjärran,
eftersom mitt folk förgäter mig och tänder offereld åt avgudar?
Se, av dem skola de bringas på fall, när de gå sin gamla stråt och vandra på villostigar, på obanade vägar.
Så göra de sitt land till ett föremål för häpnad, för begabberi evinnerligen; alla som gå där fram skola häpna och skaka huvudet.
Såsom en östanvind skall jag förskingra dem, när fienden kommer; jag skall visa dem ryggen och icke ansiktet, på deras ofärds dag.
Men de sade: »Kom, låt oss tänka ut något anslag mot Jeremia.
Ty prästerna skola icke komma till korta med undervisning, ej heller de vise med råd, ej heller profeterna med förkunnelse.
Ja, kom, låt oss fälla honom med vara tungor, vi behöva alls icke akta på vad han säger.»
HERRE, akta du på mig, och hör rad mina motståndare tala.
Skall man få vedergälla gott med ont, eftersom dessa hava grävt en grop för mitt liv?
Tänk på huru jag har stått inför ditt ansikte för att mana gott för dem, till att avvända från dem din vrede.
Därför må du överlämna deras barn åt hungersnöden och giva dem själva till pris åt svärdet, så att deras hustrur bliva barnlösa och änkor, deras män dräpta av pesten, och deras ynglingar slagna med svärd striden.
Må klagorop höras från deras hus, i det att du plötsligt låter rövarskaror komma över dem.
Ty de hava grävt en grop för att fånga mig, och snaror hava de lagt ut för mina fötter.
Men du, HERRE, känner alla deras mordiska anslag mot mig; så må du då icke förlåta dem deras missgärning eller utplåna deras synd ur din åsyn.
Må de bringas på fall inför dig; ja, utför ditt verk mot dem på din vredes tid.
Så sade HERREN: Gå åstad och köp dig en lerkruka av krukmakaren; och tag med dig några av de äldste i folket och av de äldste bland prästerna,
och gå ut till Hinnoms sons dal, som ligger framför Lerskärvsporten, och predika där de ord som jag skall tala till dig.
Du skall säga: »Hören HERRENS ord, I Juda konungar och I Jerusalems invånare: Så säger HERREN Sebaot, Israels Gud: Se, jag skall låta en sådan olycka komma över denna plats, att det skall genljuda i öronen på var och en som får höra det.
Eftersom de hava övergivit mig och icke aktat denna plats, utan där tänt offereld åt andra gudar, som varken de själva eller deras fäder eller Juda konungar hava känt, och eftersom de hava uppfyllt denna plats med oskyldigas blod,
och byggt sina Baalshöjder, för att där bränna upp sina barn i eld, till brännoffer åt Baal, fastän jag aldrig har bjudit eller talat om eller ens tänkt mig något sådant,
se, därför skola dagar komma, säger HERREN, då man icke mer skall kalla denna plats 'Tofet' eller 'Hinnoms sons dal', utan 'Dråpdalen'.
Och då skall jag på denna plats göra om intet Judas och Jerusalems råd, och jag skall låta dem falla för deras fienders svärd och för de mäns hand, som stå efter deras liv och jag skall giva deras döda kroppar till mat åt himmelens fåglar och markens djur.
Och jag skall göra denna stad till ett föremål för häpnad och begabberi; alla som gå där från skola häpna och vissla vid tanken på alla dess plågor.
Och jag skall låta dem äta sina egna söners och döttrars kött, ja, den ene skall nödgas äta den andres kött.
I sådan nöd och sådant trångmål skola de komma genom sina fiender och genom dem som stå efter deras liv.»
Och du skall slå sönder krukan inför de mäns ögon, som hava gått med dig,
och du skall säga till dem: »Så säger HERREN Sebaot: Jag skall sönderslå detta folk och denna stad, på samma sätt som man slår sönder ett krukmakarkärl, så att det icke kan bliva helt igen; och man skall begrava i Tofet, därför att ingen annan plats finnes att begrava på.
Så skall jag göra med denna plats, säger HERREN, och med dess invånare; jag skall göra denna stad lik Tofet.
Och husen i Jerusalem och Juda konungars hus, de orena, skola bliva såsom Tofetplatsen, ja, alla de hus på vilkas tak man har tänt offereld åt himmelens hela härskara och utgjutit drickoffer åt andra gudar.»
När sedan Jeremia kom igen från Tofet, dit HERREN hade sänt honom för att profetera, ställde han sig i förgården till HERRENS hus och sade till allt folket:
»Så säger HERREN Sebaot, Israels Gud: Se, över denna stad med alla dess lydstäder skall jag låta all den olycka komma, som jag har beslutit över den -- detta därför att de hava varit hårdnackade och icke velat höra mina ord.»
Då nu Pashur, Immers son, prästen, som var överuppsyningsman i HERRENS hus, hörde Jeremia profetera detta,
lät han hudflänga profeten Jeremia och satte honom i stocken i Övre Benjaminsporten till HERRENS hus.
Men när Pashur dagen därefter släppte Jeremia lös ur stocken, sade Jeremia till honom: »Pashur är icke det namn varmed HERREN benämner dig, utan Magor-Missabib;
ty så säger HERREN: Se, jag skall göra dig till skräck såväl för dig själv som för alla dina vänner; och de skola falla för sina fienders svärd, i din egen åsyn.
Och hela Juda skall jag giva i den babyloniske konungens hand, och han skall föra dem bort till Babel och dräpa dem med svärd.
Och jag skall giva denna stads alla rikedomar, allt dess gods och alla dyrbarheter däri, ja, Juda konungars alla skatter skall jag giva i deras fienders hand; och de skola göra det till sitt byte och taga det och föra det till Babel.
Och du själv, Pashur, skall gå i fångenskap, med alla som bo i ditt hus.
Du skall komma till Babel; där skall du dö, och där skall du begravas, Sjungen till HERRENS ära, jämte alla dina vänner, för vilka du har profeterat lögn.»
Du, HERRE, övertalade mig, och jag lät mig övertalas; du grep mig och blev mig övermäktig.
Så har jag blivit ett ständigt åtlöje; var man bespottar mig.
Ty' så ofta jag talar, måste jag klaga; jag måste ropa över våld och förtryck, ty HERRENS ord har blivit mig till smälek och hån beständigt.
Men när jag sade: »Jag vill icke tänka på honom eller vidare tala i hans namn», då blev det i mitt hjärta såsom brunne där en eld, instängd i mitt innersta; jag mödade mig med att uthärda den, men jag kunde det icke.
Ty jag hör mig förtalas av många; skräck från alla sidor! »Anklagen honom!» »Ja, vi vilja anklaga honom!»
Alla som hava varit mina vänner vakta på att jag skall falla: »Kanhända skall han låta locka sig, så att vi bliva honom övermäktiga och få taga hämnd på honom.»
Men HERREN är med mig såsom en väldig hjälte; därför skola mina förföljare komma på fall och intet förmå.
Ja, de skola storligen komma på skam, därför att de ej hade förstånd; de skola drabbas av en evig blygd, som icke skall varda förgäten
Ty HERREN Sebaot prövar med rättfärdighet, han ser njurar och hjärta.
Så skall jag då få se din hämnd på dem, ty för dig har jag lagt fram min sak.
Sjungen till HERRENS ära, loven HERREN; ty han räddar den fattiges själv ur de ondas hand.
Förbannad vare den dag på vilken jag föddes; utan välsignelse blive den dag då min moder födde mig.
Förbannad vare den man som förkunnade för min fader: »Ett gossebarn är dig fött», och så gjorde honom stor glädje.
Gånge det den mannen såsom det gick de städer som HERREN omstörtade utan förbarmande.
Må han få höra klagorop om morgonen och härskri om middagen.
därför att han icke dräpte mig strax i moderlivet, så att min moder fick bliva min grav och hennes liv vara havande för evigt.
Varför kom jag ut ur moderlivet och fick se olycka och bedrövelse, så att mina dagar måste försvinna i skam?
Detta är det ord som kom till Jeremia från HERREN, när konung Sidkia sände till honom Pashur, Malkias son, och prästen Sefanja, Maasejas son, och lät säga:
»Fråga HERREN för oss, då nu Nebukadressar, konungen i Babel, har angripit oss; kanhända vill HERREN handla med oss i enlighet med alla sina förra under, så att denne lämnar oss i fred.
Jeremia svarade dem: Så skolen I säga till Sidkia:
Så säger HERREN, Israels Gud Se, de vapen i eder hand, med vilka I utanför muren striden mot konungen i Babel och kaldéerna, som belägra eder, dem skall jag vända om och skall famla dem inne i denna stad.
Och jag skall själv strida mot eder med uträckt hand och stark arm, vrede och harm och stor förtörnelse.
Och jag skall slå dem som bo i denna stad, både människor och djur; i svår pest skola de dö.
Och därefter, säger HERREN, skall jag låta Sidkia, Juda konung, och hans tjänare och folket, dem som i denna stad äro kvar efter pesten svärdet och hungersnöden, falla i Nebukadressars, den babyloniske konungens, hand och i deras fienders hand, i de mäns hand, som stå efter deras liv.
Och han skall slå dem med svärdsegg; han skall icke skona dem och icke hava någon misskund eller något förbarmande.
Och till detta folk skall du säga Så säger HERREN: Se, jag förelägger eder vägen till livet och vägen till döden.
Den som stannar kvar i denna stad, han skall dö genom svärd eller hunger eller pest, men den som går ut och giver sig åt kaldéerna, som belägra eder, han skall få leva och vinna sitt liv såsom ett byte.
Ty jag har vänt mitt ansikte mot denna stad, till dess olycka och icke till dess lycka, säger HERREN.
Den skall bliva given i den babyloniske konungens hand, och han skall bränna upp den i eld.
Och till Juda konungs hus skall du säga: Hören HERRENS ord:
I av Davids hus, så säger HERREN: »Fällen var morgon rätt dom, och rädden den plundrade ur förtryckarens hand, för att icke min vrede må bryta fram såsom en eld och brinna så, att ingen kan utsläcka den» -- detta för deras onda väsendes skull.
Se, jag skall vända mig mot dig, du som bor i dalen, du bergfäste på slätten, säger HERREN, ja, mot eder som sägen: »Vem kan falla över oss, och vem kan tränga in i våra boningar?»
Jag skall hemsöka eder efter edra gärningars frukt, säger HERREN.
Ja, jag skall tända upp en eld i deras skog, och den skall förtära allt där runt omkring.
Så sade HERREN: Gå ned till Juda konungs hus och tala där följande ord;
säg: Hör HERRENS ord, du Juda konung, som sitter på Davids tron, hör det du med dina tjänare och ditt folk, I som gån in genom dessa portar.
Så säger HERREN: Öven rätt och rättfärdighet, och rädden den plundrade ur förtryckarens hand; förorätten icke främlingen, den faderlöse och änkan, gören icke övervåld mot dem, och utgjuten icke oskyldigt blod på denna plats.
Ty om I gören efter detta ord, så skola konungar som komma att sitta på Davids tron få draga in genom portarna till detta hus, på vagnar och hästar, följda av sina tjänare och sitt folk.
Men om I icke hören dessa ord, då har jag svurit vid mig själv, säger HERREN, att detta hus skall bliva ödelagt.
Ty så säger HERREN om Juda konungs hus: Väl är du för mig såsom ett Gilead, såsom Libanons topp; men jag skall sannerligen göra dig till en öken, till obebodda städer.
Och jag skall inviga fördärvare till att komma över dig, var och en med sina vapen, och de skola hugga ned dina väldiga cedrar och kasta dem i elden
Och många folk skola gå fram vid denna stad, och man skall fråga varandra: »Varför har HERREN gjort så mot denna stora stad?»
Och man skall då svara Därför att de övergåvo HERREN sin Guds, förbund och tillbådo andra gudar och tjänade dem.»
Gråten icke över en död man, och ömken honom icke; men gråten bitterligen över honom som har måst vandra bort, ty han skall icke mer komma tillbaka och återse sitt fädernesland.
Ty så säger HERREN om Sallum, Josias son, Juda konung, som blev konung efter sin fader Josia, och som har dragit bort ifrån denna plats: Han skall icke mer komma hit tillbaka,
utan på den ort dit han har blivit bortförd i fångenskap, där skall han dö; detta land skall han icke mer få återse.
Ve dig, du som bygger ditt hus med orättfärdighet och dina salar med orätt, du som låter din nästa arbeta för intet och icke giver honom hans lön,
du som säger: »Jag vill bygga mig ett stort hus med rymliga salar», och så gör åt dig vida fönster och belägger huset med cederträ och målar det rött med dyrbar färg!
Kallar du det att vara konung, att du ävlas med att bygga cederhus?
Din fader åt ju och drack, dock övade han rätt och rättfärdighet; och då gick det honom väl.
Han skaffade den betryckte och fattige rätt; och då gick det väl.
Är icke detta att känna mig? säger HERREN.
Men dina ögon och ditt hjärta stå allenast efter vinning och efter att utgjuta den oskyldiges blod och att öva förtryck och våld.
Därför säger HERREN så om Jojakim, Josias son, Juda konung: Man skall ej hålla dödsklagan efter honom och ropa: »Ack ve, min broder!
Ack ve, syster!»
Man skall ej hålla dödsklagan efter honom och ropa: »Ack ve, herre!
Ack ve, huru härlig han var!»
Såsom man begraver en åsna, så skall han begravas; han skall släpas ut och kastas bort, långt utanför Jerusalems portar.
Stig upp på Libanon och ropa, häv upp din röst i Basan, och ropa från Abarim, ty alla dina älskare äro krossade.
Jag talade till dig, när det gick dig väl, men du sade: »Jag vill icke höra.»
Sådan har din väg varit allt ifrån din ungdom, att du icke har velat höra min röst.
Alla dina herdar skola nu få en stormvind till sin herde, och dina älskare måste gå i fångenskap.
Ja, då skall du komma på skam och få blygas för all din ondskas skull.
Du som bor på Libanon, du som har ditt näste i cedrarna, huru skall du icke jämra dig, när vånda kommer över dig, ångest lik en barnaföderskas!
Så sant jag lever, säger HERREN, om du, Konja, Jojakims son, Juda konung, än vore en signetring på min högra hand, så skulle jag dock rycka dig därifrån.
Och jag skall giva dig i de mäns hand, som stå efter ditt liv, och i de mäns hans som du fruktar för, nämligen i Nebukadressars, den babyloniske konungens, hand och i kaldéernas hand.
Och dig och din moder, den som har fött dig, skall jag slunga bort till ett annat land, där I icke ären födda; och där skolen I dö.
Till det land dit deras själ längtar att återvända, dit skola de icke få vända åter.
Är då han, denne Konja, ett föraktligt, krossat beläte eller ett värdelöst kärl?
Eller varför hava de blivit bortslungade, han och hans avkomlingar, och kastade bort till ett land som de icke hava känt?
O land, land, land, hör HERRENS ord!
Så säger HERREN: Tecknen upp denne man såsom barnlös, såsom en man som ingen lycka har haft i sina livsdagar.
Ty ingen av hans avkomlingar skall vara så lyckosam att han får sitta på Davids tron och i framtiden råda över Juda.
Ve över de herdar som fördärva och förskingra fåren i min hjord! säger HERREN.
Därför säger HERREN, Israels Gud, så om de herdar som föra mitt folk i bet: Det är I som haven förskingrat mina får och drivit bort dem och underlåtit att söka deras bästa.
Men se, nu skall jag hemsöka eder för edert onda väsendes skull, säger HERREN.
Och jag skall själv församla kvarlevan av mina får ur alla de länder till vilka jag har drivit dem bort, och skall föra dem tillbaka till deras betesmarker, och de skola bliva fruktsamma och föröka sig.
Och jag skall låta herdar uppstå åt dem, vilka skola föra dem i bet; och de skola icke mer behöva frukta eller förskräckas och skola icke mer drabbas av hemsökelse, säger HERREN.
Se, dagar skola komma, säger HERREN, då jag skall låta en rättfärdig telning uppstå åt David.
Han skall regera såsom konung och hava framgång, och han skall skaffa rätt och rättfärdighet på jorden.
I hans dagar skall Juda varda frälst och Israel bo i trygghet; och detta skall vara det namn han skall få: HERREN vår rättfärdighet.
Se, därför skola dagar komma, säger HERREN, då man icke mer skall säga: »Så sant HERREN lever, han som har fört Israels barn upp ur Egyptens land»,
utan: »Så sant HERREN lever, han som har fört upp Israels hus släkt och hämtat dem ut ur nordlandet och ur alla andra länder till vilka jag hade drivit dem bort.»
Och så skola de få bo i sitt land.
Om profeterna.
Mitt hjärta vill brista i mitt bröst, alla ben i min kropp äro vanmäktiga.
Jag är såsom en drucken man, en man överväldigad av vin, inför HERREN och inför hans heliga ord.
Ty landet är fullt av äktenskapsbrytare, under förbannelse ligger landet sörjande, och betesmarkerna i öknen äro förtorkade; man hastar till vad ont är och har sin styrka i orättrådighet.
Ty både profeter och präster äro gudlösa; ända inne i mitt hus har jag mött deras ondska, säger HERREN.
Därför skall deras väg bliva för dem såsom en slipprig stig i mörkret, de skola på den stöta emot och falla.
Ty jag vill låta olycka drabba dem, när deras hemsökelses är kommer, säger HERREN.
Väl såg jag ock hos Samarias profeter vad förvänt var; de profeterade i Baals namn och förde mitt folk Israel vilse.
Men hos Jerusalems profeter har jag sett de gruvligaste ting: de leva i äktenskapsbrott och fara med lögn; de styrka modet hos dem som göra ont, så att ingen vill omvända sig från sin ondska.
De äro alla för mig såsom Sodom, och stadens invånare såsom Gomorras.
Därför säger HERREN Sebaot så om profeterna: Se, jag skall giva dem malört att äta och gift att dricka, ty från profeterna i Jerusalem har gudlöshet gått ut över hela landet.
Så säger HERREN Sebaot: Hören icke på de profeters ord, som profetera för eder, ty de bedraga eder; sina egna hjärtans syner tala de, icke vad som kommer från HERRENS mun.
De säga alltjämt till dem som förakta mig: »HERREN har så talat: Det skall gå eder väl.»
Och till var och en som vandrar i sitt hjärtas hårdhet säga de: »Ingen olycka skall komna över eder.»
Vilken av dem har då fått tillträde till HERRENS råd, så att han kan förnimma och höra hans ord?
Och vilken har aktat på hans ord och lyssnat därtill?
Se, en stormvind från HERREN är här, hans förtörnelse bryter fram, en virvlande storm!
Över de ogudaktigas huvuden virvlar den ned.
Och HERRENS vrede skall icke upphöra, förrän han har utfört och fullbordat sitt hjärtas tankar; i kommande dagar skolen I förvisso förnimma det.
Jag sände icke dessa profeter, utan själva lupo de åstad; jag talade icke till dem, utan själva profeterade de.
Om de verkligen hade tillträde till mitt råd, så borde de förkunna mina ord för mitt folk och förmå dem att vända om från sin onda väg och sitt onda väsende.
Ar jag väl en Gud allenast på nära håll, säger HERREN, och icke en Gud också i fjärran?
Eller skulle någon kunna gömma sig på ett så lönnligt ställe att jag icke skulle se honom? säger HERREN.
Är jag icke den som uppfyller himmel och jord? säger HERREN.
Jag har hört vad profeterna säga, de som profetera lögn i mitt namn; de säga: »Jag har haft en dröm, jag har haft en dröm.»
Huru länge skall detta vara?
Hava de något i sinnet, dessa profeter som profetera lögn, och som äro profeter genom sina egna hjärtans svek,
dessa som tänka att de genom sina drömmar; dem som de förtälja för varandra, skola komma mitt folk att förgäta mitt namn, likasom deras fäder glömde mitt namn för Baal?
Den profet som har haft en dröm, han må förtälja sin dröm; men den som bar undfått mitt ord, han må tala mitt ord i sanning.
Vad har halmen att skaffa med säden? säger HERREN.
Är icke mitt ord såsom en eld, säger HERREN, och likt en hammare som krossar sönder klippor?
Se, därför skall jag komma över profeterna, säger HERREN, dessa som stjäla mina ord, den ene från den andre;
ja, jag skall komma över profeterna, säger HERREN, dessa som frambära sin egen tungas ord, men säga: »Så säger HERREN.»
Ja, jag skall komma över dem som profetera lögndrömmar, säger HERREN, och som, när de förtälja dem, föra mitt folk vilse med sina lögner och sin stortalighet, fastän jag icke har sänt dem eller givit dem något uppdrag, och fastän de alls icke kunna hjälpa detta folk, säger HERREN.
Om nu detta folk eller en profet eller en präst gör dig denna fråga: »Vad förkunnar HERRENS tunga?», så skall du säga till dem vad som är den verkliga »tungan», och att jag därför skall kasta eder bort, säger HERREN.
Och den profet eller den präst eller den av folket, som säger »HERRENS tunga», den mannen och hans hus skall jag hemsöka.
Nej, så skolen I fråga varandra och säga eder emellan: »Vad har HERREN svarat?», eller: »Vad har HERREN talat?»
Men Om HERRENS »tunga» mån I icke mer orda; ty en tunga skall då vars och ens eget ord bliva för honom, eftersom I förvänden den levande Gudens, HERRENS Sebaots, vår Guds, ord.
Så skall du säga till profeten: »Vad har HERREN svarat dig?», eller: vad har HERREN talat?»
Men om I sägen »HERRENS tunga», då säger HERREN så: »Eftersom I sägen detta ord 'HERRENS tunga', fastän jag har sänt bud till eder och låtit säga: I skolen icke säga 'HERRENS tunga',
därför skall jag nu alldeles förgäta eder och kasta eder bort ifrån mitt ansikte, med den stad som jag har givit åt eder och edra fäder.
Och jag skall låta en evig smälek komma över eder, och en evig blygd, som icke skall varda förgäten.»
HERREN lät mig se följande syn: Jag fick se två korgar med fikon uppställda framför HERRENS tempel; och det var efter det att Nebukadressar, konungen i Babel, hade fört bort ifrån Jerusalem Jekonja, Jojakims son, konungen i Juda, så ock Juda furstar, jämt timmermännen och smederna, och låtit dem komma till Babel.
I den ena korgen funnos mycket goda fikon, sådana som fikon ifrån förstlingsskörden äro; och i de andra korgen funnos mycket usla fikon, så usla att de icke kunde ätas.
Och HERREN sade till mig: »Vad ser du, Jeremia?»
Jag svarade »Fikon; och de goda fikonen är mycket goda, men de usla fikonen äro mycket usla, så usla att de icke kunna ätas.»
Och HERRENS ord kom till mig han sade:
Så säger HERREN, Israels Gud: Såsom man med välbehag ser på de goda fikonen, så vill jag med välbehag se till de bortförda av Juda, dem som jag från denna plats har sänt bort till kaldéernas land.
Jag skall med välbehag vända mitt öga till dem och låta dem komma tillbaka till detta land.
Jag skall uppbygga dem och icke slå ned dem; jag skall plantera dem och icke upprycka dem.
Och jag skall giva dem hjärtan till att känna att jag är HERREN; och de skola vara mitt folk, och jag skall vara deras Gud.
Ty de skola omvända sig till mig av allt sitt hjärta.
Men såsom man gör med usla fikon, som äro så usla att de icke kunna ätas, likaså, säger HERREN, skall jag göra med Sidkia, Juda konung, och med hans furstar och med kvarlevan i Jerusalem, ja, både med dem som hava blivit kvar här i landet och med dem som hava bosatt sig i Egyptens land.
På alla orter dit jag fördriver dem skall jag göra dem till en varnagel och en skräckbild för alla riken jorden, till en smälek, till ett ordspråk och en visa, och till ett exempel som man nämner, när man förbannar.
Och jag skall sända bland dem svärd, hungersnöd och pest, till dess att de bliva utrotade ur det land som jag har givit åt dem och deras fäder.
Detta är det ord som kom till Jeremia angående hela Juda folk, i Jojakims, Josias sons, Juda konungs, fjärde regeringsår, vilket var Nebukadressars, den babyloniske konungens, första regeringsår.
Och detta ord talade profeten Jeremia till hela Juda folk och till alla Jerusalems invånare; han sade:
Allt ifrån Josias, Amons sons, Juda konungs, trettonde regeringsår ända till denna dag, eller nu under tjugutre år, har HERRENS ord kommit till mig; men fastän jag titt och ofta har talat till eder, haven I icke velat höra.
Och fastän HERREN titt och ofta har sänt till eder alla sina tjänare profeterna, haven I icke velat höra.
I böjden icke edra öron till att höra,
när de sade: »Vänden om, var och en från sin onda väg och sitt onda väsende, så skolen I för evärdliga tider få bo kvar i det land som HERREN har givit åt eder och edra fäder.
Och följen icke efter andra gudar, så att I tjänen och tillbedjen dem; och förtörnen mig icke genom edra händers verk, på det att jag icke må låta olycka komma över eder.
I villen icke höra på mig, säger HERREN, och så förtörnaden I mig genom edra händers verk, eder själva till olycka.
Därför säger HERREN Sebaot så: Eftersom I icke villen höra mina ord,
därför skall jag sända åstad och hämta alla nordens folkstammar, säger HERREN, och skall sända bud till min tjänare Nebukadressar, konungen i Babel; och jag skall låta dem komma över detta land och dess inbyggare, så ock över alla folken här runt omkring.
Och dem skall jag giva till spillo, och skall göra dem till ett föremål för häpnad och begabberi, och låta deras land bliva ödemarker för evärdlig tid.
Och jag skall i dem göra slut på fröjderop och glädjerop, på rop för brudgum och rop för brud, på buller av kvarn och ljus från lampa.
Ja, hela detta land skall bliva ödelagt och förött, och dessa folk skola vara Babels konung underdåniga i sjuttio år.
Men när sjuttio år äro till ända skall jag hemsöka konungen i Babel och folket där för deras missgärning, säger HERREN, och hemsöka kaldéernas land och göra det till en ödemark för evärdlig tid.
Och jag skall på det landet låta alla de ord fullbordas, som jag har talat mot det, allt vad som är skrivet i denna bok, och vad Jeremia har profeterat mot alla dessa folk.
Ty också dem skola mäktiga folk och stora konungar göra sig underdåniga, och jag skall vedergälla dem efter deras gärningar och deras händers verk.
Ty så sade HERREN, Israels Gud, till mig: »Tag denna kalk med vredesvin ur min hand, och giv alla de folk till vilka jag sänder dig att dricka därur.
Må de dricka, så att de ragla och mista sansen, när det svärd kommer, som jag skall sända ibland dem.»
Och jag tog kalken ur HERRENS hand och gav alla de folk att dricka, till vilka HERREN sände mig,
nämligen Jerusalem med Juda städer och med dess konungar och furstar, för att så göra dem till en ödemark, och till ett föremål för häpnad och begabberi, och till ett exempel som man nämner, när man förbannar, såsom ock nu har skett;
vidare Farao, konungen i Egypten, med hans tjänare, hans furstar och allt hans folk,
så ock allt Erebs folk med alla konungar i Us' land och alla konungar i filistéernas land, både Askelon och Gasa och Ekron och kvarlevan i Asdod;
vidare Edom, Moab och Ammons barn;
vidare alla konungar i Tyrus, alla konungar i Sidon och konungarna i kustländerna på andra sidan havet;
vidare Dedan, Tema, Bus och alla dem som hava kantklippt hår;
vidare alla konungar i Arabien och alla konungar över Erebs folk, som bo i öknen,
så ock alla konungar i Simri, alla konungar i Elam och alla konungar i Medien,
slutligen alla konungar i nordlandet -- både dem som bo nära och dem som bo fjärran, den ene såväl som den andre -- och alla övriga riken i världen, utöver jordens yta.
Och Sesaks konung skall dricka efter dem.
Och du skall säga till dem: Så säger HERREN Sebaot, Israels Gud: Dricken, så att I bliven druckna, och spyn, och fallen omkull utan att kunna stå upp; ja, fallen, när det svärd kommer, som jag skall sända bland eder. --
Men om de icke vilja taga emot kalken ur din hand och dricka, så säg till dem: Så säger HERREN Sebaot: I måsten dricka.
Ty se, med den stad som är uppkallad efter mitt namn skall jag begynna hemsökelsen.
Skullen då I bliva ostraffade?
Nej, I skolen icke bliva ostraffade, utan jag skall båda upp ett svärd mot jordens alla inbyggare, säger HERREN Sebaot.
Och du skall profetera för dem allt detta och säga till dem: HERREN upphäver ett rytande från höjden och från sin heliga boning låter han höra sin röst; ja, han upphäver ett högt rytande över sin ängd och höjer skördeskri, såsom en vintrampare, över alla jordens inbyggare.
Dånet höres intill jordens ända, ty HERREN har sak med folken, han går till rätta med allt kött; de ogudaktiga giver han till pris åt svärdet, säger HERREN.
Så säger HERREN Sebaot: Se, en olycka går fram ifrån det ena folket till det andra, och ett stort oväder stiger upp från jordens yttersta ända.
Och de som bliva slagna av HERREN på den tiden skola ligga strödda från jordens ena ända till den andra; man skall icke hålla dödsklagan efter dem eller samla dem tillhopa och begrava dem, utan de skola bliva gödsel på marken.
Jämren eder, I herdar, och klagen; vältren eder på marken, I väldige i hjorden; ty tiden är inne, att I skolen slaktas.
I skolen bliva förskingrade, I skolen komma på fall, såsom det händer jämväl ett dyrbart kärl.
Då finnes icke mer någon undflykt för herdarna, icke mer någon räddning för de väldige i hjorden.
Hör huru herdarna ropa, huru de väldige i hjorden jämra sig!
Ty HERREN ödelägger deras betesmark,
och de fredliga ängderna förgöras genom HERRENS vredes glöd.
Han drager ut såsom ett lejon ur sitt snår.
Ja, deras land bliver en ödemark under förhärjelsens glöd, under hans vredes glöd.
I begynnelsen av Jojakims, Josias sons, Juda konungs, regering kom detta ord från HERREN; han sade:
Så säger HERREN: Ställ dig i förgården till HERRENS hus och tala mot alla Juda städer, från vilka man kommer för att tillbedja i HERRENS hus, tala alla de ord som jag har bjudit dig tala till dem; tag intet därifrån.
Kanhända skola de då höra och vända om, var och en från sin onda väg; då vill jag ångra det onda som jag har i sinnet att göra med dem för deras onda väsendes skull.
Du skall säga till dem: Så säger HERREN: Om I icke viljen höra mig och vandra efter den lag som jag har förelagt eder,
och höra vad mina tjänare profeterna tala -- de som jag titt och ofta sänder till eder, fastän I icke viljen höra --
då skall jag göra med detta hus såsom jag gjorde med Silo, och skall låta denna stad för alla jordens folk bliva ett exempel som man nämner, när man förbannar.
Och prästerna och profeterna och allt folket hörde Jeremia tala dessa ord i HERRENS hus.
Och när Jeremia hade slutat att tala allt vad HERREN hade bjudit honom tala till allt folket, grepo honom prästerna och profeterna och allt folket och sade: »Du måste döden dö.
Huru djärves du profetera i HERRENS namn och säga: 'Det skall gå detta hus likasom det gick Silo, och denna stad skall ödeläggas, så att ingen mer bor däri'?»
Och allt folket församlade sig mot Jeremia i HERRENS hus.
Då nu Juda furstar hörde detta, gingo de från konungshuset upp till HERRENS hus och satte sig vid ingången till HERRENS nya port.
Då sade prästerna och profeterna till furstarna och till allt folket sålunda: »Denne man förtjänar döden, ty han har profeterat mot denna stad, såsom I haven hört med egna öron.»
Men Jeremia svarade alla furstarna och allt folket och sade: »Det är HERREN som har sänt mig att profetera mot detta hus och denna stad allt det som I haven hört.
Så bättren nu edert leverne och edert väsende, och hören HERRENS, eder Guds, röst; då vill HERREN ångra det onda som han har talat mot eder.
Och vad mig angår, så är jag i eder hand; gören med mig vad eder gott och rätt synes.
Men det skolen I veta, att om I döden mig, så dragen I oskyldigt blod över eder och över denna stad och dess invånare; ty det är i sanning HERREN som har sänt mig till eder att tala allt detta inför eder.»
Då sade furstarna och allt folket till prästerna och profeterna: »Denne man förtjänar icke döden, ty i HERRENS, vår Guds, namn har han talat till oss.
Och några av de äldste i landet stodo upp och sade till folkets hela församling sålunda:
»Morastiten Mika profeterade i Hiskias, Juda konungs, tid och sade till hela Juda folk: 'Så säger HERREN Sebaot: Sion skall varda upplöjt till en åker, och Jerusalem skall bliva en stenhop och tempelberget en skogbevuxen höjd.'
Men lät väl Hiskia, Juda konung, med hela Juda, döda honom?
Fruktade han icke i stället HERREN och bönföll inför honom, så att HERREN ångrade det onda som han hade beslutit över dem, medan tvärtom vi nu stå färdiga att draga över oss själva så mycket ont?»
Där var ock en annan man, Uria, Semajas son, från Kirjat-Hajearim, som profeterade i HERRENS namn; och han profeterade mot denna stad och detta land alldeles såsom Jeremia hade gjort.
När då konung Jojakim med alla sina hjältar och alla furstar hörde vad han sade, ville han döda honom.
Men när Uria fick höra härom, blev han förskräckt och flydde och kom till Egypten.
Då sände konung Jojakim några män till Egypten, nämligen Elnatan, Akbors son, och några andra med honom, in i Egypten.
Och dessa hämtade Uria ut ur Egypten och förde honom till konung Jojakim; och denne lät dräpa honom med svärd, och lät så kasta hans döda kropp på den allmänna begravningsplatsen.
Men Ahikam, Safans son, höll sin hand över Jeremia, så att man icke lämnade honom i folkets hand till att dödas.
I begynnelsen av Jojakims, Josias sons, Juda konungs, regering kom detta ord till Jeremia från HERREN;
han sade: Så har HERREN sagt till mig: Gör dig band och ok och sätt detta på din hals.
Sänd det sedan till konungen i Edom, konungen i Moab, konungen över Ammons barn, konungen i Tyrus och konungen i Sidon, genom de sändebud som hava kommit till Sidkia, Juda konung, i Jerusalem.
Och bjud dem med dessa ord framföra sitt budskap till sina herrar: Så säger HERREN Sebaot, Israels Gud: Så skolen I säga till edra herrar:
Jag är den som genom min stora kraft och min uträckta arm har gjort jorden, med de människor och djur som äro på jorden; och jag giver den åt vem jag vill.
Så giver jag nu alla dessa länder i min tjänare Nebukadnessars, den babyloniske konungens, hand; ja ock markens djur giver jag honom, för att de må tjäna honom.
Och alla folk skola vara honom och hans son och hans sonson underdåniga, till dess att också för hans land tiden är inne, att mäktiga folk och stora konungar skola göra honom sig underdånig.
Och det folk och det rike som icke vill vara honom, Nebukadnessar, konungen i Babel, underdånigt, och som icke vill giva sin hals under den babyloniske konungens ok, det folket skall jag hemsöka med svärd, hungersnöd och pest, säger HERREN, till dess att jag har förgjort dem genom hans hand.
Därför mån I icke höra på edra profeter och spåman, på edra drömmar, på edra teckentydare och trollkarlar, när dessa säga till eder: »I skolen icke komma att tjäna konungen i Babel»;
ty de profetera lögn för eder, och komma så åstad att I bliven förda långt undan från edert land, i det jag måste driva eder bort, så att I förgåns.
Men det folk som böjer sin hals under den babyloniske konungens ok och tjänar honom, det skall jag låta få ro i sitt land, säger HERREN, så att de kunna bruka det och bo däri.
Till Sidkia, Juda konung, talade jag på alldeles samma sätt; jag sade: Böjen eder hals under den babyloniske konungens ok, och tjänen honom och hans folk, så skolen I få leva.
Icke viljen I dö, du och ditt folk, genom svärd, hunger och pest, såsom HERREN har sagt att det skall ske med det folk som icke vill tjäna konungen i Babel?
Hören alltså icke på de profeters ord, som säga till eder »I skolen icke komma att tjäna konungen i Babel»; ty de profetera lögn för eder.
Jag har icke sänt dem, säger HERREN; det är de själva som profetera lögn i mitt namn, och de komma så åstad att jag måste driva eder bort, så att I förgåns, jämte de profeter som profetera för eder.
Och till prästerna och till hela detta folk talade jag och sade: Så säger HERREN: Hören icke på edra profeters ord, när de profetera för eder och säga: »Se, de kärl som höra till HERRENS hus skola nu snart föras tillbaka från Babel»; ty de profetera lögn för eder.
Hören icke på dem, utan tjänen konungen i Babel, så skolen I få leva.
Icke viljen I att denna stad skall bliva ödelagd?
Om de verkligen äro profeter och hava HERRENS ord, så må de lägga sig ut hos HERREN Sebaot, för att de kärl som ännu äro kvar i HERRENS hus och i Juda konungs hus och i Jerusalem icke också må föras bort till Babel
Ty så säger HERREN Sebaot om pelarna och havet och bäckenställen och det övriga som ännu är kvar här i staden,
därför att Nebukadnessar, konungen i Babel, icke tog det med sig, när han förde bort Jekonja, Jojakims son, Juda konung, från Jerusalem till Babel, jämte alla ädlingar i Juda och Jerusalem --
ja, så säger HERREN Sebaot, Israels Gud, om det som ännu är kvar här i HERRENS hus och i Juda konungs hus och i Jerusalem:
Till Babel skall det föras, och där skall det förbliva ända till den dag då jag ser därtill, säger HERREN, och för det upp till denna plats igen.
Men samma år, i begynnelsen av Sidkias, Juda konungs, regering, i femte månaden av hans fjärde regeringsår, talade profeten Hananja, Assurs son, från Gibeon, så till mig i HERRENS hus, i prästernas och allt folkets närvaro; han sade:
»Så säger HERREN Sebaot, Israels Gud: Jag skall sönderbryta den babyloniske konungens ok.
Inom två års tid skall jag föra tillbaka till denna plats alla de kärl i HERRENS hus, som Nebukadnessar, konungen i Babel, har tagit bort ifrån denna plats och fört till Babel.
Och Jekonja, Jojakims son, Juda konung, och alla fångar ifrån Juda, som hava kommit till Babel, skall jag föra tillbaka till denna plats, säger HERREN; ty jag skall sönderbryta den babyloniske konungens ok.»
Men profeten Jeremia svarade profeten Hananja, i närvaro av prästerna och allt det folk som stod i HERRENS hus;
profeten Jeremia sade: »Amen.
Så göre HERREN.
Det som du har profeterat må HERREN uppfylla, i det att han för tillbaka från Babel till denna plats de kärl som funnos i HERRENS hus, så ock alla fångarna.
Men hör dock detta ord som jag vill tala inför dig och allt folket.
Forna tiders profeter, de som hava varit före mig och dig, hava mot mäktiga länder och stora riken profeterat om krig, olycka och pest.
Därför, om nu en profet profeterar om lycka, så kan man först då när den profetens ord går i fullbordan veta att han är en profet som HERREN i sanning har sänt.»
Då tog profeten Hananja oket från profeten Jeremias hals och bröt sönder det.
Och Hananja sade i allt folkets närvaro: »Så säger HERREN: Just så skall jag inom två års tid bryta sönder den babyloniske konungen Nebukadnessars ok och taga det från alla folkens hals.»
Men profeten Jeremia gick sin väg.
Sedan, efter det att profeten Hananja hade brutit sönder oket och tagit det från profeten Jeremias hals, kom HERRENS ord till Jeremia; han sade:
»Gå åstad och säg till Hananja: Så säger HERREN: Ett ok av trä har du brutit sönder, men i dess ställe har du skaffat ett ok av järn.
Ty så säger HERREN Sebaot, Israels Gud: Ett ok av järn skall jag sätta på alla dessa folks hals, för att de må tjäna Nebukadnessar, konungen i Babel; ty honom skola de tjäna.
Ja ock markens djur har jag givit honom.»
Och profeten Jeremia sade ytterligare till profeten Hananja: »Hör, du Hananja: HERREN har icke sänt dig; du har förlett detta folk att sätta sin lit till lögn.
Därför säger HERREN så: Se, jag skall taga dig bort ifrån jorden.
I detta år skall du dö, eftersom du har predikat avfall från HERREN.»
Och samma år, i sjunde månaden, dog profeten Hananja.
Detta är vad som stod i det brev som profeten Jeremia sände från Jerusalem till de äldste som ännu levde kvar i fångenskapen, och till prästerna och profeterna och allt folket, dem som Nebukadnessar hade fört bort ifrån Jerusalem till Babel,
sedan konung Jekonja hade givit sig fången i Jerusalem, jämte konungamodern och hovmännen, Judas och Jerusalems furstar, så ock timmermännen och smederna.
Han sände brevet genom Eleasa, Safans son, och Gemarja, Hilkias son, när Sidkia, Juda konung, sände dessa till Babel, till Nebukadnessar, konungen i Babel; det lydde så:
Så säger HERREN Sebaot, Israels Gud, till alla de fångar som jag har låtit föra bort ifrån Jerusalem till Babel:
Byggen hus och bon i dem; planteren trädgårdar och äten deras frukt.
Tagen hustrur, och föden söner och döttrar; och tagen hustrur åt edra söner och given edra döttrar åt män, och må dessa föda söner och döttrar; och föröken eder där, och förminskens icke.
Och söken den stads bästa, dit jag har fört eder bort i fångenskap, och bedjen för den till HERREN; ty då det går den väl, så går det ock eder val.
Ty så säger HERREN Sebaot, Israels Gud: Låten icke bedraga eder av de profeter som äro bland eder, ej heller av edra spåman, och akten icke på de drömmar som I drömmen.
Ty man profeterar lögn för eder i mitt namn; jag har icke sänt dem, säger HERREN.
Ty så säger HERREN: Först när sjuttio år hava gått till ända i Babel, skall jag se till eder och uppfylla på eder mitt löftesord att föra eder tillbaka till denna plats.
Jag vet väl vilka tankar jag har för eder, säger HERREN, nämligen fridens tankar och icke ofärdens, till att giva eder en framtid och ett hopp.
Och I skolen åkalla mig och gå åstad och bedja till mig, och jag vill höra på eder.
I skolen söka mig, och I skolen ock finna mig, om I frågen efter mig av allt edert hjärta.
Ty jag vill låta mig finnas av eder, säger HERREN; och jag skall åter upprätta eder och skall församla eder från alla de folk och alla de arter till vilka jag har drivit eder bort, säger HERREN; och jag skall låta eder komma tillbaka till denna plats, varifrån jag har låtit föra eder bort i fångenskap.
Detta skriver jag, därför att I sägen: »HERREN har låtit profeter uppstå åt oss i Babel.»
Ty så säger HERREN om den konung som sitter på Davids tron, och om allt det folk som bor i denna stad, edra bröder som icke hava med eder gått bort i fångenskap,
ja, så säger HERREN Sebaot: Se, jag skall sända mot dem svärd, hungersnöd och pest, och låta dem räknas lika med odugliga fikon, som äro så usla att man icke kan äta dem.
Ja, jag skall förfölja dem med svärd, hungersnöd och pest, och göra dem till en varnagel för alla riken på jorden, till ett exempel som man nämner, när man förbannar, till ett föremål för häpnad, begabberi och smälek bland alla de folk till vilka jag skall driva dem bort --
detta därför att de icke ville höra mina ord, säger HERREN, när jag titt och ofta sände till dem mina tjänare profeterna.
Ty I villen ju icke höra, säger HERREN.
Men hören nu I HERRENS ord, alla I fångna som jag från Jerusalem har sänt bort till Babel:
Så säger HERREN Sebaot, Israels Gud, om Ahab, Kolajas son, och om Sidkia, Maasejas son, som i mitt namn profetera lögn för eder: Se, jag skall giva dem i Nebukadressars, den babyloniske konungens, hand, och han skall låta dräpa dem inför edra ögon.
Och alla fångar ifrån Juda, som äro i Babel, skola från dem hämta ett förbannelsens ord; de skola »HERREN göre med dig såsom med Sidkia och Ahab, vilka Babels konung lät steka i eld.»
De hava ju gjort vad som är ens galenskap i Israel, de hava begått äktenskapsbrott med varandras hustrur och hava fört lögnaktigt tal i mitt namn, sådant som jag icke hade bjudit dem.
Jag är den som vet det och betygar det, säger HERREN.
Och till nehelamiten Semaja skall du säga sålunda:
Så säger HERREN Sebaot, Israels Gud: Du har i ditt namn sänt brev till allt folket i Jerusalem och till prästen Sefanja, Maasejas son, och till alla de andra prästerna, så lydande:
»HERREN har satt dig till präst i prästen Jojadas ställe, för att i HERRENS hus skall finnas tillsyningsmän över alla vanvettingar som profetera, så att du kan sätta sådana i stock och halsjärn.
Varför har du då icke näpst Jeremia från Anatot, som profeterar för eder?
Därigenom att du har underlåtit detta har han kunnat sända bud till oss i Babel och låta säga: 'Ännu är lång tid kvar, byggen eder hus och bon i dem, och planteren trädgårdar och äten deras frukt.'»
Och prästen Sefanja har läst upp detta brev för profeten Jeremia.
Och nu har HERRENS ord kommit till Jeremia, han har sagt:
Sänd bud till alla de fångna och låt säga dem: Så säger HERREN om nehelamiten Semaja: Eftersom Semaja, utan att vara sänd av mig, har profeterat för eder och förlett eder att sätta eder lit till lögn,
därför säger HERREN så: Se, jag skall hemsöka nehelamiten Semaja och hans avkomlingar.
Ingen av dem skall få bo ibland detta folk, och han skall icke få se det goda som jag vill göra med mitt folk, säger HERREN.
Ty han har predikat avfall från HERREN.
Detta är det ord som kom till Jeremia från HERREN; han sade:
Så säger HERREN, Israels Gud: Teckna upp åt dig i en bok alla de ord som jag har talat till dig.
Ty se, dagar skola komma, säger HERREN, då jag åter skall upprätta mitt folk, Israel och Juda, säger HERREN, och låta dem komma tillbaka till det land som jag har givit åt deras fäder; och de skola taga det i besittning.
Och detta är vad HERREN har talat om Israel och Juda.
Så säger HERREN: Ett förfärans rop fingo vi höra; förskräckelse utan någon räddning!
Frågen efter och sen till: pläga då män föda barn?
Eller varför ser jag alla män hålla sina händer på länderna såsom kvinnor i barnsnöd, och varför hava alla ansikten blivit så dödsbleka?
Ve!
Detta är en stor dag, en sådan att ingen är den lik.
Ja, en tid av nöd är inne för Jakob; dock skall han bliva frälst därur.
Och det skall ske på den tiden, Säger HERREN Sebaot, att jag skall bryta sönder oket och taga det från din hals och slita av dina band.
Ja, inga främmande skola längre tvinga honom att tjäna sig,
utan han skall få tjäna HERREN, sin Gud, och David, sin konung, ty honom skall jag låta uppstå åt dem.
Så frukta nu icke, du min tjänare Jakob, säger HERREN. och var ej förfärad du Israel; ty se, jag skall frälsa dig ur det avlägsna landet, och dina barn ur deras fångenskaps land.
Och Jakob skall få komma tillbaka och leva i ro och säkerhet, och ingen skall förskräcka honom.
Ty jag är med dig, säger HERREN, till att frälsa dig.
Ja, jag skall göra ände på alla de folk; bland vilka jag har förstrött dig; men på dig vill jag icke alldeles göra ände, jag vill blott tukta dig med måtta; ty alldeles ostraffad kan jag ju ej låta dig bliva.
Ty så säger HERREN: Ohelbar är din skada, oläkligt det sår du har fått.
Ingen tager sig an din sak, så att han sköter ditt sår; ingen helande läkedom finnes för dig.
Alla dina älskare hava förgätit dig; de fråga icke efter dig.
Ty såsom man slår en fiende, så har jag slagit dig, med grym tuktan, därför att din missgärning var så stor och dina synder så många.
Huru kan du klaga över din skada, över att bot ej finnes för din plåga?
Därför att din missgärning var så stor och dina synder så många, har jag gjort dig detta.
Så skola då alla dina uppätare nu bliva uppätna, och alla dina ovänner skola allasammans gå i fångenskap; dina skövlare skola varda skövlade, och alla dina plundrare skall jag lämna till plundring.
Ty jag vill hela dina sår och läka dig från de slag du har fått, säger HERREN, då man nu kallar dig »den fördrivna», »det Sion som ingen frågar efter».
Så säger HERREN: Se, jag skall åter upprätta Jakobs hyddor och förbarma mig över hans boningar; staden skall åter bliva uppbyggd på sin höjd, och palatset skall stå på sin rätta plats.
Ifrån folket skall ljuda tacksägelse och rop av glada människor.
Jag skall föröka dem, och de skola icke förminskas; jag skall låta dem komma till ära, och de skola ej aktas ringa.
Hans söner skola varda såsom fordom, hans menighet skall bestå inför mig, jag skall hemsöka alla hans förtryckare.
Hans väldige skall stamma från honom själv, och hans herre skall utgå från honom själv, och honom skall jag låta komma mig nära och nalkas mig; ty vilken annan vill våga sitt liv med att nalkas mig? säger HERREN.
Och I skolen vara mitt folk och jag skall vara eder Gud.
Se, en stormvind från HERREN är här, hans förtörnelse bryter fram, en härjande storm!
Över de ogudaktigas huvuden virvlar den ned.
HERRENS vredes glöd skall icke upphöra, förrän han har utfört och fullbordat sitt hjärtas tankar; i kommande dagar skolen I förnimma det.
På den tiden, säger HERREN, skall jag vara alla Israels släkters Gud, och de skola vara mitt folk.
Så säger HERREN: Det folk som undslipper svärdet finner nåd i öknen; Israel får draga åstad dit där det får ro.
Fjärran ifrån uppenbarade sig HERREN för mig: »Ja, med evig kärlek har jag älskat dig; därför låter jag min nåd förbliva över dig.
Ännu en gång skall jag upprätta dig, så att du varder upprättad, du jungfru Israel; ännu en gång skall du få utrusta dig med puka och draga ut i dans bland dem som göra sig glada.
Ännu en gång skall du få plantera vingårdar på Samariens berg, och planteringsmännen skola själva skörda frukten.
Ty en dag kommer, då vaktare skola ropa på Efraims berg: 'Upp, låt oss draga till Sion, upp till HERREN, vår Gud.'»
Ty så säger HERREN: Jublen i glädje över Jakob, höjen fröjderop över honom som är huvudet bland folken, Låten lovsång ljuda och sägen: HERRE, giv frälsning åt ditt folk, åt kvarlevan av Israel.»
Ja, jag skall föra dem från nordlandet och församla dem från jordens yttersta ända -- bland dem både blinda och halta, både havande kvinnor och barnaföderskor; i en stor skara skola de komma hit tillbaka.
Under gråt skola de komma, men jag skall leda dem, där de gå bedjande fram; Jag skall föra dem till vattenbäckar, på en jämn väg, där de ej skola stappla.
Ty jag har blivit en fader för Israel, och Efraim är min förstfödde son.
Hören HERRENS ord, I hednafolk, och förkunnen det i havsländerna i fjärran; sägen: Han som förskingrade Israel skall ock församla det och bevara det, såsom en herde sin hjord.
Ty HERREN skall förlossa Jakob och lösköpa honom ur den övermäktiges hand.
Och de skola komma och jubla på Sions höjd och strömma dit där HERRENS goda är, dit där man får säd, vin och olja och unga hjordar av får och fä; deras själ skall vara lik en vattenrik trädgård, och de skola icke vidare försmäkta.
Då skola jungfrurna förlusta sig med dans; unga och gamla skola glädja sig tillsammans.
Jag skall förvandla deras sorg i fröjd, trösta dem och glädja dem efter deras bedrövelse.
Och prästerna skall jag vederkvicka med feta rätter; och mitt folk skall bliva mättat av mitt goda, säger HERREN.
Så säger HERREN: Ett rop höres i Rama, klagan och bitter gråt; det är Rakel som begråter sina barn, hon vill icke låta trösta sig i sorgen över att hennes barn icke mer äro till.
Men så säger HERREN: Hör upp med din högljudda gråt, och låt dina ögon icke mer fälla tårar; ty ditt verk skall få sin lön, säger HERREN, och de skola vända tillbaka från sina fienders land.
Ja, det finnes ett hopp för din framtid, säger HERREN; dina barn skola vända tillbaka till sitt land.
Jag har nogsamt hört huru Efraim klagar: »Du har tuktat mig, ja, jag har blivit tuktad såsom en otämd kalv; tag mig nu åter, så att jag får vända åter; du är ju HERREN, min Gud.
Ty sedan jag har vänt mitt sinne, ångrar jag mig, och sedan jag har kommit till besinning, slår jag mig på länden; jag både blyges och skämmes, då jag nu bär min ungdoms smälek.»
Är då Efraim for mig en så dyrbar son, är han mitt älsklingsbarn, eftersom jag alltjämt tänker på honom, huru ofta jag än har måst hota honom?
Ja, så mycket ömkar sig mitt hjärta över honom; jag måste förbarma mig över honom, säger HERREN.
Sätt upp vägmärken för dig, res åt dig vägvisare; giv akt på vägen, på stigen där du vandrade.
Och vänd så tillbaka, du jungfru Israel, vänd tillbaka till dessa dina städer.
Huru länge skall du göra bukter hit och dit, du avfälliga dotter?
Se, HERREN vill skapa något nytt i landet: det bliver nu kvinnan som tager mannen i sitt beskärm.
Så säger HERREN Sebaot, Israels Gud: I Juda land med dess städer skall man ännu en gång, när jag åter har upprättat det, få säga det ordet: »HERREN välsigne dig, du rättfärdighetens boning, du heliga berg.»
Och Juda folk med alla sina städer skall samlat bo däri, åkermän jämte vandrande herdar.
Ty jag skall vederkvicka trötta själar, och alla försmäktande själar skall jag mätta.
(Härvid uppvaknade jag och såg mig om, och min sömn hade varit ljuvlig.)
Se, dagar skola komma, säger HERREN, då jag skall beså Israels land och Juda land med säd av människor och med säd av djur.
Och likasom jag har vakat över dem till att upprycka, nedbryta, fördärva, förgöra och plåga, så vill jag nu vaka över dem till att uppbygga och plantera, säger HERREN.
På den tiden skall man icke mer säga: »Fäderna hava ätit sura druvor, och barnens tänder bliva ömma därav.»
Nej, var och en skall dö genom sin egen missgärning; var man som äter sura druvor, hans tänder skola bliva ömma därav.
Se, dagar skola komma, säger HERREN, då jag skall sluta ett nytt förbund med Israels hus och med Juda hus;
icke ett sådant förbund som det jag slöt med deras fäder på den dag då jag tog dem vid handen till att föra dem ut ur Egyptens land det förbund med mig, som de bröto, fastän jag var deras rätte herre, säger HERREN.
Nej, detta är det förbund som jag skall sluta med Israels hus i kommande dagar, säger HERREN: Jag skall lägga min lag i deras bröst och i deras hjärtan skall jag skriva den, och jag skall vara deras Gud, och de skola vara mitt folk.
Då skola de icke mer behöva undervisa varandra, icke den ene brodern den andre, och säga: »Lär känna HERREN»; ty de skola alla känna mig, från den minste bland dem till den störste, säger HERREN.
Ty jag skall förlåta deras missgärning, och deras synd skall jag icke mer komma ihåg.
Så säger HERREN, han som har satt solen till att lysa om dagen och månen och stjärnorna till att lysa om natten, i ordnad gång, han som rör upp havet, så att dess böljor brusa, han vilkens namn är HERREN Sebaot:
Först när denna ordning icke mer består inför mig, säger HERREN, först då skall Israels släkt upphöra att inför mig alltjämt vara ett folk.
Ja, så säger HERREN: Först när himmelen varder uppmätt därovan och jordens grundvalar utrannsakade därnere, först då skall jag förkasta all Israels släkt, till straff för allt vad de hava gjort, säger HERREN.
Se, dagar skola komma, säger HERREN, då staden åter skall varda uppbyggd till HERRENS ära, från Hananeltornet intill Hörnporten.
Och mätsnöret skall vidare dragas rätt fram mot Garebshöjden och skall sedan vändas mot Goa.
Och hela lik- och askdalen och alla fälten intill bäcken Kidron och intill hörnet vid Hästporten österut skola vara helgade åt HERREN.
Aldrig mer skall där tima någon omstörtning eller någon förstöring.
Detta är det ord som från HERREN kom till Jeremia i Sidkias, Juda konungs, tionde regeringsår, vilket var Nebukadressars adertonde regeringsår.
Vid den tiden belägrade den babyloniske konungens här Jerusalem, och profeten Jeremia låg då fången i fängelsegården i Juda konungs hus.
Ty Sidkia, Juda konung, hade låtit spärra in honom, i det han sade: »Huru djärves du profetera och säga: 'Så säger HERREN: Se, jag skall giva denna stad i de babyloniske konungens hand, och han skall intaga den.
Och Sidkia, Juda konung, skall icke undkomma kaldéernas hand, utan skall förvisso bliva given i den babyloniske konungens hand, så att han nödgas muntligen tala med honom och stå inför honom, öga mot öga.
Och Sidkia skall av honom föras till Babel och skall förbliva där, till dess jag ser till honom, säger HERREN.
När I striden mot kaldéerna, skolen I icke hava någon framgång.»
Och Jeremia sade: »HERRENS ord kom till mig; han sade:
Se, Hanamel, din farbroder Sallums son, skall komma till dig och säga: 'Köp du min åker i Anatot, ty du har såsom bördeman rätt att köpa den.'»
Och Hanamel, min farbroders son, kom till mig i fängelsegården, såsom HERREN hade sagt, och sade till mig: »Köp min åker i Anatot, i Benjamins land, ty du har arvsrätt därtill och är bördeman; så köp den då åt dig.»
Då förstod jag att det var HERRENS ord
och köpte åkern av Hanamel, min farbroders son, i Anatot, och vägde upp penningarna åt honom, sjutton siklar silver.
Jag skrev ett köpebrev och förseglade det och tillkallade vittnen och vägde upp penningarna på en våg.
Och jag tog köpebrevet, såväl det förseglade, som innehöll avtalet och de särskilda bestämmelserna, som ock det öppna brevet,
och gav köpebrevet åt Baruk, son till Neria, son till Mahaseja, i närvaro av min frände Hanamel och de vittnen som hade underskrivit köpebrevet, och alla andra judar som voro tillstädes i fängelsegården.
Och jag bjöd Baruk, i deras närvaro, och sade:
Så säger HERREN Sebaot, Israels Gud: Tag du dessa brev, både detta förseglade köpebrev och detta öppna brev, och lägg dem i ett lerkärl, för att de må vara i behåll för lång tid.
Ty så säger HERREN Sebaot, Israels Gud: Ännu en gång skall man komma att i detta land köpa hus och åkrar och vingårdar.»
Och sedan jag hade givit köpebrevet åt Baruk, Nerias son, bad jag till HERREN och sade:
»Ack Herre, HERRE, du är ju den som har gjort himmel och jord genom din stora kraft och din uträckta arm.
Intet är så underbart att du icke skulle förmå det,
du som gör nåd med tusenden och vedergäller fädernas missgärning i deras barns sköte efter dem; du store och väldige Gud, vilkens namn är HERREN Sebaot;
du som är stor i råd och mäktig i gärningar; du vilkens ögon äro öppna över människobarnens alla vägar, så att du giver åt var och en efter hans vägar och efter hans gärningars frukt;
du som gjorde tecken och under i Egyptens land, och som har gjort sådana intill denna dag, både i Israel och bland andra människor, och som har gjort dig ett namn, som är detsamma än i dag.
Du förde ditt folk Israel ut ur Egyptens land med tecken och under, med stark hand och uträckt arm, och genom stor förskräckelse.
Och du gav dem detta land, som du med ed hade lovat deras fäder att giva dem, ett land som flyter av mjölk och honung.
Och de kommo och togo det i besittning, men de ville icke höra din röst och vandrade icke efter din lag; de gjorde intet av det du hade bjudit dem att göra.
Därför lät du all denna olycka vederfaras dem.
Se, belägringsvallarna gå redan så långt fram mot staden, att man kan intaga den och genom svärd, hungersnöd och pest är staden given i de kaldeiska belägrarnas hand.
Vad du hotade med, det har skett, och du har det nu inför dina ögon.
Och likväl, fastän staden är given i kaldéernas hand, sade du, Herre HERRE, till mig: 'Köp du åkern för penningar, och tag vittnen därpå'!»
Och HERRENS ord kom till Jeremia han sade: Se,
jag är HERREN, allt kötts Gud; skulle något vara så underbart att jag icke förmådde det?
Därför säger HERREN så: Se, jag vill giva denna stad i kaldéernas och Nebukadressars, den babyloniske konungens, hand, och han skall intaga den.
Och kaldéerna, som belägra denna stad, skola komma och tända eld på staden och bränna upp den, tillika med de hus på vilkas tak man har tänt offereld åt Baal och utgjutit drickoffer åt andra gudar, till att förtörna mig.
Ty allt ifrån sin ungdom hava Israels barn och Juda barn allenast gjort vad ont är i mina ögon; ja, Israels barn hava med sina händers verk berett mig allenast förtörnelse, säger HERREN.
Ty allt ifrån den dag då denna stad byggdes ända till nu har den uppväckt min vrede och förtörnelse, så att jag måste förkasta den från mitt ansikte,
för all den ondskas skull som Israels barn och Juda barn med sina konungar, furstar, präster och profeter, både Juda män och Jerusalems invånare, hava bedrivit, till att förtörna mig.
De vände ryggen till mig och icke ansiktet; och fastän de titt och ofta blevo varnade, ville de icke höra och taga emot tuktan.
De satte upp sina styggelser i det hus som är uppkallat efter mitt namn och orenade det så;
och Baalshöjderna i Hinnoms sons dal byggde de upp, för att där offra sina söner och döttrar åt Molok, fastän jag aldrig hade bjudit dem att göra sådan styggelse eller ens tänkt mig något sådant; och så förledde de Juda till synd.
Men så säger nu HERREN, Israels Gud, om denna stad, som I menen vara genom svärd, hungersnöd och pest given i den babyloniske konungens hand:
Se, jag skall församla dem ur alla de länder till vilka jag i min vrede och harm och stora förtörnelse har fördrivit dem, och jag skall föra dem tillbaka till denna plats och låta dem bo bär i trygghet.
Och de skola vara mitt folk, och jag skall vara deras Gud.
Och jag skall giva dem alla ett och samma hjärta och lära dem en och samma väg, så att de frukta mig beständigt; för att det må gå dem väl, och deras barn efter dem.
Och jag skall sluta med dem ett evigt förbund, så att jag icke upp hör att följa dem och göra dem gott; och min fruktan skall jag ingiva i deras hjärtan, så att de icke vika av ifrån mig.
Och jag skall hava min fröjd i att göra dem gott, och skall plantera dem i detta land med trofasthet, av allt mitt hjärta och all min själ.
Ty så säger HERREN: Likasom jag har låtit all denna stora olycka komma över detta folk, så skall jag ock låta allt det goda som jag lovade dem komma dem till del.
Och man skall komma att köpa åkrar i detta land, om vilket I sägen att det är en ödemark, där varken människor eller djur kunna bo, och att det är givet i kaldéernas hand.
Ja, åkrar skall man köpa för penningar, och man skall skriva och försegla köpebrev och tillkalla vittnen i Benjamins land, i Jerusalems omnejd och i Juda städer, både i Bergsbygdens och i Låglandets och i Sydlandets städer; ty jag skall åter upprätta dem, säger HERREN.
Och HERRENS ord kom till Jeremia för andra gången, medan han ännu var inspärrad i fängelsegården; han sade:
Så säger HERREN, han som ock utför sitt verk, HERREN, som bereder det för att låta det komma till stånd, han vilkens namn är HERREN:
Ropa till mig, så vill jag svara dig och förkunna för dig stora och förunderliga ting, som du icke känner.
Ty så säger HERREN, Israels Gud, om husen i denna stad och om Juda konungars hus, som nu brytas ned för belägringsvallarna och värden:
Man har kommit hitin för att strida med kaldéerna, och man skall så fylla husen med döda kroppar av människor som jag har slagit i min vrede och förtörnelse, människor som genom all sin ondska hava vållat att jag har måst dölja mitt ansikte för denna stad.
Dock, jag skall hela dess sår och skaffa läkedom och läka dem, och jag skall låta dem skåda frid och trygghet i överflöd.
Och jag skall åter upprätta Juda och Israel och uppbygga dem, så att de bliva såsom förut.
Och jag skall rena dem från all missgärning varmed de hava syndat mot mig, och förlåta alla missgärningar genom vilka de hava syndat mot mig och avfallit från mig.
Och staden skall bliva mig till fröjd och berömmelse, och till lov och ära inför alla jordens folk, när de få höra allt det goda som jag gör med dem; och de skola förskräckas och darra vid åsynen av all den lycka och all den framgång som jag bereder henne.
Så säger HERREN: På denna plats, om vilken I sägen att den är så öde att varken människor eller djur kunna bo där, ja, här i Juda städer och på Jerusalems gator, som äro så ödelagda att inga människor, inga invånare, inga djur där finnas,
här skall man ännu en gång höra fröjderop och glädjerop, rop för brudgum och rop för brud, rop av människor som säga: »Tacken HERREN Sebaot, ty HERREN är god, ty hans nåd varar evinnerligen», och av människor som frambära lovoffer i HERRENS hus.
Ty jag vill åter upprätta landet, så att det bliver såsom förut, säger HERREN.
Så säger HERREN Sebaot: På denna plats, som nu är så öde att varken människor eller ens djur kunna bo här, ja ock i alla hithörande städer, här skola åter en gång finnas betesmarker där herdar kunna låta sina hjordar lägra sig.
I Bergsbygdens, Låglandets och Sydlandets städer, i Benjamins land i Jerusalems omnejd och i andra Juda städer skola ännu en gång hjordar draga fram, förbi herdar som räkna dem, säger HERREN.
Se, dagar skola komma, säger HERREN, då jag skall uppfylla det löftesord som jag har talat om Israels hus och angående Juda hus.
I de dagarna och på den tiden skall jag låta en rättfärdig telning växa upp åt David.
Han skall skaffa rätt och rättfärdighet på jorden.
I de dagarna skall Juda varda frälst och Jerusalem bo i trygghet; och man skall kalla det så: HERREN vår rättfärdighet.
Ty så säger HERREN: Aldrig skall den tid komma, då icke en avkomling av David sitter på Israels hus' tron,
aldrig den tid då icke en avkomling av de levitiska prästerna gör tjänst inför mig och alla dagar bär fram brännoffer och förbränner spisoffer och anställer slaktoffer.
Och HERRENS ord kom till Jeremia; han sade:
Så säger HERREN: Först när I gören om intet mitt förbund med dagen och mitt förbund med natten, så att det icke bliver dag och natt i rätt tid,
först då skall mitt förbund med min tjänare David bliva om intet, så att icke längre en avkomling av honom sitter såsom konung på hans tron, och först då mitt förbund med de levitiska prästerna, som göra tjänst åt mig.
Lika oräknelig som himmelens härskara är, och lika otalig som sanden är i havet, lika talrik skall jag låta min tjänare Davids säd bliva och lika många leviterna, som göra tjänst åt mig.
Och HERRENS ord kom till Jeremia; han sade:
Har du icke märkt huru detta folk talar och säger: »De båda släkter som HERREN utvalde, dem har han förkastat»?
Och så säga de föraktligt om mitt folk att det icke mer synes dem vara ett folk.
Men så säger HERREN: Om mitt förbund med dag och natt icke är beståndande, och om jag icke har stadgat en fast ordning för himmel och jord,
allenast då skall jag förkasta Jakobs och Davids, min tjänares, säd, så att jag icke mer av hans säd tager dem som skola råda över Abrahams, Isaks och Jakobs säd.
Ty jag skall åter upprätta dem och förbarma mig över dem.
Detta är det ord som kom till Jeremia från HERREN, när Nebukadressar, konungen i Babel, med hela sin här och med alla de riken på jorden, som lydde under hans välde, och med alla folk angrep Jerusalem och alla dess lydstäder; han sade:
Så säger HERREN, Israels Gud: Gå åstad och säg till Sidkia, Juda konung, ja, säg till honom: Så säger HERREN: Se, jag skall giva denna stad i den babyloniske konungens hand, och han skall bränna upp den i eld.
Och du själv skall icke kunna undkomma hans hand, utan skall förvisso bliva gripen och given i hans hand, så att du nödgas stå inför konungen i Babel, öga mot öga; och han skall muntligen tala med dig, och du skall komma till Babel.
Men hör HERRENS ord, du Sidkia, Juda konung: Så säger HERREN om dig: Du skall icke dö genom svärd.
Nej, i frid skall du dö; och likasom man har anställt förbränning till dina fäders, de förra konungarnas, ära, deras som hava varit före dig, så skall man ock anställa förbränning till din ära och hålla dödsklagan efter dig: »Ack ve, Herre!»
Ty detta har jag talat, säger HERREN.
Och profeten Jeremia talade till Sidkia, Juda konung, allt detta i Jerusalem,
under det att den babyloniske konungens här belägrade Jerusalem och allt som ännu återstod av städer i Juda, nämligen Lakis och Aseka; ty dessa voro de enda av Juda städer, som ännu voro kvar och voro befästa.
Detta är det ord som kom till Jeremia från HERREN, sedan konung Sidkia hade slutit ett förbund med allt folket i Jerusalem därom att de bland sig skulle utropa frihet,
så att var och en skulle släppa sin träl och sin trälinna fria, om det var en hebreisk man eller kvinna, på det att icke den ene juden skulle hava den andre till träl.
Och detta hörsammades av alla furstarna och allt folket, av dem som hade varit med om förbundet och lovat att var och en skulle släppa sin träl och sin trälinna fria, så att han icke mer skulle hava dem till trälar; de hörsammade det och släppte dem.
Men sedermera ändrade de sig och togo tillbaka de trälar och trälinnor som de hade släppt fria, och gjorde dem åter till trälar och trälinnor.
Då kom HERRENS ord till Jeremia från HERREN; han sade:
Så säger HERREN, Israels Gud: Jag själv slöt ett förbund med edra fäder på den tid då jag förde dem ut ur Egyptens land, ur träldomshuset; jag sade:
»När sju år äro förlidna, skall var och en av eder släppa sin broder, hebréen, som har sålt sig åt dig och tjänat dig i sex år; du skall då släppa honom fri ur din tjänst.»
Dock ville edra fäder icke höra på mig eller böja sina öron därtill.
Men I haven nyss vänt om och gjort vad rätt är i mina ögon, i det att I haven utropat frihet var och en för sin broder.
Och I haven härom slutit ett förbund inför mitt ansikte, i det hus som är uppkallat efter mitt namn.
Men nu haven I åter ändrat eder och ohelgat mitt namn och tagit tillbaka var och en sin träl och sin trälinna, dem som I haden släppt fria till att gå vart de ville; ja, I haven nu åter gjort dem till edra trälar och trälinnor.
Därför säger HERREN så: I haven icke hört på mig och utropat frihet var och en för sin broder och sin nästa.
Så utropar då jag, säger HERREN, för eder frihet att hemfalla åt svärd, pest och hungersnöd; ja, jag skall göra eder till en varnagel för alla riken på jorden.
Och de män som hava överträtt mitt förbund och icke hållit förpliktelserna vid det förbund de slöto inför mitt ansikte -- vid kalven som av dem blev huggen i två stycken, mellan vilka de gingo --
dessa män, nämligen Judas och Jerusalems furstar, hovmännen och prästerna och allt folket i landet, som gingo mellan styckena av kalven,
dem skall jag giva i deras fienders hand, i de mäns hand, som stå efter deras liv; och deras döda kroppar skola bliva mat åt himmelens fåglar och markens djur.
Och Sidkia, Juda konung, med hans furstar skall jag giva i deras fienders hand, i de mäns hand, som stå efter deras liv, och i händerna på den babyloniske konungens här, som nu har dragit bort ifrån eder.
Se, jag skall giva dem befallning, säger HERREN, att de åter skola draga mot denna stad och belägra den; och de skola då intaga den och bränna upp den i eld.
Och Juda städer skall jag göra till en ödemark, där ingen bor.
Detta är det ord som kom till Jeremia från HERREN i Jojakims, Josias sons, Juda konungs, tid; han sade
Gå bort till rekabiternas släkt och tala med dem, och för dem till HERRENS hus, in i en av kamrarna, och giv dem vin att dricka.
Då tog jag med mig Jaasanja, son till Jeremia, son till Habassinja, jämte hans bröder och alla hans söner och rekabiternas hela övriga släkt,
och förde dem till HERRENS hus, in i den kammare som innehades av sönerna till gudsmannen Hanan, Jigdaljas son, den kammare som ligger bredvid furstarnas, ovanom dörrvaktaren Maasejas, Sallums sons, kammare.
Och jag satte fram för rekabiternas släkt kannor, fulla med vin, så ock bägare, och sade till dem: »Dricken vin?»
Men de svarade: »Vi dricka icke vin.
Ty vår fader Jonadab, Rekabs son, har bjudit oss och sagt: 'I och edra barn skolen aldrig dricka vin;
och hus skolen I icke bygga, och säd skolen I icke så, och vingårdar skolen I icke plantera, ej heller äga sådana, utan I skolen bo i tält i all eder tid, för att I mån länge leva i det land där I bon såsom främlingar.'
Och vi hava hörsammat vår fader Jonadabs, Rekabs sons, befallning, i allt vad han har bjudit oss, så att vi med våra hustrur och våra söner och döttrar aldrig dricka vin,
ej heller bygga hus till att bo i, ej heller äga vingårdar eller åkrar eller säd.
Vi hava alltså bott i tält och hava hörsammat och gjort allt vad vår fader Jonadab har bjudit oss.
Men när Nebukadressar, konungen i Babel, drog upp och föll in i landet, sade vi: 'Välan, vi vilja begiva oss till Jerusalem, undan kaldéernas och araméernas här.'
Och så bosatte vi oss i Jerusalem.»
Och HERRENS ord kom till Jeremia; han sade:
Så säger HERREN Sebaot, Israels Gud: Gå åstad och säg till Juda män och till Jerusalems invånare: Skolen I då icke taga emot tuktan, så att I hören mina ord, säger HERREN?
Det bud som Jonadab, Rekabs son, gav sina barn, att de icke skulle dricka vin, det har blivit iakttaget, och ännu i dag dricka de icke vin, av hörsamhet mot sin faders bud.
Men själv har jag titt och ofta talat till eder, och I haven dock icke hörsammat mig.
Och titt och ofta har jag sänt till eder alla mina tjänare profeterna och låtit säga: »Vänden om, var och en från sin onda väg, och bättren edert väsende, och följen icke efter andra gudar, så att I tjänen dem; då skolen I få bo i det land som jag har givit åt eder och edra fäder.»
Men I böjden icke edert öra därtill och hörden icke på mig.
Eftersom nu detta folk icke har hörsammat mig, såsom Jonadabs, Rekabs sons, barn hava iakttagit det bud som deras fader gav dem,
därför säger HERREN, härskarornas Gud, Israels Gud, så: Se, över Juda och över alla Jerusalems invånare skall jag låta all den olycka komma, som jag har förkunnat över dem, därför att de icke hörde, när jag talade till dem, och icke svarade, när jag kallade på dem.
Och till rekabiternas släkt sade Jeremia: Så säger HERREN Sebaot, Israels Gud: Därför att I haven hörsammat eder fader Jonadabs bud och hållit alla hans bud och i alla stycken gjort såsom han har bjudit eder,
därför säger HERREN Sebaot, Israels Gud, så: Aldrig skall den tid komma, då icke en avkomling av Jonadab, Rekabs son, står inför mitt ansikte.
I Jojakims, Josias sons, Juda konungs, fjärde regeringsår kom detta ord till Jeremia från HERREN; han sade:
Tag dig en bokrulle och teckna däri upp allt vad jag har talat till dig angående Israel och Juda och alla hednafolk, från den dag då jag först talade till dig i Josias tid ända till denna dag.
Kanhända skall Juda hus, när de höra all den olycka som jag har i sinnet att göra dem, vända om, var och en från sin onda väg, och så skall jag förlåta dem deras missgärning och synd.
Då kallade Jeremia till sig Baruk, Nerias son; och efter Jeremias diktamen tecknade Baruk i en bokrulle upp alla de ord som HERREN hade talat till honom.
Och Jeremia bjöd Baruk och sade: »Jag är själv under tvång, så att jag icke kan begiva mig till HERRENS hus.
Men gå du dit; och ur den rulle som du har skrivit efter min diktamen må du därpå fastedagen läsa UPP HERRENS ord inför folket i HERRENS hus.
Inför hela Juda, så många som komma in från sina städer, må du ock läsa upp dem.
Kanhända skola de då bönfalla inför HERREN och vända om, var och en från sin onda väg.
Ty stor är den vrede och förtörnelse som HERREN har uttalat över detta folk.»
Och Baruk, Nerias son, gjorde alldeles såsom profeten Jeremia hade bjudit honom: i HERRENS hus läste han ur boken upp HERRENS ord.
I Jojakims, Josias sons, Juda konungs, femte regeringsår, i nionde månaden, utlystes nämligen en fasta inför HERREN, vilken hölls av allt folket i Jerusalem och av allt det folk som från Juda städer hade kommit till Jerusalem.
Då läste Baruk ur boken upp Jeremias ord; han läste upp dem i HERRENS hus, i sekreteraren Gemarjas, Safans sons, kammare på den övre förgården, vid ingången till nya porten på HERRENS hus, inför allt folket.
När nu Mika; son till Gemarja, son till Safan, hade hört alla HERRENS ord uppläsas ur boken,
gick han ned till konungshuset och in i sekreterarens kammare; där sutto då alla furstarna: sekreteraren Elisama, Delaja, Semajas son, Elnatan, Akbors son, Gemarja, Safans son, Sidkia, Hananjas son, och alla de andra furstarna.
Och Mika omtalade för dem allt vad han hade hört Baruk läsa upp ur boken inför folket.
Då sände alla furstarna Jehudi, son till Netanja, son till Selemja, Kusis son, åstad till Baruk och läto säga honom: »Tag med dig den rulle varur du har läst inför folket, och kom hit.»
Och Baruk, Nerias son, tog rullen med sig och kom till dem.
Då sade de till honom: »Sätt dig ned och läs den inför oss.»
Och Baruk läste inför dem.
När de då hörde allt som stod där, sågo de med förskräckelse på varandra och sade till Baruk: »Vi måste omtala för konungen allt som står här.»
Och de frågade Baruk och sade: »Tala om för oss huru det skedde att du efter hans diktamen tecknade upp allt detta.»
Baruk svarade dem: »Han dikterade för mig allt detta, och jag tecknade upp det i boken med bläck.»
Då sade furstarna till Baruk: »Gå och göm dig, du jämte Jeremia, och låten ingen veta var I ären.»
Därefter, sedan de hade lämnat rullen i förvar i sekreteraren Elisamas kammare, gingo de in till konungen på förgården och omtalade så allt för konungen.
Då sände konungen Jehudi att hämta rullen; och denne hämtade den från sekreteraren Elisamas kammare.
Sedan läste Jehudi upp den inför konungen och inför alla furstarna, som stodo omkring konungen.
Konungen bodde då i vinterhuset, ty det var den nionde månaden.
Och kolpannan stod påtänd framför honom;
och så ofta Jehudi hade läst tre eller fyra spalter, skar han av rullen med pennkniven och kastade stycket på elden i kolpannan, ända till dess att hela rullen var förtärd av elden i kolpannan.
Och varken konungen själv eller någon av hans tjänare blev förskräckt eller rev sönder sina kläder, när de hörde allt detta som upplästes.
Och fastän Elnatan, Delaja och Gemarja bådo konungen att han icke skulle bränna upp rullen, lyssnade han icke till dem.
I stället bjöd konungen Jerameel, konungasonen, och Seraja, Asriels son, och Selemja, Abdeels son, att de skulle gripa skrivaren Baruk och profeten Jeremia.
Men HERREN gömde dem undan.
Men sedan konungen hade bränt upp rullen med det som Baruk efter Jeremias diktamen hade skrivit däri, kom HERRENS ord till Jeremia; han sade:
Tag dig nu åter en annan rulle och teckna däri upp allt vad som förut stod i den förra rullen, den som Jojakim, Juda konung, brände upp.
Men angående Jojakim, Juda konung, skall du säga: Så säger HERREN: Du har bränt upp denna rulle och sagt: »Huru kunde du skriva däri att konungen i Babel förvisso skall komma och fördärva detta land, och göra slut på både människor och djur däri?»
Därför säger HERREN så om Jojakim, Juda konung: Ingen ättling av honom skall sitta på Davids tron; och hans egen döda kropp skall komma att ligga utkastad, prisgiven åt hettan om dagen och åt kölden om natten.
Och jag skall hemsöka honom och hans avkomlingar och hans tjänare för deras missgärnings skull, och över dem och över Jerusalems invånare och över Juda män skall jag låta all den olycka komma, som jag har förkunnat över dem, fastän de icke hava velat höra.
Då tog Jeremia en annan rulle och gav den åt skrivaren Baruk, Nerias son; och efter Jeremias diktamen tecknade denne däri upp allt vad som hade stått i den bok som Jojakim, Juda konung, hade bränt upp i eld.
Och till detta lades ytterligare mycket annat av samma slag.
Och Sidkia, Josias son, blev konung i stället för Konja, Jojakims son; ty Nebukadressar, konungen i Babel, gjorde honom till konung i Juda land.
Men varken han eller hans tjänare eller folket i landet hörda på HERRENS ord, dem som han talade genom profeten Jeremia.
Dock sände konung Sidkia åstad Jehukal, Selemjas son, och prästen Sefanja, Maasejas son, till profeten Jeremia och lät säga: »Bed för oss till HERREN, vår Gud.»
Jeremia gick då ännu ut och in bland folket, ty man hade ännu icke satt honom i fängelse.
Och Faraos här hade då dragit ut från Egypten; och när kaldéerna, som belägrade Jerusalem, hade fått höra ryktet därom, hade de dragit sig tillbaka från Jerusalem.
Då kom HERRENS ord till profeten Jeremia; han sade:
Så säger HERREN, Israels Gud: Så skolen I svara Juda konung, som har sänt eder till mig för att fråga mig: »Se, Faraos här, som har dragit ut till eder hjälp, skall vända tillbaka till sitt land Egypten.
Sedan skola kaldéerna komma tillbaka och belägra denna stad och de skola då intaga den och bränna upp den i eld.
Därför säger HERREN så: Bedragen icke eder själva med att tänka: 'Kaldéerna skola nu en gång för alla draga bort ifrån oss'; ty de skola icke draga bort.
Nej, om I än så slogen kaldéernas hela här, när de strida mot eder, att allenast några svårt sårade män blevo kvar av dem, så skulle dessa resa sig upp, var och en i sitt tält, och skulle bränna upp denna stad i eld.
Men när kaldéernas här hade dragit sig tillbaka från Jerusalem för Faraos har,
ville Jeremia lämna Jerusalem och begiva sig till Benjamins land, för att där taga i besittning en jordlott bland folket.
När han då kom till Benjaminsporten, stod där såsom vakthavande en man vid namn Jiria, son till Selemja, son till Hananja; denne grep profeten Jeremia och sade: »Du vill gå över till kaldéerna.»
Jeremia svarade: »Det är icke sant; jag vill icke gå över till kaldéerna», men ingen hörde på honom.
Och Jiria grep Jeremia och förde honom till furstarna.
Och furstarna förtörnades på Jeremia och läto hudflänga honom och satte honom i häkte i sekreteraren Jonatans hus, ty detta hade de gjort till fängelse.
Men när Jeremia hade kommit i fängelsehålan, ned i fångvalven, och suttit där en lång tid,
sände konung Sidkia och lät hämta honom; och hemma hos sig frågade konungen honom hemligen och sade: »Har något ord kommit från HERREN Jeremia svarade: »Ja»; och han tillade: »Du skall bliva given i den babyloniske konungens hand.
Därefter frågade Jeremia konung Sidkia: »Varmed har jag försyndat mig mot dig och dina tjänare och detta folk, eftersom I haven satt mig i fängelse?
Och var äro nu edra profeter, som profeterade för eder och sade: 'Konungen i Babel skall icke komma över eder och över detta land'?
Så hör mig nu, herre konung; värdes upptaga min bön: sänd mig icke tillbaka till sekreteraren Jonatans hus, på det att jag icke må dö där.»
På konung Sidkias befallning satte man då Jeremia i förvar i fängelsegården, och gav honom en kaka bröd om dagen från Bagargatan, till dess att det var slut på allt brödet i staden.
Så stannade Jeremia i fängelsegården.
Men Sefatja, Mattans son, och Gedalja, Pashurs son, och Jukal, Selemjas son, och Pashur, Malkias son, hörde huru Jeremia talade till allt folket och sade:
»Så säger HERREN: Den som stannar kvar i denna stad, han skall dö genom svärd eller hunger eller pest, men den som giver sig åt kaldéerna, han skall få leva, ja, han skall vinna sitt liv såsom ett byte och få leva.
Ty så säger HERREN: Denna stad skall förvisso bliva given i händerna på den babyloniske konungens här, och han skall intaga den.
Då sade furstarna till konungen: »Denne man bör dödas, eftersom han gör folket modlöst, både det krigsfolk som ännu är kvar här i staden och jämväl allt det övrig: folket, i det att han talar sådan: ord till dem.
Ty denne man söker icke folkets välfärd, utan dess olycka.
Konung Sidkia svarade: »Välan han är i eder hand; ty konungen förmår intet mot eder.»
Då togo de Jeremia och kastad honom i konungasonen Malkias brunn på fängelsegården; de släppte Jeremia ditned med tåg.
I brunnen var intet vatten, men dy, och Jeremia sjönk ned i dyn.
När nu etiopiern Ebed-Melek, en hovman, som befann sig i konungshuset, under det att konungen uppehöll sig i Benjaminsporten, fick höra att de hade sänkt Jeremia ned i brunnen,
begav han sig åstad från konungshuset och talade till konungen och sade:
»Min herre konung, dessa män hava handlat illa i allt vad de hava gjort mot profeten Jeremia; ty de hava kastat honom i brunnen, där han strax måste dö av hunger, då nu intet bröd finnes i staden.
Då bjöd konungen etiopiern Ebed-Melek och sade: »Tag med dig härifrån trettio män, och drag profeten Jeremia upp ur brunnen, innan han dör.»
Så tog då Ebed-Melek männen med sig och begav sig till konungshuset, till rummet under skattkammaren, och hämtade därifrån trasor av sönderrivna och utslitna kläder och lät sänka ned dem med tåg till Jeremia i brunnen.
Och etiopiern Ebed-Melek sade till Jeremia: »Lägg trasorna av de sönderrivna och utslitna kläderna under dina armar, mellan dem och tågen.»
Och Jeremia gjorde så.
Sedan drogo de med tågen Jeremia upp ur brunnen.
Men Jeremia måste stanna i fängelsegården.
Därefter sände konung Sidkia åstad och lät hämta profeten Jeremia till sig vid tredje ingången till HERRENS hus.
Och konungen sade till Jeremia: »Jag vill fråga dig något dölj intet för mig.»
Jeremia sade till Sidkia: »Om jag säger dig något, så kommer du förvisso att låta döda mig; och om jag giver dig ett råd, så hör du icke på mig.»
Då gav konung Sidkia Jeremia sin ed, hemligen, och sade: »Så sant HERREN lever, han som har givit oss detta vårt liv: jag skall icke låta döda dig, ej heller skall jag lämna dig i händerna på dessa män som stå efter ditt liv.»
Då sade Jeremia till Sidkia: »Så säger HERREN, härskarornas Gud, Israels Gud: Om du giver dig åt den babyloniske konungens furstar, så skall du få leva, och denna stad skall då icke bliva uppbränd i eld, utan du och ditt hus skolen få leva.
Men om du icke giver dig åt den babyloniske konungens furstar, då skall denna stad bliva given i kaldéernas hand, och de skola bränna upp den i eld, och du själv skall icke undkomma deras hand.»
Konung Sidkia svarade Jeremia: »Jag rädes för de judar som hava gått över till kaldéerna; kanhända skall man lämna mig i deras händer, och de skola då hantera mig skändligt.»
Jeremia sade: »Man skall icke göra det.
Hör blott HERRENS röst i vad jag säger dig, så skall det gå dig väl, och du skall få leva.
Men om du vägrar att giva dig, så är detta vad HERREN har uppenbarat för mig:
Se, alla de kvinnor som äro kvar i Juda konungs hus skola då föras ut till den babyloniske konungens furstar; och kvinnorna skola klaga: 'Dina vänner sökte förleda dig, och de fingo makt med dig.
Dina fötter fastnade i dyn; då drogo de sig undan'
Och alla dina hustrur och dina barn skall man föra ut till kaldéerna, och du själv skall icke undkomma deras hand, utan skall varda gripen av den babyloniske konungens hand och bliva en orsak till att denna stad brännes upp i eld.»
Då sade Sidkia till Jeremia: »Låt ingen få veta vad här har blivit talat; eljest måste du dö.
Och om furstarna få höra att jag har talat med dig, och de komma till dig och säga till dig: 'Låt oss veta vad du har sagt till konungen; dölj intet för oss, så skola vi icke döda dig; säg oss ock vad konungen har sagt till dig' --
då skall du svara dem: 'Jag bönföll inför konungen att han icke skulle sända mig tillbaka till Jonatans hus för att dö där.'»
Och alla furstarna kommo till Jeremia och frågade honom; men han svarade dem alldeles såsom konungen hade bjudit honom.
Då tego de och gingo bort ifrån honom, eftersom ingen hade hört huru det verkligen hade gått till.
Men Jeremia fick stanna i fängelsegården ända till den dag då Jerusalem blev intaget.
-- efter det att Nebukadressar, konungen i Babel, med hela sin här hade kommit till Jerusalem och begynt belägra det i Sidkia, Juda konungs, nionde regeringsår, i tionde månaden,
och efter det att staden; hade blivit stormad i Sidkias elfte regeringsår, i fjärde månaden, på nionde dagen månaden
drogo alla den babyloniske konungens furstar därin och stannade i Mellersta porten: nämligen Nergal Sareser, Samgar-Nebo, Sarsekim, överste hovmannen, Nergal-Sareser, överste magern, och alla den babyloniske konungens övriga furstar.
Och när Sidkia, Juda konung, med allt sitt krigsfolk fick se dem, flydde de och drogo om natten ut ur staden, på den väg som ledde till den kungliga trädgården, genom porten mellan de båda murarna; och han tog vägen bort åt Hedmarken till.
Men kaldéernas här förföljde dem och de hunno upp Sidkia på Jeriko hedmarker.
Och de togo fatt honom och förde honom till Nebukadressar, den babyloniske konungen, i Ribla i Hamats land; där höll denne rannsakning och dom med honom.
Och den babyloniske konungen lät i Ribla slakta Sidkias barn inför hans ögon; också alla andra Juda ädlingar lät konungen i Babel slakta.
Och på Sidkia själv lät han sticka ut ögonen och lät fängsla honom med kopparfjättrar, för att föra honom till Babel.
Och kaldéerna brände upp i eld både konungens hus och folkets hus och bröto ned Jerusalems murar.
Och återstoden av folket, dem som voro kvar i staden, och de över löpare som hade gått över till honom, och vad som för övrigt var kvar av folket, dem förde Nebusaradan, översten för drabanterna, bort till Babel.
Men av de ringaste bland folket, av dem som ingenting hade, lämnade Nebusaradan, översten för drabanterna, några kvar i Juda land, och gav dem samtidigt vingårdar och åkerfält.
Och Nebukadressar, konungen Babel, gav genom Nebusaradan, översten för drabanterna, befallning angående Jeremia och sade:
»Tag honom och se i honom till godo, och gör honom icke något ont, utan gör med honom efter som han själv begär av dig.»
Då sände Nebusaradan, översten för drabanterna, och Nebusasban, överste hovmannen, och Nergal-Sareser, överste magern, och alla den babyloniske konungens övriga väldige --
dessa sände bort och läto hämta Jeremia ifrån fängelsegården och lämnade honom åt Gedalja, son till Ahikam, son till Safan, på det att denne skulle föra honom hem; så fick han stanna där bland folket.
Men HERRENS ord hade kommit till Jeremia, medan han var inspärrad i fängelsegården; han hade sagt:
Gå och säg till etiopiern Ebed-Melek: Så säger HERREN Sebaot, Israels Gud: Se, vad jag har förkunnat, det skall jag låta komma över denna stad, till dess olycka och icke till dess lycka, och det skall uppfyllas i din åsyn på den dagen.
Men dig skall jag rädda på den dagen, säger HERREN, och du skall icke bliva given i de mäns hand, som du fruktar för.
Ty jag skall förvisso låta dig komma undan, och du skall icke falla för svärd, utan vinna ditt liv såsom ett byte, därför att du har förtröstat på mig, säger HERREN.
Detta är det ord som kom till Jeremia från HERREN, sedan Nebusaradan, översten för drabanterna, hade släppt honom lös från Rama; denne lät nämligen hämta honom, där han låg bunden med kedjor bland alla andra fångar ifrån Jerusalem och Juda, som skulle föras bort till Babel.
Översten för drabanterna lät alltså hämta Jeremia och sade till honom: »HERREN, din Gud, hade förkunnat denna olycka över denna plats;
och HERREN har låtit den komma och har gjort såsom han hade sagt.
I haden ju syndat mot HERREN och icke hört hans röst, och därför har detta vederfarits eder.
Och se, nu löser jag dig i dag ur kedjorna som dina händer hava varit bundna med.
Om du är sinnad att komma med mig till Babel, så kom, och jag skall då se dig till godo; men om du icke är sinnad att komma med mig till Babel, så gör det icke.
Se, hela landet ligger öppet för dig; dit dig synes gott och rätt att gå, dit må du gå.»
Och då han ännu dröjde att vända tillbaka, tillade han: »Vänd tillbaka till Gedalja, son till Ahikam, son till Safan, som konungen i Babel har satt över Juda städer, och stanna hos honom bland folket.
Eller gå åt vilket annat håll som helst dit det behagar dig att gå.»
Och översten för drabanterna gav honom vägkost och skänker och lät honom gå.
Så begav sig då Jeremia till Gedalja, Ahikams son, i Mispa och stannade hos honom bland folket som var kvar i landet.
När då alla krigshövitsmännen på landsbygden jämte sina män fingo höra att konungen i Babel hade satt Gedalja, Ahikams son, över landet, och att han hade anförtrott åt honom män kvinnor och barn, och dem av de ringaste i landet, som man icke hade fört bort till Babel,
kommo de till Gedalja i Mispa, nämligen Ismael, Netanjas son, Johanan och Jonatan, Kareas söner, Seraja, Tanhumets son, netofatiten Ofais söner och Jesanja, maakatitens son, med sina män.
Och Gedalja, son till Ahikam, son till Safan, gav dem och deras män sin ed och sade: »Frukten icke för att tjäna kaldéerna.
Stannen kvar i landet, och tjänen konungen i Babel, så skall det gå eder väl.
Se, själv stannar jag kvar i Mispa, för att vara till tjänst åt kaldéer som komma till oss; men I mån insamla vin och frukt och olja och lägga det i edra kärl, och stanna kvar i de städer som I haven tagit i besittning.»
Då nu också alla de judar som voro i Moabs och Ammons barns och Edoms land, och de som voro i andra länder hörde att konungen i Babel hade låtit några av judarna bliva kvar, och att han hade satt över dem Gedalja, son till Ahikam, son till Safan,
vände alla dessa judar tillbaka från alla de orter dit de hade blivit fördrivna, och kommo till Juda land, till Gedalja i Mispa.
Och de inbärgade vin och frukt i stor myckenhet.
Men Johanan, Kareas son, och alla krigshövitsmännen på landsbygden kommo till Gedalja i Mispa
och sade till honom: »Du vet väl att Baalis, Ammons barns konung, har sänt hit Ismael, Netanjas son, för att slå ihjäl dig?»
Men Gedalja, Ahikams son, trodde dem icke.
Och Johanan, Kareas son, sade i hemlighet till Gedalja i Mispa: »Låt mig gå åstad och dräpa Ismael, Netanjas son; ingen skall få veta det.
Varför skulle han få slå ihjäl dig och så bliva en orsak till att vi judar, som hava församlats till dig, allasammans förskingras, och vad som är kvar av Juda förgås?»
Men Gedalja, Ahikams son, sade till Johanan, Kareas son: »Du får icke göra detta; ty vad du säger om Ismael är icke sant.»
Men i sjunde månaden kom Ismael, son till Netanja, son till Elisama, av konungslig börd och en av konungens väldige, med tio män till Gedalja, Ahikams son, i Mispa, och de höllo måltid tillsammans i Mispa.
Och Ismael, Netanjas son, jämte de tio män som voro med honom, överföll då Gedalja, son till Ahikam, son till Safan, och slog honom till döds med svärd, honom som konungen i Babel hade satt över landet.
Därjämte dräpte Ismael alla de judar som voro hos Gedalja i Mispa, så ock alla de kaldéer som funnos där, och som tillhörde krigsfolket.
Dagen efter den då han hade dödat Gedalja, och innan ännu någon visste av detta,
kom en skara av åttio män från Sikem, Silo och Samaria; de hade rakat av sig skägget och rivit sönder sina kläder och ristat märken på sig, och hade med sig spisoffer och rökelse till att frambära i HERRENS hus.
Och Ismael, Netanjas son, gick ut emot dem från Mispa, gråtande utan uppehåll.
Och när han mötte dem, sade han till dem: »Kommen in till Gedalja, Ahikams son.»
Men när de hade kommit in i staden, blevo de nedstuckna av Ismael, Netanjas son, och de män som voro med honom, och kastade i brunnen.
Men bland dem funnos tio män som sade till Ismael: »Döda oss icke; ty vi hava förråd av vete, korn, olja och honung gömda på landsbygden.»
Då lät han dem vara och dödade dem icke med de andra.
Och brunnen i vilken Ismael kastade kropparna av alla de män som han hade dräpt, när han dräpte Gedalja, var densamma som konung Asa hade låtit göra, när Baesa, Israels konung, anföll honom; denna fylldes nu av Ismael, Netanjas son, med ihjälslagna män.
Därefter bortförde Ismael såsom fångar allt det folk som var kvar i Mispa, konungadöttrarna och allt annat folk som hade lämnats kvar i Mispa, och som Nebusaradan, översten för drabanterna, hade anförtrott åt Gedalja, Ahikams son; dem bortförde Ismael, Netanjas son; såsom fångar och drog åstad bort till Ammons barn.
Men när Johanan, Kareas son, och alla de krigshövitsmän som voro med honom fingo höra om allt det onda som Ismael, Netanjas son, hade gjort,
togo de alla sina män och gingo åstad för att strida mot Ismael, Netanjas son; och de träffade på honom vid det stora vattnet i Gibeon.
Då nu hela skaran av dem som Ismael förde med sig fick se Johanan, Kareas son, och alla de krigshövitsmän som voro med honom, blevo de glada;
och de vände om, hela skaran av dem som Ismael hade bortfört såsom fångar ifrån Mispa, och gåvo sig åstad tillbaka till Johanan, Kareas son.
Men Ismael, Netanjas son, räddade sig med åtta män undan Johanan och begav sig till Ammons barn.
Och Johanan, Kareas son, och alla de krigshövitsmän som voro med honom togo med sig allt som var kvar av folket, dem av Mispas invånare, som han hade vunnit tillbaka från Ismael, Netanjas son, sedan denne hade dräpt Gedalja, Ahikams son: både krigsmän och kvinnor och barn och hovmän, som han hade hämtat tillbaka från Gibeon.
Och de drogo åstad; men i Kimhams härbärge invid Bet-Lehem stannade de, för att sedan draga vidare och komma till Egypten,
undan kaldéerna; ty de fruktade för dessa, eftersom Ismael, Netanjas son, hade dräpt Gedalja, Ahikams son, vilken konungen i Babel hade satt över landet
Då trädde alla krigshövitsmännen fram, jämte Johanan, Kareas son, och Jesanja, Hosajas son, så ock allt folket, både små och stora,
och sade till profeten Jeremia: »Värdes upptaga vår bön: bed för oss till HERREN, din Gud, för hela denna kvarleva -- ty vi äro blott några få, som hava blivit kvar av många; du ser med egna ögon att det är så med oss.
Må så HERREN, din Gud, kungöra för oss vilken väg vi böra gå, och vad vi hava att göra.»
Profeten Jeremia svarade dem: »Jag vill lyssna till eder.
Ja, jag vill bedja till HERREN, eder Gud, såsom I haven begärt.
Och vadhelst HERREN svarar eder skall jag förkunna för eder; intet skall jag undanhålla för eder.»
Då sade de till Jeremia: »HERREN vare ett sannfärdigt och osvikligt vittne mot oss, om vi icke i alla stycken göra efter det ord varmed HERREN, din Gud, sänder dig till oss.
Det må vara gott eller ont, så vilja vi höra HERRENS, vår Guds, röst, hans som vi sända dig till; på det att det må gå oss väl, när vi höra HERRENS, vår Guds, röst.»
Och tio dagar därefter kom HERRENS ord till Jeremia.
Då kallade han till sig Johanan, Kareas son, och alla de krigshövitsmän som voro med honom, och allt folket, både små och stora,
och sade till dem: Så säger HERREN, Israels Gud, han som I haven sänt mig till, för att jag skulle hos honom bönfalla för eder:
Om I stannen kvar i detta land, så skall jag uppbygga eder och ej mer slå eder ned; jag skall plantera eder och ej mer upprycka eder.
Ty jag ångrar det onda som jag har gjort eder.
Frukten icke mer för konungen i Babel, som I nu frukten för, frukten icke för honom, säger HERREN.
Ty jag är med eder och vill frälsa eder och rädda eder ur hans hand.
Jag vill låta eder finna barmhärtighet; ja, han skall bliva barmhärtig mot eder och låta eder vända tillbaka till edert land.
Men om I sägen: »Vi vilja icke stanna i detta land», om I alltså icke hören HERRENS, eder Guds, röst,
utan tänken: »Nej, vi vilja begiva oss till Egyptens land, där vi slippa att se krig och höra basunljud och hungra efter bröd, där vilja vi bo» --
välan, hören då HERRENS ord, I kvarblivna av Juda: Så säger HERREN Sebaot, Israels Gud: Om I verkligen ställen eder färd till Egypten och kommen dit, för att bo där såsom främlingar,
så skall svärdet, som I frukten för, hinna upp eder där i Egyptens land, och hungersnöden, som I rädens för, skall följa efter eder dit till Egypten, och där skolen I dö.
Ja, de människor som ställa sin färd till Egypten, för att bo där, skola alla dö genom svärd, hunger och pest, och ingen av dem skall slippa undan och kunna rädda sig från den olycka som jag skall låta komma över dem.
Ty så säger HERREN Sebaot, Israels Gud: Likasom min vrede och förtörnelse har utgjutit sig över Jerusalems invånare, så skall ock min förtörnelse utgjuta sig över eder, om I begiven eder till Egypten, och I skolen bliva ett exempel som man nämner, när man förbannar, och ett föremål för häpnad, bannande och smälek, och I skolen aldrig mer få se denna ort.
Ja, HERREN säger till eder, I kvarblivna av Juda: Begiven eder icke till Egypten.
Märken väl att jag i dag har varnat eder.
Ty I bedrogen eder själva, när I sänden mig till HERREN, eder Gud, och saden: »Bed för oss till HERREN, vår Gud; och vadhelst HERREN, vår Gud, säger, det må du förkunna för oss, så vilja vi göra det.»
Jag har nu i dag förkunnat det för eder.
Men I haven icke velat höra HERRENS, eder Guds, röst, i allt det varmed han har sänt mig till eder.
Så veten nu att I skolen dö genom svärd, hunger och pest, på den ort dit I åstunden att komma, för att bo där såsom främlingar.
Men när Jeremia hade talat till allt folket alla HERRENS, deras Guds, ord, med vilka HERREN, deras Gud, hade sänt honom till dem, allt som sagt är,
då svarade Asarja, Hosajas son, och Johanan, Kareas son, och alla de övriga fräcka männen -- dessa svarade Jeremia: »Det är icke sant vad du säger; HERREN, vår Gud, har icke sänt dig och låtit säga: 'I skolen icke begiva eder till Egypten, för att bo där såsom främlingar.'
Nej, det är Baruk, Nerias son, som uppeggar dig mot oss, på det att vi må bliva givna i kaldéernas hand, för att dessa skola döda oss eller föra oss bort till Babel.»
Och varken Johanan, Kareas son, eller någon av krigshövitsmännen eller någon av folket ville höra HERRENS röst och stanna kvar i Juda land.
I stället togo Johanan, Kareas son, och alla krigshövitsmännen med sig alla de kvarblivna av Juda, dem som från alla de folk till vilka de hade varit fördrivna hade kommit tillbaka, för att bo i Juda land,
både män, kvinnor och barn, där till konungadöttrarna och alla andra som Nebusaradan, översten för drabanterna, hade lämnat kvar hos Gedalja, son till Ahikam, son till Safan, jämväl profeten Jeremia och Baruk, Nerias son,
och begåvo sig till Egyptens land, ty de ville icke höra HERRENS röst.
Och de kommo så fram till Tapanhes.
Och HERRENS ord kom till Jeremia i Tapanhes; han sade:
Tag dig några stora stenar och mura in dem i murbruket, där tegelgolvet lägges, vid ingången till Faraos hus i Tapanhes; gör detta inför judiska mäns ögon
och säg till dem: Så säger HERREN Sebaot, Israels Gud: Se, jag skall sända åstad och hämta min tjänare Nebukadressar, konungen i Babel, och hans tron skall jag sätta upp ovanpå de stenar som jag har låtit mura in har, och han skall på dem breda ut sin tronmatta.
Ty han skall komma och slå Egyptens land och giva i pestens våld den som hör pesten till, i fångenskapens våld den som hör fångenskapen till, i svärdets våld den som hör svärdet till.
Och jag skall tända eld på Egyptens gudahus, och han skall bränna upp dem och föra gudarna bort.
Och han skall rensa Egyptens land från ohyra, likasom en herde rensar sin mantel; sedan skall han draga därifrån i god ro.
Och han skall slå sönder stoderna i Bet-Semes i Egyptens land, och Egyptens gudahus skall han bränna upp i eld.
Detta är det ord som kom till Jeremia angående alla de judar som bodde i Egyptens land, dem som bodde i Migdol, Tapanhes, Nof och Patros' land; han sade:
»Så säger HERREN Sebaot, Israels Gud: I haven sett all den olycka som jag har låtit komma över Jerusalem och över alla Juda städer -- Se, de äro nu ödelagda, och ingen bor i dem;
detta för den ondskas skull som de bedrevo till att förtörna mig, i det att de gingo bort och tände offereld och tjänade andra gudar, som varken I själva eller edra fäder haden känt.
Och titt och ofta sände jag till eder alla mina tjänare profeterna och lät säga: 'Bedriven icke denna styggelse, som jag hatar.'
Men de ville icke höra eller böja sitt öra därtill, så att de omvände sig från sin ondska och upphörde att tända offereld åt andra gudar.
Därför blev min förtörnelse och vrede utgjuten, och den brann i Juda städer och på Jerusalems gator, så att de blevo ödelagda och förödda, såsom de nu äro.
Och nu säger HERREN, härskarornas Gud, Israels Gud, så: Varför bereden I eder själva stor olycka?
I utroten ju ur Juda både man och kvinna, både barn och spenabarn bland eder, så att ingen kvarleva av eder kommer att återstå;
I förtörnen ju mig genom edra händers verk, i det att I tänden offereld åt andra gudar i Egyptens land, dit I haven kommit, för att bo där såsom främlingar.
Härav måste ske att I varden utrotade, och bliven ett exempel som man nämner, när man förbannar, och ett föremål för smälek bland alla jordens folk.
Haven I förgätit edra fäders onda gärningar och Juda konungars onda gärningar och deras hustrurs onda gärningar och edra egna onda gärningar och edra hustrurs onda gärningar, vad de gjorde i Juda land och på Jerusalems gator?
Ännu i dag äro de icke ödmjukade; de frukta intet och vandra icke efter min lag och mina stadgar, dem som jag förelade eder och edra fäder.
Därför säger HERREN Sebaot, Israels Gud, så: Se, jag skall vända mitt ansikte mot eder till eder olycka, till att utrota hela Juda.
Och jag skall gripa de kvarblivna av Juda, som hava ställt sin färd till Egyptens land, för att bo där såsom främlingar.
Och de skola allasammans förgås, i Egyptens land skola de falla; genom svärd och hunger skola de förgås, både små och stora, ja, genom svärd och hunger skola de dö.
Och de skola bliva ett exempel som man nämner, när man förbannar, och ett föremål för häpnad, bannande och smälek.
Och jag skall hemsöka dem som bo i Egyptens land, likasom jag hemsökte Jerusalem, med svärd, hunger och pest.
Och bland de kvarblivna av Juda, som hava kommit för att bo såsom främlingar där i Egyptens land, skall ingen kunna rädda sig och slippa undan, så att han kan vända tillbaka till Juda land, dit de dock åstunda att få vända tillbaka, för att bo där.
Nej, de skola icke få vända tillbaka dit, förutom några få som bliva räddade.»
Då svarade alla männen -- vilka väl visste att deras hustrur tände offereld åt andra gudar -- och alla kvinnorna, som stodo där i en stor hop, så ock allt folket som bodde i Egyptens land, i Patros, de svarade Jeremia och sade:
»I det som du har talat till oss i HERRENS namn vilja vi icke hörsamma dig,
utan vi vilja göra allt vad vår mun har lovat, nämligen tända offereld åt himmelens drottning och utgjuta drickoffer åt henne, såsom vi och våra fader, våra konungar och furstar gjorde i Juda städer och på Jerusalems gator.
Då hade vi bröd nog, och det gick oss väl, och vi sågo icke till någon olycka.
Men från den stund då vi upphörde att tända offereld åt himmelens drottning och utgjuta drickoffer åt henne hava vi lidit brist på allt, och förgåtts genom svärd och hunger.
Och när vi nu tända offereld åt himmelens drottning och utgjuta drickoffer åt henne, är det då utan våra mäns samtycke som vi åt henne göra offerkakor, vilka äro avbilder av henne, och som vi utgjuta drickoffer åt henne?»
Men Jeremia sade till allt folket, till männen och kvinnorna och allt folket, som hade givit honom detta svar, han sade:
»Förvisso har HERREN kommit ihåg och tänkt på huru I haven tänt offereld i Juda städer och på.
Jerusalems gator, både I själva och edra fäder, både edra konungar och furstar och folket i landet.
Och HERREN kunde icke längre hava fördrag med eder för edert onda väsendes skull, och för de styggelsers skull som I bedreven, utan edert land blev ödelagt och ett föremål för häpnad och förbannelse, så att ingen kunde bo där, såsom vi nu se.
Därför att I tänden offereld och syndaden mot HERREN och icke villen höra HERRENS röst eller vandra efter hans lag, efter hans stadgar och vittnesbörd, därför har denna olycka träffat eder, såsom vi nu se».
Och Jeremia sade ytterligare till allt folket och till alla kvinnorna: »Hören HERRENS ord, I alla av Juda, som ären i Egyptens land,
Så säger HERREN Sebaot, Israels Gud: I och edra hustrur haven med edra händer fullgjort vad I taladen med eder mun, när I saden: 'Förvisso vilja vi fullgöra de löften som vi gjorde, att tända offereld åt himmelens drottning och utgjuta drickoffer åt henne.'
Välan, I mån hålla edra löften och fullgöra edra löften;
men hören då också HERRENS ord, I alla av Juda, som bon i Egyptens land: Se, jag svär vid mitt stora namn, säger HERREN, att i hela Egyptens land mitt namn icke mer skall varda nämnt av någon judisk mans mun, så att han säger: 'Så sant Herren, HERREN lever.'
Ty se, jag skall vaka över dem, till deras olycka, och icke till deras lycka, och alla män av Juda, som äro i Egyptens land, skola förgås genom svärd och hunger, till dess att de hava fått en ände.
Och allenast några som undkomma svärdet skola få vända tillbaka från Egyptens land till Juda land, en ringa hop.
Och så skola alla kvarblivna av Juda, som hava kommit till Egyptens land, för att bo där såsom främlingar, få förnimma vilkens ord det är som bliver beståndande, mitt eller deras.
Och detta skall för eder vara tecknet till att jag skall hemsöka eder på denna ort, säger HERREN, och I skolen så förnimma att mina ord om eder förvisso skola bliva beståndande, eder till olycka:
Så säger HERREN: Se, jag skall giva Farao Hofra, konungen i Egypten i hans fienders hand och i de mäns hand, som stå efter hans liv, likasom jag har givit Sidkia, Juda konung, i Nebukadressars, den babyloniske konungens, hand, hans som var hans fiende, och som stod efter hans liv.»
Detta är det ord som profeten Jeremia talade till Baruk, Nerias son, när denne efter Jeremias diktamen tecknade upp dessa tal i en bok, under Jojakims, Josias sons, Juda konungs, fjärde regeringsår; han sade:
Så säger HERREN, Israels Gud, om dig, Baruk:
Du säger: »Ve mig, ty HERREN har lagt ny sorg till min förra plåga!
Jag är så trött av suckande och finner ingen ro.»
Men så skall du svara honom: Så säger HERREN: Se, vad jag har byggt upp, det måste jag riva ned, och vad jag har planterat, det måste jag rycka upp; och detta gäller hela jorden.
Och du begär stora ting för dig!
Begär icke något sådant; ty se, jag skall låta olycka komma över all kött, säger HERREN, men dig skall jag låta vinna ditt liv såsom ett byte, till vilken ort du än må gå.
Detta är vad som kom till profeten Jeremia såsom HERRENS ord om hednafolken.
Om Egypten, angående den egyptiske konungen Farao Nekos här, som stod invid floden Frat, vid Karkemis, och som blev slagen av Nebukadressar, konungen i Babel, i Jojakims, Josias sons, Juda konungs, fjärde regeringsår.
Reden till sköld och skärm, och rycken fram till strid.
Spännen för hästarna och bestigen springarna, och ställen upp eder, med hjälmarna på.
Gören spjuten blanka, ikläden eder pansaren.
Men varav kommer detta som jag nu ser?
De äro förfärade.
De vika tillbaka; deras hjältar bliva slagna.
De taga till flykten utan att vända sig om.
Skräck från alla sidor! säger HERREN.
Ej ens den snabbaste kan fly undan, ej ens hjälten kan rädda sig.
Norrut, invid floden Frat, där stappla de och falla.
Vem är denne som stiger upp såsom Nilfloden, denne vilkens vatten svalla såsom strömmar?
Det är Egypten som stiger upp såsom Nilfloden, och såsom strömmar svalla hans vatten.
Han säger: »Jag vill stiga upp och övertäcka landet; jag vill fördärva städerna och dem som bo därinne.»
Ja, dragen ditupp, I hästar; stormen fram, I vagnar.
Må hjältarna tåga fram, etiopier och putéer, rustade med sköldar, och ludéer, rustade med bågar, bågar som de spänna.
Ty detta är Herrens; HERREN Sebaots, dag, en hämndedag, då han skall hämnas på sina motståndare; nu skall svärdet frossa sig mätt och dricka sig rusigt av deras blod.
Ty ett slaktoffer vill Herren, HERREN Sebaot, anställa i nordlandet vid floden Frat.
Drag upp till Gilead och hämta balsam, du jungfru dotter Egypten.
Men förgäves skaffar du dig läkemedel i mängd; du kan icke bliva helad.
Folken få höra om din skam, och av dina klagorop bliver jorden full; ty den ene hjälten stapplar på den andre, och de falla båda tillsammans.
Detta är det ord som HERREN talade till profeten Jeremia om att Nebukadressar, konungen i Babel, skulle komma och slå Egyptens land:
Förkunnen i Egypten och kungören i Migdol, ja, kungören i Nof, så ock i Tapanhes, och sägen: »Träd fram och gör dig redo, ty svärdet frossar runt omkring dig.»
Varför äro dina väldige slagna till marken?
De kunde ej hålla stånd, ty HERREN stötte dem bort.
Han kom många att stappla, och så föllo de, den ene över den andre; de ropade: »Upp, låt oss vända tillbaka till vårt folk och till vårt fädernesland, undan det härjande svärdet.»
Ja, man ropar där: »Farao är förlorad, Egyptens konung!
Han har förfelat sin tid.»
Så sant jag lever, säger konungen, han vilkens namn är HERREN Sebaot, en skall komma, väldig såsom Tabor ibland bergen, såsom Karmel vid havet.
Så reden nu till åt eder, I dottern Egyptens inbyggare, vad man behöver, när man skall gå i landsflykt.
Ty Nof skall bliva en ödemark och varda uppbränt, så att ingen kan bo där.
En skön kviga är Egypten; men en broms kommer farande norrifrån.
Också de legoknektar hon har i sitt land, lika gödda kalvar, ja, också de vända då om och fly allasammans, de kunna icke hålla stånd.
Ty deras ofärds dag har kommit över dem, deras hemsökelses tid.
Tyst smyger hon undan såsom en krälande orm, ty med härsmakt draga de fram, och med yxor komma de över henne, såsom gällde det att hugga ved.
De fälla hennes skog, säger HERREN, ty ogenomtränglig är den; talrikare äro de än gräshoppor, ja, de kunna ej räknas.
På skam kommer dottern Egypten; hon bliver given i nordlandsfolkets hand.
Så säger HERREN Sebaot, Israels Gud: Se, jag skall hemsöka Amon från No, så ock Farao och Egypten med dess gudar och dess konungar, ja, både Farao och dem som förlita sig på honom.
Och jag skall giva dem i de mans hand, som stå efter deras liv, i Nebukadressars, den babyloniske konungens, och i hans tjänares hand.
Men därefter skall landet bliva bebott såsom i forna dagar, säger HERREN.
Så frukta då icke, du min tjänare Jakob, och var ej förfärad, du Israel; ty se, jag skall frälsa dig ur det avlägsna landet, och dina barn ur deras fångenskaps land.
Och Jakob skall få komma tillbaka och leva i ro och säkerhet, och ingen skall förskräcka honom.
Ja, frukta icke, du min tjänare Jakob, säger HERREN, ty jag är med dig.
Och jag skall göra ände på alla de folk till vilka jag har drivit dig bort; men på dig vill jag ej alldeles göra ände, jag vill blott tukta dig med måtta; ty alldeles ostraffad kan jag ju ej låta dig bliva.
Detta är vad som kom till profeten Jeremia såsom HERRENS ord om filistéerna, förrän Farao hade intagit Gasa.
Så säger HERREN: Se, vatten stiga upp norrifrån och växa till en översvämmande ström; de översvämma landet och allt vad däri är, städerna med dem som bo därinne.
Och människorna ropa, alla landets inbyggare jämra sig
När bullret höres av hans hingstars hovslag, när hans vagnar dåna, när hans hjuldon rassla, då se ej fäderna sig om efter barnen, så maktlösa stå de
inför den dag som kommer med fördärv över alla filistéer, med undergång för alla dem som äro kvar till att försvara Tyrus och Sidon.
Ty HERREN skall fördärva filistéerna, kvarlevan från Kaftors ö.
Skallighet stundar för Gasa, det är förbi med Askelon, med kvarlevan i deras dalbygd.
Huru länge skall du rista märken på dig?
Ack ve!
Du HERRENS svärd, när skall du äntligen få ro, Drag dig tillbaka i din skida, vila dig och var stilla.
Dock, huru skulle det kunna få ro, då det är HERRENS bud det utför?
Mot Askelon, mot Kustlandet vid havet, mot dem har han bestämt det.
Om Moab.
Så säger HERREN Sebaot, Israels Gud: Ve över Nebo, ty det är förstört!
Kirjataim har kommit på skam och är intaget, fästet har kommit på skam och ligger krossat.
Moabs berömmelse är icke mer.
I Hesbon förehar man onda anslag mot det: »Upp, låt oss utrota det, så att det icke mer är ett folk.»
Också du, Madmen, skall förgöras, svärdet skall följa dig i spåren.
Klagorop höras från Horonaim, förödelse och stort brak.
Ja, Moab ligger förstört; högljutt klaga dess barn.
Uppför Halluhots höjd stiger man under gråt, och på vägen ned till Horonaim höras ångestfulla klagorop över förstörelsen.
Flyn, rädden edra liv, och bliven som torra buskar i öknen.
Ty därför att du förlitar dig på dina verk och dina skatter, skall ock du bliva intagen; och Kemos skall gå bort i fångenskap och hans präster och furstar med honom.
Och en förhärjare skall komma över var stad, så att ingen stad skall kunna rädda sig; dalen skall bliva förstörd och slätten ödelagd, såsom HERREN har sagt.
Given vingar åt Moab, ty flygande måste han fly bort.
Hans städer skola bliva mark, och ingen skall bo i dem.
Förbannad vare den som försumligt utför HERRENS verk, förbannad vare den som dröjer att bloda sitt svärd.
I säkerhet har Moab levat från sin ungdom och har legat i ro på sin drägg; han har icke varit tömd ur ett kärl i ett annat, icke vandrat bort i fångenskap; därför har hans smak behållit sig, och hans lukt har ej förvandlats.
Se, därför skola dagar komma, säger HERREN, då jag skall sända till honom vintappare, som skola tappa honom och tömma hans kärl och krossa hans krukor.