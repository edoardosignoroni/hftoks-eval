Sedan träffade de på fältet en egyptisk man; honom togo de med sig till David.
Och när de hade givit honom bröd att äta och vatten att dricka
och när de ytterligare hade givit honom ett stycke fikonkaka och två russinkakor att äta, kom livskraften tillbaka i honom igen.
På tre dygn hade han nämligen varken ätit eller druckit.
Och David frågade honom: »Vem tillhör du, och varifrån är du?»
Han svarade: »Jag är en egyptisk yngling, tjänare åt en amalekitisk man; men min herre övergav mig för tre dagar sedan, därför att jag blev sjuk.
Vi hade nämligen infallit i den del av Sydlandet, som tillhör keretéerna, och i det område som tillhör Juda, och i den del av Sydlandet, som tillhör Kaleb, och vi hade bränt upp Siklag i eld.»
David sade till honom: »Vill du föra mig ned till den rövarskaran?»
Han svarade: »Lova mig med ed vid Gud att du icke dödar mig eller utlämnar mig åt min herre, så vill jag föra dig ned till den rövarskaran.»
Så förde han honom ditned, och de lågo då kringspridda överallt på marken och åto och drucko och förlustade sig med allt det stora byte som de hade tagit ur filistéernas land och ur Juda land.
Och ända från skymningen intill nästa dags afton höll David på med att nedgöra dem; och ingen enda av dem kom undan, utom fyra hundra tjänare som satte sig upp på kamelerna och flydde.
Och David räddade allt vad amalekiterna hade tagit; sina båda hustrur räddade David också.
Ingen saknades, varken liten eller stor, ingens son och ingens dotter, ej heller något av bytet eller något av det som de hade tagit med sig; David förde alltsammans tillbaka.
David tog ock alla får och fäkreatur, och man drev dessa framför den övriga boskapen och ropade: »Detta är Davids byte.»
Och när David kom tillbaka till de två hundra man som hade varit för trötta att följa honom, och som därför hade fått stanna kvar vid bäcken Besor, gingo dessa åstad för att möta David och det folk som han hade med sig; då gick David fram till folket och hälsade dem.
Men allahanda onda och illasinnade män, bland dem som hade följt med David, togo till orda och sade: »Eftersom dessa icke följde med oss, skola vi icke giva dem något av bytet som vi hava räddat; var och en av dem må allenast taga sin hustru och sina barn med sig och gå hem.»
Men David svarade: »Så skolen I icke göra, mina bröder, med det som HERREN har givit oss, då han bevarade oss och gav i vår hand denna rövarskara, som kom över oss.
Och vem skulle för övrigt härutinnan vilja lyssna till eder?
Nej, sådan deras lott är, som draga med i striden, sådan skall deras lott vara, som stanna vid trossen; de skola dela jämnt med varandra.»
Och därvid blev det, från den dagen och allt framgent; ty han gjorde detta till lag och rätt i Israel, såsom det är ännu i dag.
När sedan David kom till Siklag, sände han en del av bytet till de äldste i Juda, sina vänner, i det han lät säga: »Detta är en skänk till eder av bytet från HERRENS fiender.»
Han sände till de äldste i Betel, de äldste i Ramot i Sydlandet och de äldste i Jattir;
till de äldste i Aroer, de äldste i Sifamot och de äldste i Estemoa;
till de äldste i Rakal, de äldste i jerameeliternas städer och de äldste i kainéernas städer;
till de äldste i Horma, de äldste i Bor-Asan och de äldste i Atak;
till de äldste i Hebron och till alla de orter där David hade vandrat omkring med sina män.
Och filistéerna stridde mot Israel; och Israels män flydde för filistéerna och föllo slagna på berget Gilboa.
Och filistéerna ansatte ivrigt Saul och hans söner.
Och filistéerna dödade Jonatan, Abinadab och Malki-Sua, Sauls söner.
När då Saul själv blev häftigt anfallen och bågskyttarna kommo över honom, greps han av stor förskräckelse för skyttarna.
Och Saul sade till sin vapendragare: »Drag ut ditt svärd och genomborra mig därmed, så att icke dessa oomskurna komma och genomborra mig och hantera mig skändligt.»
Men hans vapendragare ville det icke, ty han fruktade storligen.
Då tog Saul själv svärdet och störtade sig därpå.
Men när vapendragaren såg att Saul var död, störtade han sig ock på sitt svärd och följde honom i döden.
Så dogo då med varandra på den dagen Saul och hans tre söner och hans vapendragare, och därjämte alla hans män.
Och när israeliterna på andra sidan dalen och på andra sidan Jordan förnummo att Israels män hade flytt, och att Saul och hans söner voro döda, övergåvo de städerna och flydde; sedan kommo filistéerna och bosatte sig i dem.
Dagen därefter kommo filistéerna för att plundra de slagna och funno då Saul och hans tre söner, där de lågo fallna på berget Gilboa.
Då höggo de av hans huvud och drogo av honom hans vapen och sände dem omkring i filistéernas land och läto förkunna det glada budskapet i sitt avgudahus och bland folket.
Och de lade hans vapen i Astartetemplet, men hans kropp hängde de upp på Bet-Sans mur.
Men när invånarna i Jabes i Gilead hörde vad filistéerna hade gjort med Saul,
stodo de upp, alla stridbara män, och gingo hela natten och togo Sauls och hans söners kroppar ned från Bet-Sans mur, och begåvo sig därefter till Jabes och förbrände dem där.
Sedan togo de deras ben och begrovo dem under tamarisken i Jabes och fastade så i sju dagar.
Efter Sauls död, när David hade kommit tillbaka från segern över Amalek, och när David sedan i två dagar hade uppehållit sig i Siklag,
då hände sig på tredje dagen att en man kom från Sauls läger, med sönderrivna kläder och med jord på sitt huvud.
Och när han kom in till David, föll han ned till jorden och bugade sig.
David frågade honom: »Varifrån kommer du?»
Han svarade honom: »Jag kommer såsom flykting ifrån Israels läger.»
Då sade David till honom: »Huru har det gått?
Säg mig det.»
Han svarade: »Folket har flytt ur striden, många av folket hava också fallit och dött; Saul och hans son Jonatan äro ock döda.»
David frågade den unge mannen som berättade detta för honom: »Huru vet du att Saul och hans son Jonatan äro döda?»
Den unge mannen som hade framfört underrättelsen till honom svarade: »Jag kom av en händelse upp på berget Gilboa, och där fick jag se Saul stödja sig mot sitt spjut, under det att vagnar och ryttare ansatte honom.
När han då vände sig om och fick se mig, ropade han på mig, och jag svarade: 'Här är jag.'
Då frågade han mig vem jag var, och jag svarade honom att jag var en amalekit.
Sedan sade han till mig: 'Träd fram hit till mig och giv mig dödsstöten, ty jag är gripen av dödens vanmakt, om ock livet ännu alltjämt är kvar i mig.'
Då trädde jag fram till honom och dödade honom, ty jag visste ju att han icke skulle kunna överleva sitt fall.
Och jag tog diademet som satt på hans huvud, och ett armband som satt på hans arm, och jag bar nu detta hit till min herre.»
Då fattade David i sina kläder och rev sönder dem; så gjorde ock alla de män som voro där med honom.
Och de höllo dödsklagan och gräto och fastade ända till aftonen för Sauls och hans son Jonatans skull, och för HERRENS folks och för Israels hus' skull, därför att de hade fallit för svärd.
Och David frågade den unge mannen som hade framfört underrättelsen till honom: »Varifrån är du?»
Han svarade: »Jag är son till en amalekit som lever här såsom främling.»
David sade till honom: »Kände du då ingen fruktan för att uträcka din hand till att förgöra HERRENS smorde?»
Och David kallade på en av sina män och sade: »Kom hit och stöt ned honom.»
Och han slog honom till döds.
Och David sade till honom: »Ditt blod komme över ditt huvud, ty din egen mun har vittnat mot dig, i det att du sade: 'Jag har dödat HERRENS smorde.'»
Och David sjöng följande klagosång över Saul och hans son Jonatan,
och han befallde att man skulle lära Juda barn »Bågsången»; den är upptecknad i »Den redliges bok»:
»Din härlighet, Israel, ligger slagen på dina höjder.
Huru hava icke hjältarna fallit!
Förkunnen det icke i Gat, bebåden det ej på Askelons gator, för att filistéernas döttrar icke må glädja sig, de oomskurnas döttrar ej fröjda sig.
I Gilboa berg, på eder må ej falla dagg eller regn, ej ses offergärdsskördar.
Ty hjältarnas sköld blev där till smälek, Sauls sköld, ej sedan smord med olja.
Från slagnas blod, från hjältars hull vek Jonatans båge icke tillbaka, vände Sauls svärd ej omättat åter.
Saul och Jonatan, så kära och ljuvliga för varandra i livet, de blevo ej heller skilda i döden, de två, som voro snabbare än örnar, starka mer än lejon.
Israels döttrar, gråten över Saul, över honom som klädde eder i scharlakan och praktskrud och prydde edra kläder med gyllene smycken.
Huru hava icke hjältarna fallit i striden!
Jonatan ligger slagen på dina höjder.
Jag sörjer över dig, du min broder Jonatan; mycket ljuvlig var du mig.
Dyrbar var mig din kärlek, mer än kvinnokärlek.
Huru hava icke hjältarna fallit, de båda stridssvärden förgåtts!»
Därefter frågade David HERREN: »Skall jag draga upp till någon av Juda städer?»
HERREN svarade honom: »Drag upp.»
Då frågade David: »Vart skall jag draga upp?», Han svarade: »Till Hebron.»
Så drog då David ditupp jämte sina båda hustrur, Ahinoam från Jisreel och Abigail, karmeliten Nabals hustru.
David lät ock sina män draga ditupp, var och en med sitt husfolk; och de bosatte sig i Hebrons städer.
Dit kommo nu Juda män och smorde David till konung över Juda hus.
När man berättade för David att det var männen i Jabes i Gilead som hade begravit Saul,
skickade David sändebud till männen i Jabes i Gilead och lät säga till dem: »Varen välsignade av HERREN, därför att I haven bevisat eder herre Saul den barmhärtighetstjänsten att begrava honom!
Så må nu ock HERREN bevisa barmhärtighet och trofasthet mot eder.
Själv vill jag också göra eder gott, därför att I haven gjort detta.
Varen alltså nu vid gott mod och oförskräckta, fastän eder herre Saul är död; det är nu jag som av Juda hus har blivit smord till konung över dem.»
Men Abner, Ners son, Sauls härhövitsman, tog Sauls son Is-Boset och förde honom över till Mahanaim
och gjorde honom till konung i Gilead och asuréernas land och Jisreel, så ock över Efraim, Benjamin och hela det övriga Israel.
Sauls son Is-Boset var fyrtio år gammal, när han blev konung över Israel, och han regerade i två år.
Allenast Juda hus höll sig till David.
Den tid David var konung i Hebron över Juda hus utgjorde sammanräknat sju år och sex månader.
Och Abner, Ners son, drog ut med Sauls son Is-Bosets folk ifrån Mahanaim till Gibeon.
Joab, Serujas son, och Davids folk drogo också ut; och de mötte varandra vid Gibeons damm.
Där stannade de på var sin sida om dammen.
Och Abner sade till Joab: »Må vi låta några unga män stå upp och utföra en krigslek i vår åsyn.»
Joab svarade: »Må så ske.»
Då stodo de upp och gingo fram i lika antal: tolv för Benjamin och för Sauls son Is-Boset, och tolv av Davids folk.
Och de fattade varandra i huvudet och stötte svärdet i sidan på varandra och föllo så allasammans därför blev detta ställe kallat Helkat-Hassurim vid Gibeon.
Sedan begynte en mycket hård strid på den dagen; men Abner och Israels män blevo slagna av Davids folk.
Nu funnos där tre söner till Seruja: Joab, Abisai och Asael.
Och Asael var snabbfotad såsom en gasell på fältet.
Och Asael förföljde Abner, utan att vika undan vare sig till höger eller till vänster från Abner.
Då vände Abner sig om och sade: »Är det du, Asael?»
Han svarade: »Ja.»
Då sade Abner till honom: »Vänd dig åt annat håll, åt höger eller åt vänster.
Angrip någon av de yngre och försök att taga hans rustning.»
Men Asael ville icke låta honom vara.
Då sade Abner ännu en gång till Asael: »Låt mig vara.
Du vill väl icke att jag skall slå dig till jorden?
Huru skulle jag sedan kunna se din broder Joab i ansiktet?»
När han ändå icke ville låta honom vara, gav Abner honom med bakändan av sitt spjut en stöt i underlivet, så att spjutet gick ut baktill; och han föll ned där och dog på stället.
Och var och en som kom till platsen där Asael hade fallit ned och dött stannade där.
Och Joab och Abisai förföljde Abner.
Men när solen hade gått ned och de hade kommit till Ammahöjden, som ligger gent emot Gia, åt Gibeons öken till,
då samlade sig Benjamins barn tillhopa bakom Abner, så att de utgjorde en sluten skara, och intogo en ställning på toppen av en och samma höjd.
Och Abner ropade till Joab och sade: »Skall då svärdet få oavlåtligen frossa?
Förstår du icke att detta måste leda till ett bittert slut?»
Huru länge tänker du dröja, innan du befaller ditt folk att upphöra med att förfölja sina bröder?»
Joab svarade: »Så sant Gud lever: om du ingenting hade sagt, då hade folket först i morgon fått draga sig tillbaka och upphöra att förfölja sina bröder.»
Därefter lät Joab stöta i basunen; då stannade allt folket och förföljde icke mer Israel.
Och sedan stridde de icke vidare.
Men Abner och hans män tågade genom Hedmarken hela den natten; därefter gingo de över Jordan och tågade vidare hela förmiddagen och kommo så till Mahanaim.
Joab åter samlade tillhopa allt folket, sedan han hade upphört att förfölja Abner; då fattades av Davids folk nitton man utom Asael.
Davids folk hade däremot slagit till döds tre hundra sextio man av Benjamin och av Abners folk.
Och de togo upp Asael och begrovo honom i hans faders grav i Bet-Lehem.
Därefter tågade Joab och hans män hela natten och kommo i dagningen till Hebron.
Kriget mellan Sauls hus och Davids hus blev långvarigt.
Därunder blev David allt starkare och starkare, men Sauls hus allt svagare och svagare.
I Hebron föddes söner åt David. hans förstfödde var Amnon, som han fick med Ahinoam från Jisreel.
Hans andre son var Kilab, som han fick med Abigal, karmeliten Nabals hustru, och den tredje var Absalom, son till Maaka, som var dotter till Talmai, konungen i Gesur.
Den fjärde var Adonia, Haggits son, och den femte var Sefatja, Abitals son.
Den sjätte var Jitream, som David fick med sin hustru Egla.
Dessa föddes åt David i Hebron.
Så länge kriget varade mellan Sauls hus och Davids hus, bistod Abner kraftigt Sauls hus.
Men Saul hade haft en bihustru vid namn Rispa, Ajas dotter; och Is-Boset sade till Abner: »Varför har du gått in till min faders bihustru?»
För dessa hans ord blev Abner mycket vred och sade: »Är jag då ett hundhuvud från Juda land?
Just då jag bevisar barmhärtighet mot din fader Sauls hus, mot hans bröder och hans vänner, och icke har låtit dig falla i Davids hand, just då tillvitar du mig att hava begått en missgärning med denna kvinna.
Gud straffe Abner nu och framgent, om jag icke hädanefter handlar så mot David som HERREN med ed har lovat honom:
jag vill göra så, att konungadömet tages ifrån Sauls hus, och att i stället Davids tron bliver upprest över både Israel och Juda, från Dan ända till Beer-Seba.»
Då tordes han icke säga ett ord mer åt Abner, av fruktan för honom.
Men Abner skickade strax sändebud till David och lät säga: »Vem tillhör landet?», och lät vidare säga: »Slut förbund med mig, så skall jag bistå dig och göra så, att hela Israel går över till dig.»
Han svarade: »Gott!
Jag vill sluta förbund med dig.
Men en sak fordrar jag av dig, nämligen att du icke träder fram inför mitt ansikte utan att hit medföra Mikal, Sauls dotter, när du kommer för att träda fram inför mitt ansikte.»
Därefter skickade David sändebud till Is-Boset, Sauls son, och lät säga: »Giv mig åter min hustru Mikal, som jag förvärvade mig för ett hundra filistéers förhudar.»
Då sände Is-Boset åstad och lät taga henne ifrån hennes man, Paltiel, Lais' son.
Men hennes man gick med henne och följde henne under beständig gråt ända till Bahurim.
Här sade Abner till honom: »Vänd om och gå dina färde.»
Då vände han om.
Och Abner hade underhandlat med de äldste i Israel och sagt: »Sedan lång tid tillbaka haven I sökt att få David till konung över eder.
Fullborden nu edert uppsåt, ty så har HERREN sagt om David: Genom min tjänare Davids hand skall jag frälsa mitt folk Israel ifrån filistéernas hand och ifrån alla dess fienders hand.»
Likaledes talade Abner härom med benjaminiterna.
Därefter gick Abner ock åstad for att tala med David i Hebron om allt vad Israel och hela Benjamins hus hade funnit lämpligt att svara.
När då Abner, åtföljd av tjugu man, kom till David i Hebron, gjorde David ett gästabud för Abner och hans män.
Och Abner sade till David: »Jag vill stå upp och gå åstad och församla hela Israel till min herre konungen, för att de må sluta förbund med dig, så att du bliver konung på vad villkor dig lyster.»
Sedan lät David Abner gå, och han drog bort i frid.
Just då kommo Davids folk och Joab hem från ett strövtåg och förde med sig ett stort byte; men Abner var nu icke längre kvar hos David i Hebron, ty denne hade låtit honom gå, och han hade dragit bort i frid.
Men när Joab och hela hans här kom hem, berättade man för honom och sade: »Abner, Ners son, kom till konungen, och denne lät honom gå, och han drog bort i frid.»
Då gick Joab in till konungen och sade: »Vad har du gjort!
Då nu Abner hade kommit till dig, varför lät du då honom gå, så att han fritt kunde draga sina färde?
Du känner väl Abner, Ners son?
Han kom hit för att bedraga dig.
Han ville utforska ditt görande och låtande, och utforska allt vad du förehar.
Sedan, när Joab hade gått ut från David, sände han bud efter Abner, och sändebuden förde denne tillbaka från Bor-Hassira.
Men David visste intet därom.
När Abner så hade kommit tillbaka till Hebron, förde Joab honom avsides till mitten av porten, under förevändning att tala enskilt med honom; där sårade han honom till döds med en stöt i underlivet -- detta for att hämnas sin broder Asaels blod.
När David sedan fick höra detta, sade han: »Jag och mitt konungadöme äro oskyldiga inför HERREN evinnerligen till Abners, Ners sons blod.
Må det komma över Joabs huvud och över hela hans faders hus; och må i Joabs hus aldrig fattas män som hava flytning, eller som äro spetälska, eller som stödja sig på krycka, eller som falla för svärd, eller som lida brist på bröd.»
Så hade nu Joab och hans broder Abisai dräpt Abner, därför att denne hade dödat deras broder Asael vid Gibeon, under striden.
Och David sade till Joab och allt folket som var med honom: »Riven sönder edra kläder och höljen eder i sorgdräkt och hållen dödsklagan efter Abner.»
Och konung David gick själv bakom båren.
Så begrovo; de Abner i Hebron; och konungen brast ut i gråt vid Abners grav, och allt folket grät.
Och konungen sjöng följande klagosång över Abner: »Måste då Abner dö en gudlös dåres död?
Dina händer voro ju ej bundna, dina fötter ej slagna i fjättrar.
Du föll såsom man faller för ogärningsmän.»
Då begrät allt folket honom ännu mer.»
Och allt folket kom för att förmå David att äta något under dagens lopp; men David betygade med ed och sade: »Gud straffe mig nu och framgent, om jag smakar bröd eller något annat, förrän solen har gått ned.»
När folket hörde detta, behagade det dem alla väl, likasom allt annat som konungen gjorde behagade allt folket väl.
Och allt folket och hela Israel insåg då att konungen ingen del hade haft i att Abner, Ners son, hade blivit dödad.
Och konungen sade till sina tjänare: »I veten nogsamt att en furste och en stor man i dag har fallit i Israel.
Men jag är ännu svag, fastän jag är smord till konung, och dessa män, Serujas söner, äro starkare än jag.
HERREN vedergälle den som ont gör, efter hans ondska.»
Då nu Sauls son hörde att Abner var död i Hebron, sjönk allt hans mod, och hela Israel var förskräckt.
Men Sauls son hade till hövitsmän för sina strövskaror två män, av vilka den ene hette Baana och den andre Rekab, söner till Rimmon från Beerot, av Benjamins barn.
Ty också Beerot räknas till Benjamin;
men beerotiterna flydde till Gittaim och bodde där sedan såsom främlingar, vilket de göra ännu i dag.
(Också Jonatan, Sauls son, hade lämnat efter sig en son, som nu var ofärdig i fötterna.
Han var nämligen fem år gammal, när budskapet om Saul och Jonatan kom från Jisreel, och då tog hans sköterska honom och flydde; men under hennes bråda flykt föll han omkull och blev därefter halt; och han hette Mefiboset.)
Nu gingo beerotiten Rimmons söner Rekab och Baana åstad och kommo till Is-Bosets hus, då det var som hetast på dagen, medan han låg i sin middagssömn.
När de så, under förevändning att hämta vete, hade kommit in i det inre av huset, sårade de honom med en stöt i underlivet; därefter flydde Rekab och hans broder Baana undan.
De kommo alltså in i huset, när han låg på sin vilobädd i sovkammaren, och sårade honom till döds och höggo huvudet av honom; därpå togo de hans huvud och färdades genom Hedmarken hela natten.
Och de förde så Is-Bosets huvud till David i Hebron och sade till konungen: »Se här är Is-Bosets, Sauls sons, din fiendes, huvud, hans som stod efter ditt liv.
HERREN har i dag givit min herre konungen hämnd på Saul och hans efterkommande.»
Då svarade David Rekab och hans broder Baana, beerotiten Rimmons söner, och sade till dem: »Så sant HERREN lever, han som har förlossat mig från all nöd:
den som förkunnade för mig och sade: 'Nu är Saul död', och som menade sig vara en glädjebudbärare, honom lät jag gripa och dräpa i Siklag, honom som jag eljest skulle hava givit budbärarlön;
huru mycket mer skall jag icke då nu, när ogudaktiga män hava dräpt en oskyldig man i hans eget hus, på hans säng, utkräva hans blod av eder hand och utrota eder från jorden!»
På Davids befallning dräpte hans män dem sedan och höggo av deras händer och fötter och hängde upp dem vid dammen i Hebron.
Men Is-Bosets huvud togo de, och de begrovo det i Abners grav i Hebron.
Sedan; kommo alla Israels stammar till David i Hebron och sade så: »Vi äro ju ditt kött och ben.
Redan för länge sedan, då Saul ännu var konung över oss, var det du som var ledare och anförare för Israel.
Och till dig har HERREN sagt: Du skall vara en herde för mitt folk Israel, ja, du skall vara en furste över Israel.»
När så alla de äldste i Israel kommo till konungen i Hebron, slöt konung David ett förbund med dem där i Hebron, inför HERREN; och sedan smorde de David till konung över Israel.
David var trettio år gammal, när han blev konung, och han regerade i fyrtio år.
I Hebron regerade han över Juda i sju år och sex månader, och i Jerusalem regerade han i trettiotre år över hela Israel och Juda.
Och konungen drog med sina män till Jerusalem, mot jebuséerna, som bodde där i landet.
De sade då till David: »Hitin kommer du icke; blinda och halta skola driva dig bort, de mena att David icke skall komma hitin.»
Men David intog likväl Sions borg, det är Davids stad.
Och David sade på den dagen: »Vemhelst som slår ihjäl en jebusé och tränger fram till vattenledningen, han slår ihjäl just dessa halta och blinda, som David hatar.»
Därför plägar man säga: »Ingen blind och halt må komma in i huset.»
Sedan tog David sin boning på borgen och kallade den Davids stad.
Där uppförde David byggnader runt omkring, från Millo och vidare inåt.
Och David blev allt mäktigare och mäktigare, och HERREN, härskarornas Gud, var med honom.
Och Hiram, konungen i Tyrus, skickade sändebud till David med cederträ, därjämte ock timmermän och stenhuggare; och de byggde ett hus åt David.
Och David märkte att HERREN hade befäst honom såsom konung över Israel, och att han hade upphöjt hans konungadöme, för sitt folk Israels skull.
Och David tog sig ännu flera bihustrur och hustrur från Jerusalem, sedan han hade kommit från Hebron; och åt David föddes ännu flera söner och döttrar.
Dessa äro namnen på de söner som föddes åt honom i Jerusalem: Sammua, Sobab, Natan, Salomo,
Jibhar, Elisua, Nefeg, Jafia,
Elisama, Eljada och Elifelet.
Men när filistéerna hörde att David hade blivit smord till konung över Israel, drogo de allasammans upp för att fånga David.
När David hörde detta, drog han ned till borgen.
Och sedan filistéerna hade kommit fram, spridde de sig i Refaimsdalen.
Då frågade David HERREN: »Skall jag draga upp mot filistéerna?
Vill du då giva dem i min hand?»
HERREN svarade David: »Drag upp; ty jag skall giva filistéerna i din hand.
Och David kom till Baal-Perasim, och där slog David dem.
Då sade han: »HERREN har brutit ned mina fiender inför mig, likasom en vattenflod bryter ned.»
Därav fick det stället namnet Baal-Perasim.
De lämnade där efter sig sina avgudabilder, och David och hans män togo dessa med sig.
Men filistéerna drogo upp ännu en gång och spridde sig i Refaimsdalen.
När David då frågade HERREN, svarade han: »Du skall icke draga ditupp; du må kringgå dem bakifrån, så att du kommer över dem från det håll där bakaträden stå.
Så snart du sedan hör ljudet av steg i bakaträdens toppar, skynda då raskt fram, ty då har HERREN dragit ut framför dig till att slå filistéernas här.»
David gjorde såsom HERREN hade bjudit honom; och han slog filistéerna och förföljde dem från Geba ända fram emot Geser.
Åter församlade David allt utvalt manskap i Israel, trettio tusen man.
Och David bröt upp och drog åstad med allt sitt folk ifrån Baale-Juda, för att därifrån föra upp Guds ark, som hade fått sitt namn efter HERREN Sebaot, honom som tronar på keruberna.
Och de satte Guds ark på en ny vagn och förde den bort ifrån Abinadabs hus på höjden; och Ussa och Ajo, Abinadabs söner, körde den nya vagnen.
Så förde de Guds ark bort ifrån Abinadabs hus på höjden, och följde själva med, och Ajo gick därvid framför arken.
Och David och hela Israels hus fröjdade sig inför HERREN, med allahanda instrumenter av cypressträ, med harpor, psaltare, pukor, skallror och cymbaler.
Men när de kommo till Nakonslogen, räckte Ussa ut sin hand mot Guds ark och fattade i den, ty oxarna snavade.
Då upptändes HERRENS vrede mot Ussa, och Gud slog honom där för hans förseelse, så att han föll ned död där vid Guds ark.
Men det gick David hårt till sinne att HERREN så hade brutit ned Ussa; och han kallade det ställe Peres-Ussa, såsom det heter ännu i dag.
Och David betogs av sådan fruktan för HERREN på den dagen, att han sade: »Huru skulle jag töras låta HERRENS ark komma till mig?»
Därför ville David icke låta flytta in HERRENS ark till sig i David stad, utan lät sätta in den i gatiten Obed-Edoms hus.
Sedan blev HERRES ark kvar i gatiten Obed-Edoms hus i tre månader; men HERREN välsignade Obed-Edom och hela hans hus.
När det nu blev berättat för konung David att HERREN hade välsignat Obed-Edoms hus och allt vad han hade, för Guds arks skull, då gick David åstad och hämtade Guds ark ur Obed-Edoms hus upp till Davids stad under jubel.
Och när de som buro HERRENS ark hade gått sex steg framåt, offrade han en tjur och en gödkalv.
Själv dansade David med all makt inför HERREN, och därvid var David iklädd en linne-efod.
Så hämtade David och hela Israel HERRENS ark ditupp under jubel och basuners ljud.
När då HERRENS ark kom in i Davids stad, blickade Mikal, Sauls dotter, ut genom fönstret, och när hon såg konung David hoppa och dansa inför HERREN fick hon förakt för honom i sitt hjärta.
Sedan de hade fört HERRENS ark ditin, ställde de den på dess plats i tältet som David hade slagit upp åt den; och därefter offrade David brännoffer inför HERREN, så ock tackoffer.
När David hade offrat brännoffret och tackoffret välsignade han folket i HERREN Sebaots namn.
Och åt allt folket, åt var och en i hela hopen av israeliter, både man och kvinna, gav han en kaka bröd, ett stycke kött och en druvkaka.
Sedan gick allt folket hem, var och en till sitt.
Men när David kom tillbaka för att hälsa sitt husfolk, gick Mikal, Sauls dotter, ut emot honom och sade: »Huru härlig har icke Israels konung visat sig i dag, då han i dag har blottat sig för sina tjänares tjänstekvinnors ögon, såsom löst folk plägar göra!»
Då sade David till Mikal: »Inför HERREN, som har utvalt mig framför din fader och hela hans hus, och som har förordnat mig till furste över HERRENS folk, över Israel -- inför HERREN fröjdade jag mig.
Dock kände jag mig rätteligen för ringa till detta, ja, jag var i mina ögon allt för låg därtill.
Skulle jag då söka ära hos tjänstekvinnorna, om vilka du talade?»
Och Mikal, Sauls dotter, fick inga barn, så länge hon levde.
Då nu konungen satt i sitt hus, sedan HERREN hade låtit honom få ro runt omkring för alla hans fiender,
sade han till profeten Natan: »Se, jag bor i ett hus av cederträ, under det att Guds ark bor i ett tält.
Natan sade till konungen: »Välan, gör allt vad du har i sinnet; ty HERREN är med dig.»
Men om natten kom HERRENS ord till Natan; han sade:
»Gå och säg till min tjänare David: Så säger HERREN: Skulle du bygga mig ett hus att bo i?
Jag har ju icke bott i något hus, allt ifrån den dag då jag förde Israels barn upp ur Egypten ända till denna dag, utan jag har flyttat omkring i ett tält, i ett tabernakel.
Har jag då någonsin, varhelst jag flyttade omkring med alla Israels barn, talat och sagt så till någon enda av Israels stammar, som jag har förordnat till herde för mitt folk Israel: 'Varför haven I icke byggt mig ett hus av cederträ?'
Och nu skall du säga så till min tjänare David: Så säger HERREN Sebaot: Från betesmarken, där du följde fåren, har jag hämtat dig, för att du skulle bliva en furste över mitt folk Israel.
Och jag har varit med dig på alla dina vägar och utrotat alla dina fiender för dig.
Och jag vill göra dig ett namn, så stort som de störstes namn på jorden.
Jag skall bereda en plats åt mitt folk Israel och plantera det, så att det får bo kvar där, utan att vidare bliva oroat.
Orättfärdiga människor skola icke mer förtrycka det, såsom fordom skedde,
och såsom det har varit allt ifrån den tid då jag förordnade domare över mitt folk Israel; och jag skall låta dig få ro för alla dina fiender.
Så förkunnar nu HERREN för dig att HERREN skall uppbygga ett hus åt dig.
När din tid är ute och du vilar hos dina fäder, skall jag efter dig upphöja den son som skall utgå ur ditt liv; och jag skall befästa hans konungadöme.
Han skall bygga ett hus åt mitt namn, och jag skall befästa hans konungatron för evig tid.
Jag skall vara hans fader, och han skall vara min son, så att jag visserligen, om han gör något illa, skall straffa honom med ris, såsom människor pläga tuktas, och med plågor, sådana som hemsöka människors barn;
men min nåd skall icke vika ifrån honom, såsom jag lät den vika ifrån Saul, vilken jag lät vika undan för dig.
Ditt hus och ditt konungadöme skola bliva beståndande inför dig till evig tid; ja, din tron skall vara befäst för evig tid.»
Alldeles i överensstämmelse med dessa ord och med denna syn talade nu Natan till David.
Då gick konung David in och satte sig ned inför HERRENS ansikte och sade: »Vem är jag, Herre, HERRE, och vad är mitt hus, eftersom du har låtit mig komma härtill?
Och detta har ändå synts dig vara för litet, Herre, HERRE; du har ock talat angående din tjänares hus om det som ligger långt fram i tiden. och härom har du talat på människosätt, Herre, HERRE!
Vad skall nu David vidare tala till dig?
Du känner ju din tjänare, Herre, HERRE.
För ditt ords skull och efter ditt hjärta har du gjort allt detta stora och förkunnat det för din tjänare.
Därför är du ock stor HERRE Gud, ty ingen är dig lik, och ingen Gud finnes utom dig, efter allt vad vi hava hört med våra öron.
Och var finnes på jorden något enda folk likt ditt folk Israel, något folk som en Gud själv har gått åstad att förlossa åt sig till ett folk, för att så göra sig ett namn -- ja, för att göra dessa stora ting med eder och dessa fruktansvärda gärningar med ditt land, inför ditt folk, det som du förlossade åt dig från Egypten, från hedningarna och deras gudar.
Och du har berett åt dig ditt folk Israel, dig till ett folk för evig tid, och du, HERRE, har blivit deras Gud.
Så uppfyll nu, HERRE Gud, för evig tid vad du har talat om din tjänare och om hans hus; gör såsom du har talat.
Då skall ditt namn bliva stort till evig tid, så att man skall säga: 'HERREN Sebaot är Gud över Israel.'
Och så skall din tjänare Davids hus bestå inför dig.
Ty du, HERRE Sebaot, Israels Gud, har uppenbarat för din tjänare och sagt: 'Jag vill bygga dig ett hus.'
Därför har din tjänare fått frimodighet att bedja till dig denna bön.
Och nu, Herre, HERRE, du är Gud, och dina ord äro sanning; och du du har lovat din tjänare detta goda,
så värdes nu välsigna din tjänares hus, så att det förbliver evinnerligen inför dig.
Ja, du, Herre, HERRE, har lovat det, och genom din välsignelse skall din tjänares hus bliva välsignat evinnerligen.»
En tid härefter slog David filistéerna och kuvade dem.
Därvid bemäktigade sig David huvudstaden och tog den ur filistéernas hand.
Han slog ock moabiterna och mätte dem med snöre, i det att han lät dem lägga sig ned på jorden: med två snörlängder mätte han ut den del av dem, som skulle dödas, och med en full snörlängd den del som han låt leva.
Så blevo moabiterna David underdåniga och förde till honom skänker.
Likaledes slog David Hadadeser, Rehobs son, konungen i Soba, när denne hade dragit åstad för att utsträcka sitt välde till floden.
Och David tog till fånga av han folk ett tusen sju hundra ryttare och tjugu tusen man fotfolk; och David lät avskära fotsenorna på alla vagnshästarna, utom på ett hundra hästar, som han skonade.
När sedan araméerna från Damaskus kommo för att hjälpa Hadadeser, konungen i Soba, nedgjorde David tjugutvå tusen man av dem.
Och David insatte fogdar bland araméerna i Damaskus, och araméerna blevo David underdåniga och förde till honom skänker.
Så gav HERREN seger åt David, varhelst han drog fram.
Och David tog de gyllene sköldar som Hadadesers tjänare hade burit och förde dem till Jerusalem.
Och från Hadadesers städer Beta och Berotai tog konung David koppar i stor myckenhet.
Då nu Toi, konungen i Hamat, hörde att David hade slagit Hadadesers hela här,
sände han sin son Joram till konung David för att hälsa honom och lyckönska honom, därför att han hade givit sig i strid med Hadadeser och slagit honom; ty Hadadeser hade varit Tois fiende.
Och han hade med sig kärl av silver, av guld och av koppar.
Också dessa helgade konung David åt HERREN, likasom han hade gjort med det silver och guld han hade tagit från alla de folk som han hade underlagt sig:
från araméerna, moabiterna, Ammons barn, filistéerna och amalekiterna, så ock med det byte han hade tagit från Hadadeser, Rehobs son, konungen i Soba.
Och när David kom tillbaka från sin seger över araméerna, gjorde han sig ytterligare ett namn i Saltdalen, där han slog aderton tusen man.
Och han insatte fogdar i Edom, i hela Edom insatte han fogdar; och alla edoméer blevo David underdåniga.
Så gav HERREN seger åt David, varhelst han drog fram.
David regerade nu över hela Israel; och David skipade lag och rätt åt allt sitt folk.
Joab, Serujas son, hade befälet över krigshären, och Josafat Ahiluds son, var kansler.
Sadok, Ahitubs son, och Ahimelek, Ebjatars son, voro präster, och Seraja var sekreterare.
Benaja, Jojadas son, hade befälet över keretéerna och peletéerna; dessutom voro Davids söner präster.
Och David sade: »Finnes ännu någon kvar av Sauls hus, mot vilken jag kan bevisa barmhärtighet för Jonatans skull?»
Nu hade Sauls hus haft en tjänare vid namn Siba; honom hämtade man till David.
Då sade konungen till honom: »Är du Siba?»
Han svarade: »Ja, din tjänare.»
Konungen frågade: »Finnes ingen kvar av Sauls hus, mot vilken jag kan bevisa barmhärtighet, såsom Gud är barmhärtig?»
Siba svarade konungen: »Ännu finnes kvar en son till Jonatan, en som är ofärdig i fötterna.»
Konungen frågade honom »Var är han?»
Siba svarade konungen: »Han är nu i Makirs, Ammiels sons, hus i Lo-Debar.»
Då sände konung David och lät hämta honom från Makirs, Ammiels sons, hus i Lo-Debar.
När så Mefiboset, Sauls son Jonatans son, kom in till David, föll han ned på sitt ansikte och bugade sig.
Då sade David: »Mefiboset!»
Han svarade: »Ja, din tjänare hör.»
David sade till honom: »Frukta icke, ty jag vill bevisa barmhärtighet mot dig för din fader Jonatans skull, och jag vill giva dig allt din faders Sauls jordagods tillbaka, och du skall äta vid mitt bord beständigt.»
Då bugade han sig och sade: »Vad är jag, din tjänare, eftersom du vänder dig till en sådan död hund som jag är?»
Därefter tillkallade konungen Siba, Sauls tjänare, och sade till honom; »Allt som Saul och hela hans hus har ägt giver jag åt din herres son.
Och du med dina söner och dina tjänare skall bruka jorden åt honom och inbärga skörden, för att din herres son må hava bröd att äta, dock skall Mefiboset, din herres son, beständigt äta vid mitt bord.»
Siba hade nämligen femton söner och tjugu tjänare.
Då sade Siba till konungen: »Din tjänare skall i alla stycken göra såsom min herre konungen bjuder sin tjänare.» »Ja», svarade han, »Mefiboset skall äta vid mitt bord, såsom vore han en av konungens söner.»
Mefiboset hade en liten son, som hette Mika.
Och alla som bodde i Sibas hus blevo Mefibosets tjänare.
Själv bodde Mefiboset i Jerusalem, eftersom han beständigt skulle äta vid konungens bord.
Och han var halt på båda fötterna.
En tid härefter dog Ammons barns konung, och hans son Hanun blev konung efter honom.
Då sade David: »Jag vill bevisa Hanun, Nahas' son, vänskap, likasom hans fader bevisade mig vänskap.»
Och David sände några av sina tjänare för att trösta honom i hans sorg efter fadern.
När så Davids tjänare kommo till Ammons barns land,
sade Ammons barns furstar till sin herre Hanun: »Menar du att David därmed att han sänder tröstare till dig vill visa dig att han ärar din fader?
Nej, för att undersöka staden, för att bespeja och sedan fördärva den har David sänt sina tjänare till dig.»
Då tog Hanun Davids tjänare och lät raka av dem halva skägget och skära av deras kläder mitt på, ända uppe vid sätet, och lät dem så gå.
När man berättade detta för David, sände han bud emot dem; ty männen voro ju mycket vanärade.
Och konungen lät säga: »Stannen i Jeriko, till dess edert skägg hinner växa ut, och kommen så tillbaka.»
Då nu Ammons barn insågo att de hade gjort sig förhatliga för David, sände de bort och lejde från Aram-Bet-Rehob och Aram-Soba tjugu tusen man fotfolk, av konungen i Maaka ett tusen man och av Tobs män tolv tusen.
När David hörde detta, sände han åstad Joab med hela hären, de tappraste krigarna.
Och Ammons barn drogo ut och ställde upp sig till strid framför stadsporten; men de från Aram-Soba och Rehob, ävensom Tobs män och maakatéerna, ställde upp sig för sig själva på fältet.
Då Joab nu såg att han hade fiender både framför sig och bakom sig, gjorde han ett urval bland allt Israels utvalda manskap och ställde sedan upp sig mot araméerna.
Men det övriga folket överlämnade han åt sin broder Absai, vilken med dem ställde upp sig mot Ammons barn.
Och han sade: »Om araméerna bliva mig övermäktiga, så skall du komma mig till hjälp; och om Ammons barn bliva dig övermäktiga, så vill jag tåga till din hjälp.
Var nu vid gott mod; ja, låt oss visa mod i striden för vårt folk och för vår Guds städer.
Sedan må HERREN göra vad honom täckes.»
Därefter ryckte Joab fram med sitt folk till strid mot araméerna och de flydde för honom.
Men när Ammons barn sågo att araméerna flydde, flydde också de för Abisai och begåvo sig in i staden.
Då drog Joab bort ifrån Ammons barn och begav sig tillbaka till Jerusalem.
Då alltså araméerna sågo att de hade blivit slagna av Israel, församlade de sig allasammans.
Och Hadadeser sände bud att de araméer som bodde på andra sidan floden skulle rycka ut; dessa kommo då till Helam, anförda av Sobak, Hadadesers härhövitsman.
När detta blev berättat för David, församlade han hela Israel och gick över Jordan och kom till Helam; och araméerna ställde upp sig i slagordning mot David och gåvo sig i strid med honom.
Men araméerna flydde för Israel, och David dräpte av araméerna manskapet på sju hundra vagnar, så ock fyrtio tusen ryttare; deras härhövitsman Sobak slog han ock där till döds.
Då alltså Hadadesers alla lydkonungar sågo att de hade blivit slagna av israeliterna, ingingo de fred med dem och blevo dem underdåniga.
Efter detta fruktade araméerna för att vidare hjälpa Ammons barn.
Följande år, vid den tid då konungarna plägade draga i fält, sände David åstad Joab och med honom sina tjänare och hela Israel; och de härjade Ammons barns land och belägrade Rabba, medan David stannade kvar i Jerusalem.
Då hände sig en afton, när David hade stått upp från sitt läger och gick omkring på konungshusets tak, att han från taket fick se en kvinna som badade; och kvinnan var mycket fager att skåda.
David sände då åstad och förfrågade sig om kvinnan, och man sade: »Det är Bat-Seba, Eliams dotter, hetiten Urias hustru.»
Då sände David några män med uppdrag att hämta henne, och hon kom till honom, och han låg hos henne, när hon hade helgat sig från sin orenhet.
Sedan återvände hon hem.
Men kvinnan blev havande; hon sände då åstad och lät underrätta David därom och säga: »Jag är havande.»
Då sände David till Joab detta bud: »Sänd till mig hetiten Uria.»
Så sände då Joab Uria till David.
Och när Uria kom till David, frågade denne om det stod väl till med Joab och med folket, och huru kriget gick.
Därefter sade David till Uria: »Gå nu ned till ditt hus och två dina fötter.»
När då Uria gick ut ur konungens hus, sändes en gåva från konungen efter honom.
Men Uria lade sig till vila vid ingången till konungshuset, jämte hans herres alla andra tjänare, och gick icke ned till sitt eget hus.
Detta berättade man för David och sade: »Uria har icke gått ned till sitt hus.»
Då sade David till Uria: »Du kommer ju från resan; varför har du då icke gått ned till ditt hus?»
Uria svarade David: »Arken och Israel och Juda bo nu i lägerhyddor, och min herre Joab och min herres tjänare äro lägrade ute på marken: skulle jag då gå in i mitt hus för att äta och dricka och ligga hos min hustru?
Så sant du lever, så sant din själ lever: jag vill icke göra så.»
Då sade David till Uria: »Stanna här också i dag, så vill jag i morgon sända dig åstad.»
Så stannade då Uria i Jerusalem den dagen och den följande.
Och David inbjöd honom till sig och lät honom äta och dricka med sig och gjorde honom drucken.
Men om aftonen gick han ut och lade sig på sitt läger tillsammans med sin herres tjänare, och gick icke ned till sitt hus.
Följande morgon skrev David ett brev till Joab och sände det med Uria.
I brevet skrev han så: »Ställen Uria längst fram, där striden är som häftigast, och dragen eder sedan tillbaka från honom, så att han bliver slagen till döds.»
Under belägringen av staden skickade då Joab Uria till den plats där han visste att de tappraste männen funnos.
Och männen i staden gjorde ett utfall och gåvo sig i strid med Joab, och flera av folket, av Davids tjänare, föllo; också hetiten Uria dödades.
Då sände Joab och lät berätta för David allt vad som hade hänt under striden.
Och han bjöd budbäraren och sade: »När du har omtalat för konungen allt vad som har hänt under striden,
då upptändes kanske konungens vrede, och han säger till dig: 'Varför gingen I under striden så nära intill staden?
Vissten I icke att de skulle skjuta uppifrån muren?
Vem var det som slog ihjäl Abimelek, Jerubbesets son?
Var det icke en kvinna som kastade en kvarnsten ned på honom från muren, så att han dödades, där i Tebes?
Varför gingen I då så nära intill muren?'
Men då skall du säga: 'Din tjänare Uria, hetiten, är ock död.'»
Budbäraren gick åstad och kom och berättade för David allt vad Joab hade sänt honom att säga;
budbäraren sade till David: »Männen blevo oss övermäktiga och drogo ut mot oss på fältet, men vi slogo dem tillbaka ända till stadsporten.
Då sköto skyttarna uppifrån muren på dina tjänare, så att flera av konungens tjänare dödades; din tjänare Uria, hetiten, är ock död.»
Då sade David till budbäraren: »Så skall du säga till Joab: 'Låt icke detta förtryta dig, ty svärdet förtär än den ene, än den andre; fortsatt med kraft stadens belägring och förstör den.'
Och intala honom så mod.»
Då nu Urias hustru hörde att hennes man Uria var död, höll hon dödsklagan efter sin man.
Och när sorgetiden var förbi, sände David och lät hämta henne hem till sig, och hon blev hans hustru; därefter födde hon honom en son.
Men vad David hade gjort misshagade HERREN.
Och HERREN sände Natan till David.
När han kom in till honom, sade han till honom: »Två män bodde i samma stad; den ene var rik och den andre fattig.
Den rike hade får och fäkreatur i stor myckenhet.
Men den fattige hade icke mer än ett enda litet lamm, som han hade köpt; han uppfödde det, och det växte upp hos honom och hans söner, tillsammans med dem: det åt av hans brödstycke och drack ur hans bägare och låg i hans famn och var för honom såsom en dotter.
Så kom en vägfarande till den rike mannen; då nändes han icke taga av sina får och fäkreatur för att tillreda åt den resande som hade kommit till honom, utan han tog den fattige mannens lamm och tillredde det åt mannen som hade kommit till honom.»
Då upptändes Davids vrede storligen mot den mannen, och han sade till Natan: »Så sant HERREN lever: dödens barn är den man som har gjort detta.
Och lammet skall han ersätta fyradubbelt, därför att han gjorde sådant, och eftersom han var så obarmhärtig.»
Men Natan sade till David: »Du är den mannen.
Så säger HERREN, Israels Gud: Jag har smort dig till konung över Israel, och jag har räddat dig ur Sauls hand.
Jag har givit dig din herres hus och lagt din herres hustrur i din famn; ja jag har givit dig Israels hus och Juda.
Och om detta skulle vara för litet, så vore jag villig att ytterligare giva dig både ett och annat.
Varför har du då föraktat HERRENS ord och gjort vad ont är i hans ögon?
Hetiten Uria har du låtit slå ihjäl med svärd, och hans hustru har du tagit till hustru åt dig själv; ja, honom har du dräpt med Ammons barns svärd.
Så skall nu icke heller svärdet vika ifrån ditt hus till evig tid, därför att du har föraktat mig och tagit hetiten Urias hustru till hustru åt dig.
Så säger HERREN: Se, jag skall låta olyckor komma över dig från ditt eget hus, och jag skall taga dina hustrur inför dina ögon och giva dem åt en annan, och han skall ligga hos dina hustrur mitt på ljusa dagen.
Ty väl har du gjort sådant i hemlighet, men jag vill låta detta ske inför hela Israel, och det på ljusa dagen.»
Då sade David till Natan: »Jag har syndat mot HERREN.»
Natan sade till David: »Så har ock HERREN tillgivit dig din synd; du skall icke dö.
Men eftersom du genom denna gärning har kommit HERRENS fiender att förakta honom, skall ock den son som har blivit född åt dig döden dö.»
Sedan gick Natan hem igen.
Och HERREN slog barnet som Urias hustru hade fött åt David, han slog det, så att det blev dödssjukt.
Då sökte David Gud för gossens skull; och David höll fasta, och när han kom hem, låg han på bara marken över natten.
Då stodo de äldste i hans hus upp och gingo till honom, för att förmå honom att stiga upp från marken; men han ville icke, och han åt icke heller något med dem.
Men på sjunde dagen dog barnet.
Då fruktade Davids tjänare att om tala för honom att barnet hade dött, ty de tänkte: »När vi talade till honom, medan barnet ännu levde, ville han ju icke lyssna till våra ord.
Huru skulle vi då kunna säga till honom att barnet har dött?
Han kunde göra något ont.»
Men när David såg att hans tjänare viskade med varandra, förstod han att barnet hade dött.
Då frågade David sina tjänare: »Har barnet dött?»
De svarade: »Ja.»
Då stod David upp från marken och tvådde sig och smorde sig och bytte om kläder och gick in i HERRENS hus och tillbad.
Och när han kom hem igen, begärde han att man skulle sätta fram mat åt honom, och han åt.
Då sade hans tjänare till honom: »Varför gör du på detta sätt?
Medan barnet levde, fastade du och grät för dess skull; men så snart barnet har dött, står du upp och äter!»
Han svarade: så länge barnet ännu levde, fastade och grät jag, ty jag tänkte: 'Vem vet, kanhända bliver HERREN mig nådig och låter barnet få leva.'
Men nu, när det har dött, varför skulle jag då fasta?
Kan jag väl skaffa honom tillbaka igen?
Jag går bort till honom, men han kommer icke tillbaka till mig.»
Och David tröstade sin hustru Bat-Seba och gick in till henne och låg hos henne.
Och hon födde en son, åt vilken han gav namnet Salomo.
Och HERREN älskade honom
och sände ett budskap med profeten Natan, och denne gav honom namnet Jedidja, för HERRENS skull.
Och Joab angrep Rabba i Ammons barns land och intog konungastaden.
Sedan sände Joab bud till David och lät säga honom: »Jag har angripit Rabba och har redan intagit Vattenstaden.
Så församla du nu det övriga folket och belägra staden och intag den, så att det icke bliver jag som intager staden och får bära namnet därför.»
Då församlade David allt folket och tågade till Rabba och angrep det och intog det.
Och han tog deras konungs krona från hans huvud; den vägde en talent guld och var prydd med en dyrbar sten.
Den sattes nu på Davids huvud.
Och han förde ut byte från staden i stor myckenhet.
Och folket därinne förde han ut och lade dem under sågar och tröskvagnar av järn och bilor av järn och överlämnade dem åt Molok.
Så gjorde han mot Ammons barns alla städer.
Sedan vände David med allt folket tillbaka till Jerusalem.
Därefter tilldrog sig följande Davids son Absalom hade en skön syster som hette Tamar, och Davids son Amnon fattade kärlek till henne.
Ja, Amnon kom för sin syster Tamars skull i en sådan vånda att han blev sjuk; ty hon var jungfru, och det syntes Amnon icke vara möjligt att göra henne något.
Men Amnon hade en vän, som hette Jonadab, en son till Davids broder Simea; och Jonadab var en mycket klok man.
Denne sade nu till honom: »Varför ser du var morgon så avtärd ut, du konungens son?
Vill du icke säga mig det?»
Amnon svarade honom: »Jag har fattat kärlek till min broder Absaloms syster Tamar.»
Jonadab sade till honom: »Lägg dig på din säng och gör dig sjuk.
När då din fader kommer för att besöka dig, så säg till honom: 'Låt min syster Tamar komma och giva mig något att äta, men låt henne tillreda maten inför mina ögon; så att jag ser det och kan få den ur hennes hand att äta.'»
Då lade Amnon sig och gjorde sig sjuk.
När nu konungen kom för att besöka honom, sade Amnon till konungen: »Låt min syster Tamar komma hit och tillaga två kakor inför mina ögon, så att jag kan få dem ur hennes hand att äta.»
Då sände David bud in i huset till Tamar och lät säga: »Gå till din broder Amnons hus och red till åt honom något att äta.»
Tamar gick då åstad till sin broder Amnons hus, där denne låg till sängs.
Och hon tog deg och knådade den och gjorde därav kakor inför hans ögon och gräddade kakorna.
Därefter tog hon pannan och lade upp dem därur inför hans ögon; men han ville icke äta.
Och Amnon sade: »Låt alla gå ut härifrån.
Då gingo alla ut därifrån.
Sedan sade Amnon till Tamar: »Bär maten hitin i kammaren, så att jag får den ur din hand att äta.»
Då tog Tamar kakorna som hon hade tillrett och bar dem in i kammaren till sin broder Amnon.
Men när hon kom fram med dem till honom, för att han skulle äta, fattade han i henne och sade till henne: »Kom hit och ligg hos mig, min syster.»
Hon sade till honom: »Ack nej, min broder, kränk mig icke; ty sådant får icke ske i Israel.
Gör icke en sådan galenskap.
Vart skulle jag då taga vägen med min skam?
Och du själv skulle ju sedan i Israel hållas för en dåre.
Tala nu med konungen; han vägrar nog icke att giva mig åt dig.»
Men han ville icke lyssna till hennes ord och blev henne övermäktig och kränkte henne och låg hos henne.
Men därefter fick Amnon en mycket stor motvilja mot henne; ja, den motvilja han fick mot henne var större än den kärlek han hade haft till henne.
Och Amnon sade till henne: »Stå upp och gå din väg.»
Då sade hon till honom: »Gör dig icke skyldig till ett så svårt brott som att driva bort mig; det vore värre än det andra som du har gjort med mig.»
Men han ville icke höra på henne, utan ropade på den unge man som han hade till tjänare och sade: »Driven denna kvinna ut härifrån, och rigla du dörren efter henne.»
Och hon hade en fotsid livklädnad på sig; ty i sådana kåpor voro konungens döttrar klädda, så länge de voro jungfrur.
När tjänaren nu hade fört ut Tamar och riglat dörren efter henne,
tog hon aska och strödde på sitt huvud, och den fotsida livklädnaden som hon hade på sig rev hon sönder; och hon lade handen på sitt huvud och gick där ropande och klagande.
Då sade hennes broder Absalom till henne: »Har din broder Aminon varit hos dig?
Tig nu stilla, min syster; han är ju din broder.
Lägg denna sak icke så på sinnet.»
Så stannade då Tamar i sin broder Absaloms hus i svår sorg.
Men när konung David fick höra allt detta, blev han mycket vred.
Och Absalom talade intet med Amnon, varken gott eller ont, ty Absalom hatade Amnon, därför att denne hade kränkt hans syster Tamar.
Två år därefter hade Absalom fårklippning i Baal-Hasor, som ligger vid Efraim.
Och Absalom inbjöd då alla konungens söner.
Absalom kom till konungen och sade: »Din tjänare skall nu hava fårklippning; jag beder att konungen ville jämte sina tjänare gå med din tjänare.»
Men konungen svarade Absalom »Nej, min son, vi må icke allasammans gå med, ty vi vilja icke vara dig till besvär.»
Och fastän han bad honom enträget, ville han icke gå, utan gav honom sin avskedshälsning.
Då sade Absalom: »Om du icke vill, så låt dock min broder Amnon gå med oss.»
Konungen frågade honom: »Varför skall just han gå med dig?»
Men Absalom bad honom så enträget, att han lät Amnon och alla de övriga konungasönerna gå med honom.
Och Absalom bjöd sina tjänare och sade: »Sen efter, när Amnons hjärta bliver glatt av vinet; och när jag då säger till eder: 'Huggen ned Amnon', så döden honom utan fruktan.
Det är ju jag som bjuder eder det, varen frimodiga och skicken eder såsom käcka män.»
Och Absaloms tjänare gjorde med Amnon såsom Absalom hade bjudit.
Då stodo alla konungens söner upp och satte sig var och en på sin mulåsna och flydde.
Medan de ännu voro på väg, kom till David ett rykte om att Absalom hade huggit ned alla konungens söner, så att icke en enda av dem fanns kvar.
Då stod konungen upp och rev sönder sina kläder och lade sig på marken, under det att alla hans tjänare stodo där med sönderrivna kläder.
Men Jonadab, som var son till Davids broder Simea, tog till orda och sade: »Min herre må icke tänka att de hava dödat alla de unga männen, konungens söner, det är Amnon allena som är död.
Ty Absaloms uppsyn har bådat olycka ända ifrån den dag då denne kränkte hans syster Tamar.
Så må nu min herre konungen icke akta på detta som har blivit sagt, att alla konungens söner äro döda; nej, Amnon allena är död.»
Emellertid flydde Absalom. -- När nu mannen som stod på vakt lyfte upp sina ögon, fick han se mycket folk komma från vägen bakom honom, vid sidan av berget.
Då sade Jonadab till konungen: »Se, där komma konungens söner.
Såsom din tjänare sade, så har det gått till.»
Just när han hade sagt detta, kommo konungens söner; och de brusto ut i gråt.
Också konungen och alla hans tjänare gräto häftigt och bitterligen.
Men Absalom hade flytt och begivit sig till Talmai, Ammihurs son, konungen i Gesur.
Och David sörjde hela tiden sin son.
Sedan Absalom hade flytt och begivit sig till Gesur, stannade han där i tre år.
Och konung David avstod ifrån att draga ut mot Absalom, ty han tröstade sig över att Amnon var död.
Men Joab, Serujas son, märkte att konungens hjärta var vänt mot Absalom.
Då sände Joab till Tekoa och lät därifrån hämta en klok kvinna och sade till henne: »Låtsa att du har sorg, och kläd dig i sorgkläder och smörj dig icke med olja, utan skicka dig såsom en kvinna som i lång tid har haft sorg efter en död.
Gå så in till konungen och tala till honom såsom jag säger dig.»
Joab lade nu orden i hennes mun.
Och kvinnan från Tekoa talade med konungen; hon föll ned till jorden på sitt ansikte och bugade sig och sade: »Hjälp, o konung!»
Konungen sade till henne: »Vad fattas dig?»
Hon svarade: »Ack, jag är änka; min man är död.
Och din tjänarinna hade två söner; dessa båda kommo i träta med varandra ute på marken, där ingen fanns, som kunde träda emellan och hindra dem; den ene slog då ned den andre och dödade honom.
Och nu har hela släkten rest sig upp mot din tjänarinna, och de säga: 'Giv hit honom som slog ned sin broder, så att vi få döda honom, därför att han har tagit sin broders liv och dräpt honom; på det sättet förgöra vi ock arvingen.'
På det att efter min man varken namn eller efterkommande må finnas på jorden, vilja de utsläcka den gnista av mig, som ännu är kvar.»
Då sade konungen till kvinnan: »Gå hem igen; jag vill giva befallning om dig.»
Kvinnan från Tekoa sade till konungen: »På mig, o min herre konung, och på min faders hus vile missgärningen, men konungen och hans tron vare utan skuld.»
Konungen sade: »Om någon säger något åt dig, så för honom till mig; han skall sedan icke mer antasta dig.
Hon sade: »Ja, må konungen tänka på HERREN, sin Gud, så att blodshämnaren icke får göra olyckan större, och så att de icke förgöra min son.»
Då sade han: »Så sant HERREN lever, icke ett hår av din son skall falla på jorden.»
Men kvinnan sade: »Låt din tjänarinna tala ännu ett ord till min herre konungen.»
Han sade: »Tala.»
Då sade kvinnan: »Varför är du då så sinnad mot Guds folk?
När konungen talar så, då ligger ju däri att han själv bär på skuld, eftersom konungen icke låter sin förskjutne son komma tillbaka.
Vi måste ju alla dö och äro då såsom vatten som spilles på jorden, vilket icke kan samlas upp igen.
Men Gud tager icke livet bort, utan han tänker ut vad göras kan, för att den förskjutne icke må förbliva förskjuten och skild från honom.
Och att jag nu har kommit för att tala detta till min herre konungen, det har skett därför att folket förskräckte mig.
Då tänkte din tjänarinna: Jag vill dock tala med konungen; kanhända skall konungen uppfylla sin trälinnas önskan.
Ja, konungen skall lyssna till sin trälinna och rädda mig från den mans hand, som vill förgöra både mig och min son från Guds arvedel.
Och din tjänarinna tänkte: Min herre konungens ord skall giva mig ro.
Ty min herre konungen är lik Guds ängel däri att han hör allt, både gott och ont.
Och nu vare HERREN, din Gud, med dig.
Då svarade konungen och sade till kvinnan: »Dölj icke för mig något av det varom jag nu vill fråga dig.»
Kvinnan sade: »Min herre konungen tale.»
Då sade konungen: »Har icke Joab sin hand med i allt detta?»
Kvinnan svarade och sade: »Så sant du lever, min herre konung: om min Herre konungen talar något, så kan ingen komma undan det, vare sig åt höger eller åt vänster.
Ja, det är din tjänare Joab som har bjudit mig detta, och han har lagt i din tjänarinnas mun allt vad jag har sagt.
För att giva saken ett annat utseende har din tjänare Joab handlat på detta sätt; men min herre liknar i vishet Guds ängel och vet allt som sker på jorden.»
Så sade då konungen till Joab: »Välan, jag vill göra såsom du önskar.
Gå nu och för tillbaka den unge mannen Absalom.»
Då föll Joab ned till jorden på sitt ansikte och bugade sig och välsignade konungen; och Joab sade: »I dag märker din tjänare att jag har funnit nåd för dina ögon, min herre konung, eftersom konungen uppfyller sin tjänares önskan.»
Och Joab stod upp och begav sig till Gesur och förde Absalom till Jerusalem.
Men konungen sade: »Han får begiva sig till sitt hus, men han får icke komma inför mitt ansikte.
Då begav sig Absalom till sitt hus, och kom icke inför konungens ansikte.
Men i hela Israel fanns ingen så skön man som Absalom, ingen som man så mycket prisade: från hans fotblad upp till hans hjässa fanns icke något fel på honom
Och när han lät klippa håret på sitt huvud -- vid slutet av vart år lät han klippa det, ty det blev honom då så tungt att han måste låta klippa det -- så befanns det, att när man vägde håret från hans huvud, då vägde det två hundra siklar, efter konungsvikt.
Och åt Absalom föddes tre söner och en dotter, som fick namnet Tamar; hon var en skön kvinna.
När Absalom hade bott två hela år i Jerusalem utan att få komma inför konungens ansikte,
sände han bud efter Joab, i avsikt att skicka denne till konungen; men han ville icke komma till honom.
Och han sände bud ännu en gång, men han ville ändå icke komma.
Då sade han till sina tjänare: »I sen att Joab där har ett åkerstycke vid sidan av mitt, och på det har han korn; gån nu dit och tänden eld därpå.»
Så tände då Absaloms tjänare eld på åkerstycket.
Då stod Joab upp och gick hem till Absalom och sade till honom: »Varför hava dina tjänare tänt eld på mitt åkerstycke?»
Absalom svarade Joab: »Jag sände ju till dig och lät säga: Kom hit, så att jag kan skicka dig till konungen och låta säga: 'Varför fick jag komma hem från Gesur?
Det hade varit bättre för mig, om jag ännu vore kvar där.'
Nu vill jag komma inför konungens ansikte; och finnes någon missgärning hos mig, så må han döda mig.
Då gick Joab till konungen och sade honom detta.
Denne kallade då till sig Absalom, och han kom till konungen; och han föll ned för honom på sitt ansikte och bugade sig till jorden inför konungen.
Och konungen kysste Absalom.
En tid härefter skaffade Absalom sig vagn och hästar, därtill ock femtio man som löpte framför honom.
Och Absalom plägade bittida om morgonen ställa sig vid sidan av vägen som ledde till porten, och så ofta någon då var på väg till konungen med en rättssak som han ville hava avdömd, kallade Absalom honom till sig och frågade: »Från vilken stad är du?»
När han då svarade: »Din tjänare är från den och den av Israels stammar»,
sade Absalom till honom: »Din sak är visserligen god och rätt, men du har ingen som hör på dig hos konungen.»
Och Absalom tillade: »Ack om jag bleve satt till domare i landet!
Om då var och en som hade någon rätts- och domssak komme till mig, så skulle jag skaffa honom rättvisa.»
Och när någon gick fram för att buga sig för honom, räckte han ut sin hand och fattade i honom och kysste honom.
På detta sätt gjorde Absalom med alla israeliter som kommo för att få någon sak avdömd hos konungen.
Så förledde Absalom Israels män.
Fyrtio år voro nu förlidna, då Absalom en gång sade till konungen: »Låt mig begiva mig till Hebron för att där infria det löfte som jag har gjort åt HERREN.
Ty din tjänare gjorde ett löfte, när jag bodde i Gesur i Aram; jag sade: 'Om HERREN låter mig komma tillbaka till Jerusalem, så vill jag hålla en gudstjänst åt HERREN.'»
Konungen sade till honom: »Gå i frid.»
Då stod han upp och begav sig till Hebron.
Men Absalom sände ut hemliga budbärare till alla Israels stammar och lät säga: »När I hören basunen ljuda, så sägen: 'Nu har Absalom blivit konung i Hebron.'»
Och med Absalom hade följt två hundra män från Jerusalem, som voro inbjudna och följde med i all oskuld, utan att veta om någonting.
Medan Absalom offrade slaktoffren, sände han också och lät hämta giloniten Ahitofel, Davids rådgivare, från hans stad Gilo.
Och sammansvärjningen växte i styrka, och i allt större myckenhet gick folket över till Absalom.
Men en budbärare kom till David och sade: »Israels män hava vänt sina hjärtan till Absalom.»
Då sade David till alla sina tjänare, dem som han hade hos sig i Jerusalem: »Upp, låt oss fly, ty ingen annan räddning finnes för oss undan Absalom.
Skynden eder åstad, så att han icke med hast kommer över oss och för olycka över oss och slår stadens invånare med svärdsegg.»
Konungens tjänare svarade konungen: »Till allt vad min herre konungen behagar äro dina tjänare redo.
Då drog konungen ut, och allt hans husfolk följde honom; dock lämnade konungen kvar tio av sina bihustrur för att vakta huset.
Så drog då konungen ut, och allt folket följde honom; men de stannade vid Bet-Hammerhak.
Och alla hans tjänare tågade förbi på sidan om honom, så ock alla keretéerna och peletéerna; och alla gatiterna, sex hundra man, som hade följt med honom från Gat, tågade likaledes förbi framför konungen.
Då sade konungen till gatiten Ittai: »Varför går också du med oss?
Vänd om och stanna hos den som nu är konung; du är ju en främling och därtill landsflyktig från ditt hem.
I går kom du; skulle jag då i dag låta dig irra omkring med oss på var färd, nu då jag själv går jag vet icke vart?
Vänd tillbaka och för dina bröder tillbaka med dig; må nåd och trofasthet bevisas eder.»
Men Ittai svarade konungen och sade: »Så sant HERREN lever, och så sant min herre konungen lever: på den plats där min herre konungen är, där vill ock din tjänare vara, det må gälla liv eller död.»
Då sade David till Ittai: »Kom då och drag med.»
Och gatiten Ittai drog med jämte alla sina män och alla kvinnor och barn som han hade med sig.
Och hela landet grät högljutt, när allt folket drog fram.
Och då nu konungen gick över bäcken Kidron, gick ock allt folket över och tog vägen åt öknen.
Bland de andra såg man ock Sadok jämte alla leviterna, och de buro med sig Guds förbundsark; men de satte ned Guds ark -- varvid också Ebjatar kom ditupp -- till dess att allt folket hade hunnit draga fram ur staden.
Då sade konungen till Sadok: »För Guds ark tillbaka in i staden.
Om jag finner nåd för HERRENS ögon, låter han mig komma tillbaka, så att jag åter får se honom och hans boning.
Men om han säger så: 'Jag har icke behag till dig' -- se, då är jag redo; han göre då med mig såsom honom täckes.»
Och konungen sade till prästen Sadok: »Du är ju siare; vänd tillbaka till staden i frid.
Och din son Ahimaas och Ebjatars son Jonatan, båda edra söner, må följa med eder.
Se, jag vill dröja vid färjställena i öknen, till dess att ett budskap kommer från eder med underrättelser till mig.
Då förde Sadok och Ebjatar Guds ark tillbaka till Jerusalem och stannade där.
Men David gick gråtande uppför Oljeberget med överhöljt huvud ock bara fötter; och allt folket som följde med honom hade ock höljt över sina huvuden och gingo ditupp under gråt.
Och när man berättade för David att Ahitofel var med bland dem som hade sammansvurit sig med Absalom, sade David: »HERRE, gör Ahitofels råd till dårskap.»
När sedan David hade kommit upp på bergstoppen, där man plägade tillbedja Gud, då kom arkiten Husai emot honom, med sönderriven livklädnad och med jord på sitt huvud.
David sade till honom: »Om du går med mig, så bliver du mig till besvär.
Men om du vänder tillbaka till staden och säger till Absalom: 'Din tjänare vill jag vara, o konung; jag har förut varit din faders tjänare, men nu vill jag vara din tjänare', så kan du gagna mig med att göra Ahitofels råd om intet.
Där har du ju ock prästerna Sadok och Ebjatar; allt vad du får höra från konungens hus må du meddela prästerna Sadok och Ebjatar.
De hava ju ock där sina båda söner hos sig: Sadok har Ahimaas, och Ebjatar Jonatan; genom dem kunnen I sända mig bud om allt vad I fån höra.»
Så gick då Husai, Davids vän, in i staden.
Och jämväl Absalom drog in i Jerusalem.
När David hade gått framåt ett litet stycke från bergstoppen, då mötte honom Siba, Mefibosets tjänare, med ett par lastade åsnor, som buro två hundra bröd, ett hundra russinkakor, ett hundra fruktkakor och en vinlägel.
Då sade konungen till Siba: »Vad vill du med detta?»
Siba svarade: »Åsnorna skola vara för konungens husfolk till att rida på, brödet och fruktkakorna skola tjänarna hava att äta, och vinet skola de törstande hava att dricka i öknen.»
Konungen sade: »Men var är din herres son?»
Siba svarade konungen: »Han är kvar i Jerusalem; ty han tänkte: 'Nu skall Israels hus giva mig tillbaka min faders rike.'»
Då sade konungen till Siba: »Se, allt vad Mefiboset äger skall vara ditt.»
Siba svarade: »Jag faller ned för dig; låt mig finna nåd för dina ögon, min herre konung.»
När sedan konung David hade kommit till Bahurim, då trädde därifrån ut en man som var besläktad med Sauls hus och hette Simei, Geras son; han trädde fram och for ut i förbannelser.
Och han kastade stenar på David och på alla konung Davids tjänare, fastän allt folket och alla hjältarna omgåvo denne, både till höger och till vänster.
Och Simeis ord, när han förbannade honom, voro dessa: »Bort, bort, du blodsman, du ogärningsman!
HERREN låter nu allt Sauls hus' blod komma tillbaka över dig, du som har blivit konung i hans ställe; HERREN giver nu konungadömet åt din son Absalom.
Se, nu har du kommit i den olycka du förtjänade, ty en blodsman är du.»
Då sade Abisai, Serujas son, till konungen: »Varför skall den döda hunden där få förbanna min herre konungen?
Låt mig gå dit och hugga huvudet av honom.»
Men konungen svarade: »Vad haven I med mig att göra, I Serujas söner?
Om han förbannar, och om det är HERREN som har bjudit honom att förbanna David, vem törs då fråga: 'Varför gör du så?'
Och David sade ytterligare till Abisai och till alla sina tjänare: »Min son, han som har utgått från mitt eget liv, står mig ju efter livet; med huru mycket mer skäl då denne benjaminit!
Låten honom vara, må han förbanna; ty HERREN har befallt honom det.
Kanhända skall HERREN se till den orätt mig sker, så att HERREN åter giver mig lycka, till gengäld för den förbannelse som i dag uttalas över mig.»
Och David gick med sina män vägen fram, under det att Simei gick längs utmed berget, jämsides med honom, och for ut i förbannelser och kastade stenar och grus, där han gick jämsides med honom.
När så konungen, med allt folket som följde honom, hade kommit till Ajefim, rastade han där.
Men Absalom hade med allt sitt folk, Israels män, kommit till Jerusalem; han hade då också Ahitofel med sig.
När nu arkiten Husai, Davids vän, kom till Absalom, ropade Husai till Absalom: »Leve konungen!
Leve konungen!»
Absalom sade till Husai: »Är det så du visar din kärlek mot din vän?
Varför har du icke följt med din vän?»
Husai svarade Absalom: »Nej, den som HERREN och detta folk och alla Israels män hava utvalt, honom vill jag tillhöra, och hos honom vill jag stanna.
Och dessutom, vilken bör jag tjäna?
Bör jag icke tjäna inför hans son?
Jo, såsom jag har tjänat inför din fader, så vill jag ock göra det inför dig.»
Och Absalom sade till Ahitofel: »Given nu ett råd om vad vi skola göra.»
Ahitofel sade till Absalom: »Gå in till din faders bihustrur, som han har lämnat kvar för att vakta huset.
Då får hela Israel höra att du har gjort dig förhatlig för din fader, och så styrkes modet hos alla dem som hålla med dig.
Därefter slog man upp ett tält åt Absalom ovanpå taket, och så gick Absalom in till sin faders bihustrur inför hela Israels ögon.
Den tiden gällde nämligen ett råd som Ahitofel gav lika mycket som om man hade frågat Gud till råds; så mycket gällde vart råd av Ahitofel både för David och för Absalom.
Och Ahitofel sade till Absalom: »Låt mig utvälja tolv tusen män, så vill jag bryta upp och förfölja David i natt.
Då kan jag komma över honom och förskräcka honom, medan han är utmattad och modlös, och allt hans folk skall då taga till flykten; sedan kan jag döda konungen, när han står där övergiven.
Därefter skall jag föra allt folket tillbaka till dig.
Ty om det så går den man du söker, så är detta som om alla vände tillbaka; allt folket får då frid.»
Detta behagade Absalom och alla de äldste i Israel.
Likväl sade Absalom: »Kalla ock arkiten Husai hit, så att vi också få höra vad han har att säga.
När då Husai kom in till Absalom, sade Absalom till honom: »Så och så har Ahitofel talat. »Skola vi göra såsom han har sagt?
Varom icke, så tala du.»
Husai svarade Absalom: Det råd som Ahitofel denna gång har givit är icke gott.»
Och Husai sade ytterligare: »Du känner din fader och hans män, och vet att de äro hjältar och bistra såsom en björninna från vilken man har tagit ungarna ute på marken.
Och din fader är ju en krigsman som icke vilar med sitt folk under natten.
Nu har han säkerligen gömt sig i någon håla eller på något annat ställe.
Om nu redan i början några av folket här fölle, så skulle var och en som finge höra talas därom säga att det folk som följer Absalom har lidit ett nederlag;
och då skulle till och med den tappraste, den som hade mod såsom ett lejon, bliva högeligen förfärad; ty hela Israel vet att din fader är en hjälte, och att de som följa honom äro tappra män.
Därför är nu mitt råd: Låt hela Israel från Dan ända till Beer-Seba församla sig till dig, så talrikt som sanden vid havet; och själv må du draga med i striden.
När vi så drabba ihop med honom, varhelst han må påträffas, skola vi slå ned på honom, såsom daggen faller över marken; och då skall intet bliva kvar av honom och alla de män som äro med honom
Ja, om han också droge sig tillbaka in i någon stad, så skulle hela Israel kasta linor omkring den staden, och vi skulle draga den ned i dalen, till dess att icke minsta sten vore att finna därav.
Då sade Absalom och alla Israels män: »Arkiten Husais råd är bättre än Ahitofels råd.»
HERREN hade nämligen skickat det så, att Ahitofels goda råd gjordes om intet, för att HERREN skulle låta olycka komma över Absalom.
Och Husai sade till prästerna Sadok och Ebjatar: »Det och det rådet har Ahitofel givit Absalom och de äldste i Israel, men jag har givit det och det rådet.
Så sänden nu med hast bud och låten säga David: 'Stanna icke över natten vid färjställena i öknen, utan gå hellre över, för att icke konungen och allt hans folk må drabbas av fördärv.'»
Nu hade Jonatan och Ahimaas sitt tillhåll vid Rogelskällan, och en tjänstekvinna gick dit med budskap; sedan plägade de själva gå med budskapet till konung David.
Ty de tordes icke gå in i staden och visa sig där.
Men en gosse fick se dem och berättade det för Absalom.
Då gingo båda med hast sin väg och kommo in i en mans hus i Bahurim, som på sin gård hade en brunn; i den stego de ned.
Och hans hustru tog ett skynke och bredde ut det över brunnshålet och strödde gryn därpå, så att man icke kunde märka något.
Då nu Absaloms tjänare kommo in i huset till hustrun och frågade var Ahimaas och Jonatan voro, svarade hon dem: »De gingo över bäcken där.»
Då sökte de, men utan att finna, och vände så tillbaka till Jerusalem.
Men sedan de hade gått sin väg, stego de andra upp ur brunnen och gingo med sitt budskap till konung David; de sade till David: »Bryten upp och gån med hast över vattnet, ty det och det rådet har Ahitofel givit, till eder ofärd.»
Då bröt David upp med allt det folk han hade hos sig, och de gingo över Jordan; och om morgonen, när det blev dager, saknades ingen enda, utan alla hade kommit över Jordan.
Men när Ahitofel såg att man icke följde hans råd, sadlade han sin åsna och stod upp och for hem till sin stad, och sedan han hade beställt om sitt hus, hängde han sig.
Och när han var död, blev han begraven i sin faders grav.
Så hade nu David kommit till Mahanaim, när Absalom med alla Israels män gick över Jordan.
Men Absalom hade satt Amasa i Joabs ställe över hären.
Och Amasa var son till en man vid namn Jitra, en israelit, som hade gått in till Abigal, Nahas' dotter och Serujas, Joabs moders, syster.
Och Israel och Absalom lägrade sig i Gileads land.
Men när David kom till Mahanaim, hade Sobi, Nahas' son, från Rabba i Ammons barns land, och Makir, Ammiels son, från Lo-Debar, och Barsillai, en gileadit från Rogelim,
låtit föra dit sängar, skålar, lerkärl, så ock vete, korn, mjöl och rostade ax, ävensom bönor, linsärter och annat rostat,
därjämte honung, gräddmjölk, får och nötostar till mat åt David och hans folk; ty de tänkte: »Folket är hungrigt, trött och törstigt i öknen.
Och David mönstrade sitt folk och satte över- och underhövitsmän över dem.
Därefter lät David folket tåga åstad: en tredjedel under Joabs befäl, en tredjedel under Abisais, Serujas sons, Joabs broders, befäl, och en tredjedel under gatiten Ittais befäl.
Och konungen sade till folket: »Jag vill ock själv draga ut med eder.»
Men folket svarade: »Du får icke draga ut; ty om vi måste fly, aktar ingen på oss, och om hälften av oss bliver dödad, aktar man icke heller på oss, men du är nu så god som tio tusen av oss.
Därför är det nu bättre att du står redo att komma oss till hjälp från staden.
Då sade konungen till dem: »Vad I ansen vara bäst vill jag göra.»
Och konungen ställde sig vid sidan av porten, under det att allt folket drog ut i avdelningar på hundra och tusen.
Men konungen bjöd Joab, Abisai och Ittai och sade: »Faren nu varligt med den unge mannen Absalom.»
Och allt folket hörde huru konungen så bjöd alla hövitsmännen angående Absalom.
Så drog då folket ut på fältet mot Israel, och striden stod i Efraims skog.
Där blev Israels folk slaget av Davids tjänare, och många stupade där på den dagen: tjugu tusen man.
Och striden utbredde sig över hela den trakten; och skogen förgjorde mer folk, än svärdet förgjorde på den dagen.
Och Absalom kom i Davids tjänares väg.
Absalom red då på sin mulåsna; och när mulåsnan kom under en stor terebint med täta grenar, fastnade hans huvud i terebinten, så att han blev hängande mellan himmel och jord, ty mulåsnan som han satt på sprang sin väg.
Och en man fick se det och berättade för Joab och sade: »Jag såg där borta Absalom hänga i en terebint.»
Då sade Joab till mannen som berättade detta för honom: »Om du såg det, varför slog du honom då icke strax till jorden?
Jag skulle då gärna hava givit dig tio siklar silver och ett bälte.»
Men mannen svarade Joab: »Om jag ock finge väga upp tusen siklar silver i mina händer, skulle jag dock icke vilja uträcka min hand mot konungens son, ty konungen bjöd ju dig och Abisai och Ittai, så att vi hörde det: 'Tagen vara, I alla, på den unge mannen Absalom.'
Dessutom, om jag lömskt hade förgripit mig på hans liv, så hade du säkerligen lämnat mig i sticket, eftersom intet kan förbliva dolt för konungen.»
Joab sade: »Jag vill icke på detta sätt förhala tiden med dig.»
Därefter tog han tre spjut i sin hand och stötte dem i Absaloms bröst, medan denne ännu var vid liv, där han hängde under terebinten.
Sedan kommo tio unga män, Joabs vapendragare, ditfram, och av dem blev Absalom till fullo dödad.
Och Joab lät stöta i basunen, och folket upphörde att förfölja Israel, ty Joab ville skona folket.
Och de togo Absalom och kastade honom i en stor grop i skogen och staplade upp ett mycket stort stenröse över honom.
Men hela Israel flydde, var och en till sin hydda.
Och Absalom hade, medan han ännu levde, låtit resa åt sig en stod som står i Konungsdalen; ty han tänkte: »Jag har ingen son som kan bevara mitt namns åminnelse.
Den stoden hade han uppkallat efter sitt namn, och den heter ännu i dag Absaloms minnesvård.
Och Ahimaas, Sadoks son, sade: »Låt mig skynda åstad och förkunna för konungen glädjebudskapet att HERREN har dömt honom fri ifrån hans fienders hand.»
Men Joab svarade honom: »I dag bliver du ingen glädjebudbärare; en annan dag må du förkunna glädjebudskap, men denna dag förkunnar du icke något glädjebudskap, eftersom nu konungens son är död.»
Därefter sade Joab till en etiopier: »Gå och berätta för konungen vad du har sett.»
Då föll etiopiern ned för Joab och skyndade därpå åstad.
Men Ahimaas, Sadoks son; sade ännu en gång till Joab: »Låt också mig, vad än må ske, få skynda åstad, efter etiopiern.»
Joab sade: »Varför vill du skynda åstad, min son, då detta ju icke kan vara ett glädjebudskap som skaffar dig någon lön?»
Han svarade: »Vad än må ske vill jag skynda åstad.»
Då sade han till honom: »Så skynda då.»
Och Ahimaas skyndade åstad och tog vägen över Jordanslätten och hann om etiopiern.
Under tiden satt David inne i porten.
Och väktaren gick upp på porttaket invid muren; när han där lyfte upp sina ögon, fick han se en man komma ensam springande.
Väktaren ropade och förkunnade det för konungen.
Då sade konungen: »Är han ensam, så har han ett glädjebudskap att kungöra.»
Och han kom allt närmare.
Därefter fick väktaren se en annan man komma springande; då ropade väktaren till portvaktaren och sade: »Nu ser jag åter en man komma ensam springande.»
Konungen sade: »Denne är ock en glädjebudbärare.»
Och väktaren sade: »Efter sitt sätt att springa tyckes mig den förste vara Ahimaas, Sadoks son.»
Då sade konungen: »Det är en god man; han kommer säkerligen med ett gott glädjebudskap.»
Och Ahimaas ropade och sade till konungen: »Allt väl!»
Därefter föll han ned till Jorden på sitt ansikte inför konungen och sade: »Lovad vare HERREN, din Gud, som har prisgivit de människor som hade upplyft sin hand mot min herre konungen!»
Då frågade konungen: »Står det väl till med den unge mannen Absalom?»
Ahimaas svarade: »Jag såg en stor hop folk, när Joab avsände konungens andre tjänare och mig, din tjänare; men jag vet icke vad det var.»
Konungen sade: »Gå åt sidan och ställ dig där.»
Då gick han åt sidan och blev stående där
Just då kom etiopiern.
Och etiopiern sade: »Mottag, min herre konung, det glädjebudskapet att HERREN i dag har dömt dig fri ifrån alla de mäns hand, som hava rest sig upp mot dig.»
Konungen frågade etiopiern: »Står det väl till med den unge mannen Absalom?»
Etiopiern svarade: »Må det så gå med min herre konungens fiender och med alla som resa sig upp mot dig för att göra dig ont, såsom det har gått med den unge mannen.
Då blev konungen häftigt upprörd och gick upp i salen över porten och grät.
Och under det att han gick, ropade han så: »Min son Absalom, min son, min son Absalom!
Ack, att jag hade fått dö i ditt ställe!
Absalom, min son, min son!»
Och det blev berättat för Joab att konungen grät och sörjde Absalom.
Och segern blev på den dagen förbytt till sorg för allt folket, eftersom folket på den dagen fick höra sägas att konungen var bedrövad för sin sons skull.
Och folket smög sig på den dagen in i staden, såsom människor pläga göra, vilka hava vanärat sig, därigenom att de hava flytt under striden.
Men konungen hade skylt sitt ansikte; och konungen klagade med hög röst: »Min son Absalom!
Absalom, min son, min son!»
Då gick Joab in i huset till konungen och sade: »Du kommer i dag alla dina tjänares ansikten att rodna av skam, fastän de i dag hava räddat både ditt eget liv och dina söners och döttrars liv och dina hustrurs liv och dina bihustrurs liv.
Ty du älskar ju dem som hata dig, och hatar dem som älska dig.
I dag har du nämligen gjort kunnigt att dina hövitsmän och tjänare äro intet for dig, ty i dag märker jag, att om Absalom vore vid liv, men alla vi andra i dag hade omkommit, så skulle detta hava varit dig mer till behag.
Men stå nu upp, och gå ut och tala vänligt med dina tjänare; ty jag svär vid HERREN, att om du icke gör det, så skall icke en enda man stanna kvar hos dig över denna natt, och detta skall för dig bliva en större olycka än alla de olyckor som hava övergått dig från din ungdom ända till nu.»
Då stod konungen upp och satte sig i porten.
Och man gjorde kunnigt för allt folket och sade: »Konungen sitter nu i porten.»
Då kom allt folket inför konungen.
Men Israel hade flytt, var och en till sin hydda.
Och allt folket i alla Israels stammar begynte därefter förebrå varandra och säga: »Konungen har räddat oss från vara fienders hand och hjälpt oss ifrån filistéernas hand, och nu har han måst fly ur landet för Absalom.
Men Absalom, som vi hade smort till konung över oss, har blivit dödad i striden.
Varför sägen I då icke ett ord om att föra konungen tillbaka?»
Under tiden hade konung David sänt bud till prästerna Sadok och Ebjatar och låtit säga: »Talen så till de äldste i Juda: 'Varför skolen I vara de sista att hämta konungen tillbaka hem?
Ty vad hela Israel talar har redan kommit för konungen, där han bor.
I ären ju mina bröder, I ären ju mitt kött och ben.
Varför skolen I då vara de sista att hämta konungen tillbaka?'
Och till Amasa skolen I säga: 'Är du icke mitt kött och ben?
Gud straffe mig nu och framgent, om du icke för all din tid skall bliva härhövitsman hos mig i Joabs ställe.'»
Härigenom vann han alla Juda mäns hjärtan utan undantag, så att de sände detta budskap till konungen: »Vänd tillbaka, du själv med alla dina tjänare.»
Då vände konungen tillbaka och kom till Jordan; men Juda hade kommit till Gilgal för att möta konungen och föra konungen över Jordan.
Också Simei, Geras son, benjaminiten, som var från Bahurim, skyndade sig och drog ned med Juda män for att möta konung David.
Och med honom följde tusen man från Benjamin, ävensom Siba, vilken hade varit tjänare i Sauls hus, jämte hans femton söner och tjugu tjänare.
Dessa hade nu hastat ned till Jordan före konungen.
Och färjan gick över för att överföra konungens familj, och för att användas efter hans gottfinnande.
Men Simei, Geras son, föll ned inför konungen, när han skulle fara över Jordan,
och sade till konungen: »Må min herre icke tillräkna mig min missgärning, och icke tänka på huru illa din tjänare gjorde på den dag då min herre konungen drog ut från Jerusalem; må konungen icke akta därpå.
Ty din tjänare inser att jag då försyndade mig; därför har jag nu i dag först av hela Josefs hus kommit hitned för att möta min herre konungen.
Då tog Abisai, Serujas son, till orda och sade: »Skulle icke Simei dödas för detta?
Han har ju förbannat HERRENS smorde.»
Men David svarade: »Vad haven I med mig att göra, I Serujas söner, eftersom I i dag ären mig till hinders?
Skulle väl i dag någon dödas i Israel?
Vet jag då icke att jag i dag har blivit konung över Israel?»
Därefter sade konungen till Simei: »Du skall icke dö.»
Och konungen gav honom sin ed därpå.
Mefiboset, Sauls son, hade ock kommit ned för att möta konungen.
Han hade varken ansat sina fötter eller sitt skägg, ej heller hade han låtit två sina kläder allt ifrån den dag då konungen drog bort, ända till den dag då han kom igen i frid.
När han nu kom till Jerusalem för att möta konungen, sade konungen till honom: »Varför följde du icke med mig, Mefiboset?»
Han svarade: »Min herre konung, min tjänare bedrog mig.
Ty din tjänare sade: 'Jag vill sadla min åsna och sätta mig på den och så begiva mig till konungen'; din tjänare är ju halt.
Men han har förtalat din tjänare hos min herre konungen.
Min herre konungen är ju dock såsom Guds ängel; så gör nu vad dig täckes.
Ty hela min faders hus förtjänade intet annat än döden av min herre konungen, och likväl lät du din tjänare sitta bland dem som få äta vid ditt bord.
Vad har jag då rätt att ytterligare begära, och varom kan jag väl ytterligare ropa till konungen?»
Konungen sade till honom: »Varför ordar du ytterligare härom?
Jag säger att du och Siba skolen dela jordagodset.»
Då sade Mefiboset till konungen: »Han må gärna taga alltsammans, sedan nu min herre konungen har kommit hem igen i frid.»
Gileaditen Barsillai hade ock farit ned från Rogelim och drog sedan med konungen till Jordan, för att få ledsaga honom över Jordan.
Barsillai var då mycket gammal: åttio år.
Han hade sörjt för konungens behov, medan denne uppehöll sig i Mahanaim, ty han var en mycket rik man.
Konungen sade nu till Barsillai: »Du skall draga med mig, så skall jag sörja för dina behov hemma hos mig i Jerusalem.»
Men Barsillai svarade konungen: »Huru många år kan jag väl ännu hava att leva, eftersom jag skulle följa med konungen upp till Jerusalem?
Jag är nu åttio år gammal; kan jag då känna skillnad mellan bättre och sämre, eller har väl din tjänare någon smak för vad jag äter eller för vad jag dricker?
Eller kan jag ännu njuta av att höra sångare och sångerskor sjunga?
Varför skulle din tjänare då ytterligare bliva min herre konungen till besvär?
Allenast för en stund vill din tjänare fara med konungen över Jordan.
Varför skulle väl konungen giva mig en sådan vedergällning?
Låt din tjänare vända tillbaka, så att jag får dö i min stad, där jag har min faders och min moders grav.
Men se här är din tjänare Kimham, låt honom få draga med min herre konungen; och gör för honom vad dig täckes.»
Då sade konungen: »Så må då Kimham draga med mig, och jag skall göra för honom vad du vill.
Och allt vad du begär av mig skall jag göra dig.»
Därefter gick allt folket över Jordan, och konungen själv gick också över.
Och konungen kysste Barsillai och tog avsked av honom.
Sedan vände denne tillbaka hem igen.
Så drog nu konungen till Gilgal, och Kimham följde med honom, så ock allt Juda folk.
Och de, jämte hälften av Israels folk, förde konungen ditöver.
Men då kommo alla de övriga israeliterna till konungen och sade till honom: »Varför hava våra bröder, Juda män, fått hemligen bemäktiga sig dig och föra konungen och hans familj, tillika med alla Davids män, över Jordan?»
Alla Juda män svarade Israels män: »Konungen står ju oss närmast; varför vredgens I då häröver?
Hava vi levat på konungen eller skaffat oss någon vinning genom honom?»
Då svarade Israels män Juda män och sade: »Tio gånger större del än I hava vi i den som är konung, alltså ock i David.
Varför haven I då ringaktat oss?
Och voro icke vi de som först talade om att hämta vår konung tillbaka?»
Men Juda män läto ännu hårdare ord falla än Israels män.
Nu hände sig att där fanns en illasinnad man vid namn Seba, Bikris son, en benjaminit.
Denne stötte i basun och sade: »Vi hava ingen del i David och ingen arvslott i Isais son.
Israel drage hem, var och en till sin hydda.»
Då övergåvo alla Israels män David och följde Seba, Bikris son; men Juda män höllo sig till sin konung och följde honom från Jordan ända till Jerusalem.
Så kom David hem igen till Jerusalem.
Och konungen tog då de tio bihustrur som han hade lämnat kvar för att vakta huset, och satte in dem i ett särskilt hus till att där förvaras; och han gav dem underhåll, men gick icke in till dem.
Där förblevo de nu instängda till sin dödsdag och levde redan under hans livstid såsom änkor.
Och konungen sade till Amasa: »Båda upp åt mig Juda män inom tre dagar, och inställ dig sedan själv här.»
Amasa begav sig då åstad för att uppbåda Juda; men när han dröjde utöver den tid som hade blivit honom förelagd,
sade David till Abisai: »Nu kommer Seba, Bikris son, att bliva farligare för oss än Absalom.
Tag du din herres tjänare och sätt efter honom, så att han icke bemäktigar sig några befästa städer och tillfogar oss för stor skada.»
Alltså drogo Joabs män tillika med keretéerna och peletéerna och alla hjältarna ut efter honom; de drogo ut från Jerusalem för att sätta efter Seba, Bikris son.
Men när de hade hunnit till den stora stenen vid Gibeon, kom Amasa emot dem.
Joab var då klädd i livrocken som plägade utgöra hans dräkt, och ovanpå den hade han ett bälte, med ett svärd i skidan, bundet över sina länder; men när han gick fram, föll det ut.
Och Joab sade till Amasa: »Står det väl till med dig, min broder?»
Därvid fattade Joab Amasa i skägget med högra handen såsom för att kyssa honom.
Och då Amasa icke tog sig till vara för det svärd som Joab hade i sin andra hand, gav denne honom därmed en stöt i underlivet, så att hans inälvor runno ut på jorden.
Så dog han, utan att den andre behövde giva honom någon ytterligare stöt.
Därefter fortsatte Joab och hans broder Abisai att förfölja Seba, Bikris son.
Men en av Joabs tjänare stod kvar därbredvid och ropade: »Var och en som är Joabs vän och håller med David, han följe efter Joab.»
Nu låg Amasa sölad i sitt blod mitt på vägen; och mannen såg allt folket stannade.
Då förde han Amasa undan från vägen in på åkern och kastade ett kläde över honom, eftersom han såg huru alla de som kommo därförbi stannade.
Så snart han var bortskaffad från vägen, drogo alla förbi och följde Joab för att sätta efter Seba, Bikris son.
Denne drog emellertid genom alla Israels stammar till Abel och Bet-Maaka och genom hela Habberim; och folk samlade sig och följde honom ända ditin.
Men de kommo och belägrade honom där i Abel vid Bet-Hammaaka och kastade upp mot staden en vall, som reste sig inemot yttermuren.
Och allt Joabs folk arbetade på att förstöra muren och kullstöta den.
Då ropade en klok kvinna från staden: »Hören!
Hören!
Sägen till Joab att han kommer hit, så att jag får tala med honom.»
När han då kom fram till kvinnan, frågade hon: »Är du Joab?»
Han svarade: »Ja.»
Hon sade till honom: »Hör din tjänarinnas ord.»
Han svarade: »Jag hör.»
Då sade hon: »Fordom plägade man säga så: 'I Abel skall man fråga till råds'; sedan kunde man utföra sina planer.
Vi äro de fridsammaste och trognaste i Israel, och du söker att förgöra en stad som är en moder i Israel.
Varför vill du förstöra HERRENS arvedel?»
Joab svarade och sade: »Bort det, bort det, att jag skulle vilja förstöra och fördärva!
Det är icke så, utan en man från Efraims bergsbygd vid namn Seba, Bikris son, har rest sig upp mot konung David; utlämnen allenast honom, så vill jag draga bort ifrån staden.»
Kvinnan svarade Joab: »Hans huvud skall strax bliva utkastat till dig över muren.»
Sedan vände sig kvinnan med sitt kloka råd till allt folket, och de höggo huvudet av Seba, Bikris son, och kastade ut det till Joab.
Då stötte denne i basunen, och krigsfolket skingrade sig och drog bort ifrån staden, var och en till sin hydda.
Och Joab vände tillbaka till konungen i Jerusalem.
Joab hade nu befälet över hela krigshären i Israel, och Benaja, Jojadas son, hade befälet över keretéerna och peletéerna.
Adoram hade uppsikten över de allmänna arbetena, och Josafat, Ahiluds son, var kansler.
Seja var sekreterare, och Sadok och Ebjatar voro präster.
Dessutom var ock jairiten Ira präst hos David.
Men under Davids tid uppstod en hungersnöd, som varade oavbrutet i tre år; då sökte David HERRENS ansikte.
HERREN svarade: »För Sauls och hans blodbefläckade hus' skull sker detta, därför att han dödade gibeoniterna.
Då kallade konungen till sig gibeoniterna och talade med dem.
Men gibeoniterna voro icke israeliter, utan en kvarleva av amoréerna och fastän Israels barn hade givit dem sin ed, hade Saul, i sin nitälskan för Israels barn och för Juda, försökt att nedgöra dem.
David sade nu till gibeoniterna: »Vad skall jag göra för eder, och varmed skall jag bringa försoning, så att I välsignen HERRENS arvedel?»
Gibeoniterna svarade honom: »Vi fordra icke silver och guld av Saul och hans hus, ej heller hava vi rätt att döda någon man i Israel.»
Han frågade: »Vad begären I då att jag skall göra för eder?»
De svarade konungen: »Den man som ville förgöra oss, och som stämplade mot oss, för att vi skulle bliva utrotade och icke mer hava bestånd någonstädes inom Israels land,
av hans söner må sju utlämnas till oss, så att vi få upphänga dem för HERREN i Sauls, HERRENS utvaldes, Gibea.»
Konungen sade: »Jag skall utlämna dem.»
Men konungen skonade Mefiboset, Sauls son Jonatans son, för den ed vid HERREN, som de, David och Jonatan, Sauls son, hade svurit varandra.
Däremot tog konungen de två söner, Armoni och Mefiboset, som Rispa, Ajas dotter, hade fött åt Saul, och de fem söner som Mikal, Sauls dotter, hade fött åt meholatiten Adriel, Barsillais son
och överlämnade dem åt gibeoniterna, och dessa upphängde dem på berget inför HERREN, så att de omkommo, alla sju på en gång.
Och det var under de första skördedagarna, när kornskörden begynte, som de blevo dödade.
Då tog Rispa, Ajas dotter, sin sorgdräkt och hade den till sitt läger ovanpå klippan från det att skörden begynte, ända till dess att vattnet strömmade ned över dem från himmelen; och hon tillstadde icke himmelens fåglar att slå ned på dem om dagen, ej heller markens vilda djur att göra det om natten.
När det blev berättat för David vad Rispa, Ajas dotter, Sauls bihustru, hade gjort
begav sig David åstad och hämtade Sauls och hans son Jonatans ben från borgarna i Jabes i Gilead.
Dessa hade nämligen i hemlighet tagit deras kroppar bort ifrån den öppna platsen i Bet-San, där filistéerna hade hängt upp dem, när filistéerna slogo Saul på Gilboa.
Och då han hade fört Sauls och hans son Jonatans ben upp därifrån, samlade man ock ihop de upphängdas ben.
Sedan begrov man Sauls och hans son Jonatans ben i Benjamins land, i Sela, i hans fader Kis' grav; man gjorde allt vad konungen hade bjudit.
Och därefter hörde Gud landets bön.
Åter uppstod krig mellan filistéerna och Israel.
Och David drog ned med sina tjänare, och de stridde mot filistéerna.
Men David blev trött;
och Jisbo-Benob, en av rafaéernas avkomlingar, vilkens lans vägde tre hundra siklar koppar, och som var iklädd en ny rustning, tänkte då döda David.
Men Abisai, Serujas son, kom honom till hjälp och slog filistéen till döds.
Då besvuro Davids män honom att han icke mer skulle draga ut med dem i striden, så att han icke utsläckte Israels lampa.
Därefter stod åter en strid med filistéerna vid Gob; husatiten Sibbekai slog då ned Saf, en av rafaéernas avkomlingar.
Åter stod en strid med filistéerna vid Gob; Elhanan, Jaare-Oregims son, betlehemiten, slog då ned gatiten Goljat, som hade ett spjut vars skaft liknade en vävbom.
Åter stod en strid vid Gat.
Där var en reslig man som hade sex fingrar på var hand och sex tår på var fot, eller tillsammans tjugufyra; han var ock en avkomling av rafaéerna.
Denne smädade Israel; då blev han nedgjord av Jonatan, son till Simeai, Davids broder.
Dessa fyra voro avkomlingar av rafaéerna i Gat; och de föllo för Davids och hans tjänares hand.
Och David talade till HERREN denna sångs ord, när HERREN hade räddat honom från alla hans fienders hand och från Sauls hand.
Han sade: HERRE, du mitt bergfäste, min borg och min räddare,
Gud, du min klippa, till vilken jag tager min tillflykt, min sköld och min frälsnings horn, mitt värn och min tillflykt, min frälsare, du som frälsar mig från våldet!
HERREN, den högtlovade, åkallar jag, och från mina fiender bliver jag frälst.
Ty dödens bränningar omvärvde mig, fördärvets strömmar förskräckte mig,
dödsrikets band omslöto mig, dödens snaror föllo över mig.
Men jag åkallade HERREN i min nöd, ja, jag gick med min åkallan till min Gud.
Och han hörde från sin himmelska boning min röst, och mitt rop kom till hans öron.
Då skalv jorden och bävade, himmelens grundvalar darrade; de skakades, ty hans vrede var upptänd.
Rök steg upp från hans näsa och förtärande eld från hans mun, eldsglöd ljungade från honom.
Och han sänkte himmelen och for ned och töcken var under hans fötter.
Han for på keruben och flög, han sågs komma på vindens vingar
Och han gjorde mörker till en hydda som omslöt honom: vattenhopar, tjocka moln.
Ur glansen framför honom ljungade eldsglöd.
HERREN dundrade från himmelen den Högste lät höra sin röst.
Han sköt pilar och förskingrade dem, ljungeld och förvirrade dem.
Havets bäddar kommo i dagen, jordens grundvalar blottades, för HERRENS näpst, för hans vredes stormvind.
Han räckte ut sin hand från höjden och fattade mig, han drog mig upp ur de stora vattnen.
Han räddade mig från min starke fiende, från mina ovänner, ty de voro mig övermäktiga.
De överföllo mig på min olyckas dag, men HERREN blev mitt stöd.
Han förde mig ut på rymlig plats han räddade mig, ty han hade behag till mig.
HERREN lönar mig efter min rättfärdighet; efter mina händers renhet vedergäller han mig.
Ty jag höll mig på HERRENS vägar och avföll icke från min Gud i ogudaktighet;
nej, alla hans rätter hade jag för ögonen, och från hans stadgar vek jag icke av.
Så var jag ostrafflig för honom och tog mig till vara för missgärning.
Därför vedergällde mig HERREN efter min rättfärdighet, efter min renhet inför hans ögon.
Mot den fromme bevisar du dig from, mot en ostrafflig hjälte bevisar du dig ostrafflig.
Mot den rene bevisar du dig ren, men mot den vrånge bevisar du dig avog.
och du frälsar ett betryckt folk, men dina ögon äro emot de stolta, till att ödmjuka dem.
Ja, du, HERRE, är min lampa; ty HERREN gör mitt mörker ljust.
Ja, med dig kan jag nedslå härskaror, med min Gud stormar jag murar.
Guds väg är ostrafflig, HERRENS tal är luttrat.
En sköld är han för alla som taga sin tillflykt till honom.
Ty vem är Gud förutom HERREN, och vem är en klippa förutom vår Gud?
Gud, du som var mitt starka värn och ledde den ostrafflige på hans väg,
du som gjorde hans fötter såsom hindens och ställde mig på mina höjder,
du som lärde mina händer att strida och mina armar att spänna kopparbågen!
Du gav mig din frälsnings sköld och din bönhörelse gjorde mig stor,
du skaffade rum för mina steg, där jag gick, och mina fötter vacklade icke.
Jag förföljde mina fiender och förgjorde dem; jag vände icke tillbaka, förrän jag hade gjort ände på dem.
Ja, jag gjorde ände på dem och slog dem, så att de icke mer reste sig; de föllo under mina fötter.
Du omgjordade mig med kraft till striden, du böjde mina motståndare under mig.
Mina fiender drev du på flykten för mig, dem som hatade mig förgjorde jag.
De sågo sig omkring, men det fanns ingen som frälste; efter HERREN, men han svarade dem icke.
Och jag stötte dem sönder till stoft på jorden, jag krossade och förtrampade dem såsom orenlighet på gatan.
Du räddade mig ur mitt folks strider, du bevarade mig till ett huvud över hedningar; folkslag som jag ej kände blevo mina tjänare.
Främlingar visade mig underdånighet; vid blotta ryktet hörsammade de mig.
Ja, främlingarnas mod vissnade bort; de omgjordade sig och övergåvo sina borgar.
HERREN lever!
Lovad vare min klippa, upphöjd vare Gud, min frälsnings klippa!
Gud, som har givit mig hämnd och lagt folken under mig;
du som har fört mig ut från mina fiender och upphöjt mig över mina motståndare, räddat mig från våldets man!
Fördenskull vill jag tacka dig, HERRE, bland hedningarna, och lovsjunga ditt namn.
Ty du giver din konung stor seger och gör nåd mot din smorde, mot David och hans säd till evig tid.
Dessa voro Davids sista ord: Så säger David, Isais son, så säger den man som blev högt upphöjd, Jakobs Guds smorde, Israels ljuvlige sångare:
HERRENS Ande har talat genom mig, och hans ord är på min tunga;
Israels Gud har så sagt, Israels klippa har så talat till mig: »Den som råder över människorna rätt, den som råder i Guds fruktan,
han är lik morgonens ljus, när solen går upp, en morgon utan moln, då jorden grönskar genom solsken efter regn.
Ja, är det icke så med mitt hus inför Gud?
Han har ju upprättat med mig ett evigt förbund, i allo stadgat och betryggat.
Ja, visst skall han låta all frälsning och glädje växa upp åt mig.
Men de onda äro allasammans lika bortkastade törnen, som man ej vill taga i med handen.
Och måste man röra vid dem, så rustar man sig med järn och med spjutskaft, och bränner sedan upp dem i eld på stället.
Dessa äro namnen på Davids hjältar: Joseb-Bassebet, en takemonit, den förnämste bland kämparna, han som svängde sitt spjut över åtta hundra som hade blivit slagna på en gång.
Och näst honom kom Eleasar, son till Dodi, son till en ahoait.
Han var en av de tre hjältar som voro med David, när de blevo smädade av filistéerna, som där hade församlat sig till strid; Israels män drogo sig då tillbaka.
Men han höll stånd och högg in på filistéerna, till dess att hans hand blev så trött att den var såsom faststelnad vid svärdet; och HERREN beredde så en stor seger på den dagen.
Sedan hade folket allenast att vända om och följa med honom för att plundra.
Och efter honom kom Samma, son till Age, en hararit.
En gång hade filistéerna församlat sig, så att de utgjorde en hel skara.
Och där var ett åkerstycke, fullt med linsärter.
Och folket flydde för filistéerna.
Då ställde han sig mitt på åkerstycket och försvarade det och slog filistéerna; och HERREN beredde så en stor seger.
En gång drogo tre av de trettio förnämsta männen ned och kommo vid skördetiden till David vid Adullams grotta, medan en skara filistéer var lägrad i Refaimsdalen.
Men David var då på borgen, under det att en filisteisk utpost fanns i Bet-Lehem.
Och David greps av lystnad och sade: »Ack att någon ville giva mig vatten att dricka från brunnen vid Bet-Lehems stadsport!»
Då bröto de tre hjältarna sig igenom filistéernas läger och hämtade vatten ur brunnen vid Bet-Lehems stadsport och togo det och buro det till David.
Men han ville icke dricka det, utan göt ut det såsom ett drickoffer åt HERREN.
Han sade nämligen: »Bort det, HERRE, att jag skulle göra detta!
Skulle jag dricka de mäns blod, som gingo åstad med fara för sina liv?»
Och han ville icke dricka det.
Sådana ting hade de tre hjältarna gjort.
Abisai, broder till Joab, Serujas son, var den förnämste av tre andra; han svängde en gång sitt spjut över tre hundra som hade blivit slagna.
Och han hade ett stort namn bland de tre.
Han var visserligen mer ansedd än någon annan i detta tretal, och han var de andras hövitsman, men upp till de tre första kom han dock icke.
Och Benaja, son till Jojada, som var son till en tapper, segerrik man från Kabseel; han slog ned de två Arielerna i Moab, och det var han som en snövädersdag steg ned och slog ihjäl lejonet i brunnen.
Han slog ock ned den egyptiske mannen som var så ansenlig att skåda.
Fastän egyptiern hade ett spjut i handen, gick han ned mot honom, väpnad allenast med sin stav.
Och han ryckte spjutet ur egyptierns hand och dräpte honom med hans eget spjut.
Sådana ting hade Benaja, Jojadas son, gjort.
Och han hade ett stort namn bland de tre hjältarna.
Han var mer ansedd än någon av de trettio, men upp till de tre första kom han icke.
Och David insatte honom i sin livvakt.
Till de trettio hörde: Asael, Joabs broder; Elhanan, Dodos son, från Bet-Lehem;
haroditen Samma; haroditen Elika;
peletiten Heles; tekoaiten Ira, Ickes' son;
anatotiten Abieser; husatiten Mebunnai;
ahoaiten Salmon; netofatiten Maherai;
netofatiten Heleb, Baanas son; Ittai, Ribais son, från Gibea i Benjamins barns stam;
Benaja, en pirgatonit; Hiddai från Gaas' dalar;
arabatiten Abi-Albon; barhumiten Asmavet;
saalboniten Eljaba; Bene-Jasen; Jonatan;
harariten Samma; arariten Ahiam, Sarars son;
Elifelet, son till Ahasbai, maakatitens son; giloniten Eliam, Ahitofels son;
Hesro från Karmel; arabiten Paarai;
Jigeal, Natans son, från Soba; gaditen Bani;
ammoniten Selek; beerotiten Naharai, vapendragare åt Joab, Serujas son;
jeteriten Ira; jeteriten Gareb;
hetiten Uria.
Tillsammans utgjorde de trettiosju.
Men HERRENS vrede upptändes åter mot Israel, så att han uppeggade David mot dem och sade: »Gå åstad och räkna Israel och Juda.»
Då sade konungen till Joab, hövitsmannen för hans här: »Far igenom alla Israels stammar, från Dan ända till Beer-Seba, och anställen en folkräkning, så att jag får veta huru stor folkmängden är.»
Joab svarade konungen: »Må HERREN, din Gud, föröka detta folk hundrafalt, huru talrikt det än är, och må min herre konungen få se detta med egna ögon.
Men varför har min herre konungen fått lust till sådant?»
Likväl blev konungens befallning gällande, trots Joab och härens andra hövitsmän; alltså drog Joab jämte härens andra hövitsmän ut i konungens tjänst för att anställa folkräkning i Israel.
Och de gingo över Jordan och lägrade sig vid Aroer, på högra sidan om staden i Gads dal, och åt Jaeser till.
Därifrån kommo de till Gilead och Tatim-Hodsis land; sedan kommo de till Dan-Jaan och så runt omkring till Sidon.
Därefter kommo de till Tyrus' befästningar och till hivéernas och kananéernas alla städer; slutligen drogo de till Beer-Seba i Juda sydland.
Och sedan de så hade farit igenom hela landet, kommo de efter nio månader och tjugu dagar hem till Jerusalem.
Och Joab uppgav för konungen vilken slutsumma folkräkningen utvisade: i Israel funnos åtta hundra tusen stridbara, svärdbeväpnade män, och Juda män voro fem hundra tusen.
Men Davids samvete slog honom, sedan han hade låtit räkna folket, och David sade till HERREN: »Jag har syndat storligen i vad jag har gjort; men tillgiv nu, HERRE, din tjänares missgärning, ty jag har handlat mycket dåraktigt.»
Då nu David stod upp om morgonen, hade HERRENS ord kommit till profeten Gad, Davids siare; han hade sagt:
»Gå och tala till David: Så säger HERREN: Tre ting förelägger jag dig; välj bland dem ut åt dig ett som du vill att jag skall göra dig.»
Då gick Gad in till David och förkunnade detta för honom.
Han sade till honom: »Vill du att hungersnöd under sju år skall komma i ditt land?
Eller att du i tre månader skall nödgas fly för dina ovänner, medan de förfölja dig?
Eller att pest i tre dagar skall hemsöka ditt land?
Betänk nu och eftersinna vilket svar jag skall giva honom som har sänt mig.»
David svarade Gad: »Jag är i stor vånda.
Men låt oss då falla i HERRENS hand, ty hans barmhärtighet är stor; i människohand vill jag icke falla.»
Så lät då HERREN pest komma i Israel, från morgonen intill den bestämda tiden; därunder dogo av folket, ifrån Dan ända till Beer-Seba, sjuttio tusen män.
Men när ängeln räckte ut sin hand över Jerusalem för att fördärva det, ångrade HERREN det onda, och han sade till ängeln, folkets fördärvare: »Det är nog; drag nu din hand tillbaka.»
Och HERRENS ängel var då vid jebuséen Araunas tröskplats.
Men när David fick se ängeln som slog folket, sade han till HERREN så: »Det är ju jag som har syndat, det är jag som har gjort illa; men dessa, min hjord, vad hava de gjort?
Må din hand vända sig mot mig och min faders hus.»
Och Gad kom till David samma dag och sade till honom: »Gå åstad och res ett altare åt HERREN på jebuséen Araunas tröskplats.»
Och David gick åstad efter Gads ord, såsom HERREN hade bjudit.
När Arauna nu blickade ut och fick se att konungen och hans tjänare kommo till honom, gick han ut och föll ned till jorden på sitt ansikte för konungen.
Och Arauna sade: »Varför kommer min herre konungen till sin tjänare?»
David svarade: »För att köpa tröskplatsen av dig och där bygga ett altare åt HERREN; och må så hemsökelsen upphöra bland folket.»
Då sade Arauna till David: »Min herre konungen tage till sitt offer vad honom täckes.
Se här äro fäkreaturen till brännoffer, och här äro tröskvagnarna, jämte fäkreaturens ok, till ved.
Alltsammans, o konung, giver Arauna åt konungen.»
Och Arauna sade ytterligare till konungen: »Må HERREN, din Gud, vara dig nådig.»
Men konungen svarade Arauna: »Nej, jag vill köpa det av dig för ett bestämt pris; ty jag vill icke offra åt HERREN, min Gud, brännoffer som jag har fått för intet.»
Och David köpte tröskplatsen och fäkreaturen för femtio siklar silver.
Och David byggde där ett altare åt HERREN och offrade brännoffer och tackoffer.
Och HERREN lyssnade till landets bön, och hemsökelsen upphörde bland Israel.
Konung David var nu gammal och kommen till hög ålder; och ehuru man höljde täcken över honom, kunde han dock icke hålla sig varm.
Då sade hans tjänare till honom: »Må man för min herre konungens räkning söka upp en ung kvinna, en jungfru, som kan bliva konungens tjänarinna och sköta honom.
Om hon får ligga i din famn, så bliver min herre konungen varm»
Så sökte de då över hela Israels land efter en skön flicka; och de funno Abisag från Sunem och förde henne till konungen.
Hon var en mycket skön flicka, och hon skötte nu konungen och betjänade honom, men konungen hade intet umgänge med henne.
Men Adonia, Haggits son, hov sig upp och sade: »Det är jag som skall bliva konung.»
Och han skaffade sig vagnar och ryttare, därtill ock femtio man som löpte framför honom.
Hans fader hade aldrig velat bedröva honom med att säga: »Varför gör du så?»
Han var ock mycket fager; och hans moder hade fött honom näst efter Absalom.
Och han begynte underhandla med Joab, Serujas son, och med prästens Ebjatar, och dessa slöto sig till Adonia och understödde honom.
Men prästen Sadok och Benaja, Jojadas son, samt profeten Natan, Simei, Rei och Davids hjältar höllo icke med Adonia.
Och Adonia slaktade får och fäkreatur och gödkalvar vid Soheletstenen, som ligger vid Rogelskällan; och han inbjöd dit alla sina bröder, konungens söner, och alla de Juda män som voro i konungens tjänst.
Men profeten Natan, Benaja, hjältarna och sin broder Salomo inbjöd han icke.
Då sade Natan så till Bat-Seba, Salomos moder: »Du har väl hört att Adonia, Haggits son, har blivit konung, utan att vår herre David vet därom?
Men jag vill nu giva dig ett råd, för att du må kunna rädda ditt liv och din son Salomos liv.
Gå in till konung David och säg till honom: 'Har du icke, min herre konung, själv med ed lovat din tjänarinna och sagt: Din son Salomo skall bliva konung efter mig; han skall sitta på min tron?
Varför har då Adonia blivit konung?'
Och medan du ännu är där och talar med konungen, skall jag efter dig komma in och bekräfta dina ord.»
Så gick då Bat-Seba in till konungen, i kammaren.
Konungen var nu mycket gammal; och Abisag från Sunem betjänade konungen.
Och Bat-Seba bugade sig och föll ned för konungen.
Då frågade konungen: »Vad önskar du?»
Hon sade till honom: »Min herre, du har ju själv lovat din tjänarinna med en ed vid HERREN, din Gud: 'Din son Salomo skall bliva konung efter mig; han skall sitta på min tron.'
Men se, nu har Adonia blivit konung, fastän du, min herre konung, ännu icke har fått veta det.
Och han har slaktat tjurar och gödkalvar och får i myckenhet, och han har inbjudit alla konungens söner och prästen Ebjatar och härhövitsmannen Joab; men din tjänare Salomo har han icke inbjudit.
På dig, min herre konung, äro nu hela Israels ögon riktade, i förväntan att du skall kungöra för dem vem som skall sitta på min herre konungens tron efter honom.
Eljest torde hända, att när min herre konungen har gått till vila hos sina fäder, då bliva jag och min son Salomo hållna såsom brottslingar.»
Medan hon ännu höll på att tala med konungen, kom profeten Natan.
Och man anmälde det för konungen och sade: »Profeten Natan är här.»
När han så kom inför konungen, föll han ned till jorden på sitt ansikte för konungen.
Och Natan sade: »Min herre konung, är det väl du som har sagt att Adonia skall bliva konung efter dig, och att han skall sitta på din tron?
Ty han har i dag gått ned och slaktat tjurar och gödkalvar och får i myckenhet, och har inbjudit alla konungens söner och härhövitsmännen och prästen Ebjatar, och de hålla nu på med att äta och dricka hos honom; och de ropa: 'Leve konung Adonia!'
Men mig, din tjänare, och prästen Sadok och Benaja, Jojadas son, och din tjänare Salomo har han icke inbjudit.
Kan väl detta hava utgått från min herre konungen, utan att du har låtit dina tjänare vet vem som skall sitta på min herre konungens tron efter honom?»
Då svarade konung David och sade: »Kallen hit till mig Bat-Seba.»
När hon nu kom inför konungen och stod inför konungen,
betygade konungen med ed och sade: »Så sant HERREN lever, han som har förlossat mig från all nöd:
såsom jag lovade dig med ed vid HERREN, Israels Gud, då jag sade: 'Din son Salomo skall bliva konung efter mig; han skall sitta på min tron i mitt ställe', så vill jag denna dag göra.»
Då bugade sig Bat-Seba, med ansiktet mot jorden, och föll ned för konungen och sade: »Må min herre, konung David, leva evinnerligen!»
Och konung David sade: »Kallen till mig prästen Sadok och profeten Natan och Benaja, Jojadas son.
När dessa kommo inför konungen,
sade konungen till dem: »Tagen eder herres tjänare med eder och sätten min son Salomo på min egen mulåsna och fören honom med till Gihon.
Där må prästen Sadok och profeten Natan smörja honom till konung över Israel; sedan skolen I stöta i basun och ropa: 'Leve konung Salomo!'
Därefter skolen I följa honom hitupp, och när han kommer hit, skall han sätta sig på min tron, och så skall han vara konung i mitt ställe.
Ty det är honom jag har förordnat att vara furste över Israel och Juda.»
Då svarade Benaja, Jojadas son, konungen och sade: »Amen.
Så bjude ock HERREN, min herre konungens Gud.
Såsom HERREN har varit med min herre konungen, så vare han ock med Salomo.
Ja, må han göra hans tron ännu mäktigare än min herres, konung Davids, tron.»
Så gingo nu prästen Sadok och profeten Natan och Benaja, Jojadas son, ditned, jämte keretéerna och peletéerna, och satte Salomo på konung Davids mulåsna och förde honom till Gihon.
Och prästen Sadok tog oljehornet ur tältet och smorde Salomo.
Därefter stötte de i basun, och allt folket ropade: »Leve konung Salomo!»
Sedan följde allt folket honom upp, under det att de blåste på flöjter och visade sin glädje med ett så stort jubel, att jorden kunde rämna av deras rop.
Men Adonia och alla de inbjudna som han hade hos sig hörde detta, just då de hade slutat att äta.
När Joab nu hörde basunljudet, sade han: »Varför höres detta larm från staden?»
Medan han ännu talade, kom Jonatan, prästen Ebjatars son; och Adonia sade: »Kom hit, ty du är en rättskaffens man och har nog ett gott glädjebudskap att förkunna.»
Jonatan svarade och sade till Adonia: »Nej, vår herre, konung David, har gjort Salomo till konung.
Och konungen har med honom sänt åstad prästen Sadok och profeten Natan och Benaja, Jojadas son, jämte keretéerna och peletéerna, och de hava satt honom på konungens mulåsna.
Därefter hava prästen Sadok och profeten Natan i Gihon smort honom till konung, och sedan hava de dragit upp därifrån under jubel, och hela staden har kommit i rörelse.
Härav kommer det buller som I haven hört.
Salomo sitter nu ock på konungatronen.
Vidare hava konungens tjänare kommit och lyckönskat vår herre konung David, och sagt: 'Din Gud låte Salomos namn bliva ännu större än ditt namn, och hans tron ännu mäktigare än din tron.'
Och konungen har tillbett, nedböjd på sin säng;
ja, konungen har sagt så: 'Lovas vare HERREN, Israels Gud, som i dag har satt en efterträdare på min tron, så att jag med egna ögon har fått se det!»
Då blevo alla de inbjudna som voro hos Adonia förskräckta och stodo upp och gingo bort, var och en sin väg.
Men Adonia fruktade så för Salomo, att han stod upp och gick bort och fattade i hornen på altaret.
Och det blev berättat för Salomo: »Se, Adonia fruktar för konung Salomo; därför har han fattat i hornen på altaret och sagt: 'Konung Salomo måste lova mig i dag med ed att han icke skall döda sin tjänare med svärd.'»
Då sade Salomo: »Om han vill vara en rättskaffens man, så skall icke ett hår av hans huvud falla till jorden; men om något ont bliver funnet hos honom, så skall han dö.»
Därefter sände konung Salomo åstad och lät hämta honom från altaret; och han kom och föll ned för konung Salomo.
Då sade Salomo till honom: »Gå hem till ditt.»
Då nu tiden tillstundade att David skulle dö, bjöd han sin son Salomo och sade:
»Jag går nu all världens väg; så var då frimodig och visa dig såsom en man.
Och håll vad HERREN, din Gud, bjuder dig hålla, så att du vandrar på hans vägar och håller hans stadgar, hans bud och rätter och vittnesbörd, såsom det är skrivet i Moses lag, på det att du må hava framgång i allt vad du gör, och överallt dit du vänder dig;
så att HERREN får uppfylla det ord som han talade om mig, då han sade: 'Om dina barn hava akt på sin väg, så att de vandra inför mig i trohet och av allt sitt hjärta och av all sin själ, då' -- sade han -- 'skall på Israels tron aldrig saknas en avkomling av dig.'
Vidare: du vet väl vad Joab, Serujas son, har gjort mot mig, huru han gjorde mot de två härhövitsmännen i Israel, Abner, Ners son, och Amasa, Jeters son, huru han dräpte dem, så att han i fredstid utgöt blod, likasom hade det varit krig, och, likasom hade det varit krig, lät blod komma på bältet som han hade omkring sina länder, och på skorna som han hade på sina fötter.
Så gör nu efter din vishet, och låt icke hans grå hår få med frid fara ned i dödsriket.
Men mot gileaditen Barsillais söner skall du bevisa godhet, så att de få vara med bland dem som äta vid ditt bord; ty på sådant sätt bemötte de mig, när jag flydde för din broder Absalom.
Vidare har du hos dig Simei, Geras son, benjaminiten från Bahurim, som for ut mot mig i gruvliga förbannelser på den dag då jag gick till Mahanaim, men som sedan kom ned till Jordan mig till mötes, varvid jag med en ed vid HERREN lovade honom och sade: 'Jag skall icke döda dig med svärd.'
Men nu må du icke låta honom bliva ostraffad, ty du är en vis man och vet väl vad du bör göra med honom, så att du låter hans grå hår med blod fara ned i dödsriket.»
och David gick till vila hos sina fäder och blev begraven i Davids stad.
Den tid David regerade över Israel var fyrtio år; i Hebron regerade han i sju år, och i Jerusalem regerade han i trettiotre år.
Och Salomo satte sig på sin fader Davids tron, och han konungamakt blev starkt befäst.
Men Adonia, Haggits son, kom till Bat-Seba, Salomos moder.
Hon frågade då: »Har du gott att meddela?»
Han svarade: »Ja.»
Därefter sade han: »Jag har något att tala med dig om.»
Hon svarade: »Tala.»
Då sade han: »Du vet själv att konungadömet tillhörde mig, och att hela Israel fäste sina blickar på mig, i förväntan att jag skulle bliva konung.
Men så gick konungadömet ifrån mig och blev min broders; genom HERRENS skickelse blev det hans.
Nu har jag en enda bön till dig.
Visa icke bort mig.»
Hon svarade honom: »Tala.»
Då sade han: »Säg till konung Salomo -- dig visar han ju icke bort -- att han giver mig Abisag från Sunem till hustru.»
Bat-Seba svarade: »Gott!
Jag skall själv tala med konungen om dig.»
Så gick då Bat-Seba in till konung Salomo för att tala med honom om Adonia.
Då stod konungen upp och gick emot henne och bugade sig för henne och satte sig därefter på sin stol; man ställde ock fram en stol åt konungens moder, och hon satte sig på hans högra sida.
Därefter sade hon: »Jag har en enda liten bön till dig.
Visa icke bort mig.»
Konungen svarade henne: »Framställ din bön, min moder; jag vill ingalunda visa bort dig.»
Då sade hon: »Låt giva Abisag från Sunem åt din broder Adonia till hustru.»
Men konung Salomo svarade och sade till sin moder: »Varför begär du endast Abisag från Sunem åt Adonia?
Du kunde lika gärna begära konungadömet åt honom -- han är ju min äldste broder -- ja, åt honom och åt prästen Ebjatar och åt Joab, Serujas son.»
Och konung Salomo betygade med ed vid HERREN och sade: »Gud straffe mig nu och framgent, om icke Adonia med sitt liv skall få umgälla att han har talat detta.
Och nu, så sant HERREN lever, han som har utsett mig och uppsatt mig på min fader Davids tron, och som, enligt sitt löfte, har uppbyggt åt mig ett hus: i dag skall Adonia dödas.»
Därefter sände konung Salomo åstad och lät utföra detta genom Benaja, Jojadas son; denne stötte ned honom, så att han dog.
Och till prästen Ebjatar sade konungen: »Gå bort till ditt jordagods i Anatot, ty du har förtjänat döden; men i dag vill jag icke döda dig, eftersom du har burit Herrens, HERRENS ark framför min fader David, och eftersom du med min fader har lidit allt vad han har fått lida.
Så drev Salomo bort Ebjatar och lät honom icke längre vara HERRENS präst, för att HERRENS ord skulle uppfyllas, det som han hade talat i Silo över Elis hus.
Då nu ryktet härom kom till Joab -- som ju hade slutit sig till Adonia, om han ock icke hade slutit sig till Absalom -- flydde han till HERRENS tält och fattade i hornen på altaret.
Men när det blev berättat för konung Salomo att Joab hade flytt till HERRENS tält, och att han stod invid altaret, sände Salomo åstad Benaja, Jojadas son, och sade: »Gå och stöt ned honom.»
När Benaja så kom till HERRENS tält, sade han till honom: »Så säger konungen: Gå bort härifrån.»
Men han svarade: »Nej; här vill jag dö.»
När Benaja framförde detta till konungen och sade: »Så och så har Joab sagt, så har han svarat mig»,
sade konungen till honom: »Gör såsom han har sagt, stöt ned honom och begrav honom, så att du befriar mig och min faders hus från skulden för det blod som Joab utan sak har utgjutit.
Och må HERREN låta hans blod komma tillbaka över hans eget huvud, därför att han stötte ned två män som voro rättfärdigare och bättre än han själv, och dräpte dem med svärd, utan att min fader David visste det, nämligen Abner, Ners son, härhövitsmannen i Israel, och Amasa, Jeters son, härhövitsmannen i Juda.
Ja, deras blod skall komma tillbaka över Joabs och hans efterkommandes huvud för evigt.
Men åt David och hans efterkommande, hans hus och hans tron skall HERREN giva frid till evig tid.
Så gick då Benaja, Jojadas son, ditupp och stötte ned honom och dödade honom; och han blev begraven där han bodde i öknen.
Och konungen satte Benaja, Jojadas son, i hans ställe över hären; och prästen Sadok hade konungen satt i Ebjatars ställe.
Därefter sände konungen och lät kalla till sig Simei och sade till honom: »Bygg dig ett hus i Jerusalem och bo där, och därifrån får du icke gå ut, varken hit eller dit.
Ty det må du veta, att på den dag du går ut och går över bäcken Kidron skall du döden dö.
Ditt blod kommer då över ditt eget huvud.»
Simei sade till konungen: »Vad du har talat är gott; såsom min herre konungen har sagt, så skall din tjänare göra.»
Och Simei bodde i Jerusalem en lång tid.
Men tre år därefter hände sig att två tjänare flydde ifrån Simei till Akis, Maakas son, konungen i Gat.
Och man berättade för Simei och sade: »Dina tjänare äro i Gat.»
Då stod Simei upp och sadlade sin åsna och begav sig till Akis i Gat för att söka efter sina tjänare.
Simei begav sig alltså åstad och hämtade sina tjänare från Gat.
Men när det blev berättat för Salomo att Simei hade begivit sig från Jerusalem till Gat och kommit tillbaka,
sände konungen och lät kalla till sig Simei och sade till honom: »Har jag icke bundit dig med ed vid HERREN och varnat dig och sagt till dig: 'Det må du veta, att på den dag du går ut och begiver dig hit eller dit skall du döden dö'?
Och du svarade mig: 'Vad du har sagt är gott, och jag har hört det.'
Varför har du då icke aktat på din ed vid HERREN och på det bud som jag har givit dig?»
Och konungen sade ytterligare till Simei: »Du känner själv allt det onda som ditt hjärta vet med sig att du har gjort min fader David.
HERREN skall nu låta din ondska komma tillbaka över ditt eget huvud.
Men konung Salomo skall bliva välsignad, och Davids tron skall bliva befäst inför HERREN till evig tid.»
På konungens befallning gick därefter Benaja, Jojadas son, fram och stötte ned honom, så att han dog.
Och konungadömet blev befäst i Salomos hand.
Och Salomo befryndade sig med Farao, konungen i Egypten; han tog Faraos dotter till hustru och förde henne in i Davids stad, och där fick hon bo, till dess han hade byggt sitt hus färdigt, så ock HERRENS hus och muren runt omkring Jerusalem.
Emellertid offrade folket på höjderna, eftersom ännu vid denna tid intet hus hade blivit byggt åt HERRENS namn.
Och Salomo älskade HERREN och vandrade efter sin fader Davids stadgar, utom att han frambar offer på höjderna och tände offereld där.
Och konungen begav sig till Gibeon för att offra där, ty detta var den förnämsta offerhöjden; tusen brännoffer offrade Salomo på altaret där.
I Gibeon uppenbarade sig nu HERREN för Salomo i en dröm om natten; Gud sade: »Bed mig om vad du vill att jag skall giva dig.»
Salomo svarade: »Du har gjort stor nåd med din tjänare, min fader David, eftersom han vandrade inför dig i trohet, rättfärdighet och rättsinnighet mot dig.
Och du bevarade åt honom denna stora nåd och gav honom en son till efterträdare på hans tron, såsom ju nu har skett.
Ja, nu har du, HERRE, min Gud, gjort din tjänare till konung efter min fader David; men jag är en helt ung man, som icke rätt förstår att vara ledare och anförare.
Och din tjänare är här bland ditt folk, det som du har utvalt, ett folk som är så talrikt att det icke kan räknas eller täljas för sin myckenhets skull.
Så giv nu din tjänare ett hörsamt hjärta, så att han kan vara domare för ditt folk och skilja mellan gott och ont; ty vem förmår väl eljest att vara domare för detta ditt stora folk?»
Detta, att Salomo bad om sådant, täcktes Herren.
Och Gud sade till honom: »Eftersom du har bett om sådant och icke bett om ett långt liv, ej heller bett om rikedom eller bett om dina fienders liv, utan har bett om att få förstånd till att akta på vad rätt är,
se, därför vill jag göra såsom du önskar; se, jag giver dig ett så vist och förståndigt hjärta, att din like icke har funnits före dig, och att din like ej heller skall uppstå efter dig.
Därtill giver jag dig ock vad du icke har bett om, nämligen både rikedom och ära, så att i all din tid ingen konung skall vara din like.
Och om du vandrar på mina vägar, så att du håller mina stadgar och bud, såsom din fader David gjorde, då skall jag låta dig länge leva.»
Därefter vaknade Salomo och fann att det var en dröm.
Och när han kom till Jerusalem, trädde han fram inför Herrens förbundsark och offrade brännoffer och frambar tackoffer; och därefter gjorde han ett gästabud för alla sina tjänare.
Vid den tiden kommo två skökor till konungen och trädde fram inför honom.
Och den ena kvinnan sade: »Hör mig, herre.
Jag och denna kvinna bo i samma hus.
Och jag födde barn där i huset hos henne.
Sedan, på tredje dagen efter det jag hade fött mitt barn, födde ock denna kvinna ett barn.
Och vi voro tillsammans, utan att någon främmande var hos oss i huset; allenast vi båda voro i huset.
Men en natt dog denna kvinnas son, ty hon hade legat ihjäl honom.
Då stod hon upp om natten och tog min son från min sida, under det att din tjänarinna sov, och lade honom i sin famn, men sin döde son lade hon i min famn.
När jag då om morgonen reste mig upp för att giva min son di, fick jag se att han var död.
Men när jag såg nogare på honom om morgonen, fick jag se att det icke var min son, den som jag hade fött.»
Då sade den andra kvinnan: »Det är icke så.
Min son är den som lever, och din son är den som är död.»
Men den första svarade: »Det är icke så.
Din son är den som är död, och min son är den som lever.»
Så tvistade de inför konungen.
Då sade konungen: »Den ena säger: 'Denne, den som lever, är min son, och din son är den som är död.'
Och den andra säger: 'Det är icke så.
Din son är den som är död, och min son är den som lever.'»
Därefter sade konungen: »Tagen hit ett svärd.»
Och när man hade burit svärdet fram till konungen,
sade konungen: »Huggen det levande barnet i två delar, och given den ena hälften åt den ena och den andra hälften åt den andra.»
Men då sade den kvinna vilkens son det levande barnet var till konungen -- ty hennes hjärta upprördes av kärlek till sonen -- hon sade: »Hör mig, herre; given henne det levande barnet; döden det icke.»
Men den andra sade: »Må det vara varken mitt eller ditt; huggen det itu.»
Då tog konungen till orda och sade: »Given henne det levande barnet; döden det icke.
Hon är dess moder.»
När nu hela Israel fick höra talas om den dom som konungen hade fällt, häpnade de över konungen, ty de sågo att Guds vishet var i honom till att skipa rätt.
Konung Salomo var nu konung över hela Israel.
Och dessa voro hans förnämsta män: Asarja, Sadoks son, var präst;
Elihoref och Ahia, Sisas söner, voro sekreterare; Josafat, Ahiluds son, var kansler;
Benaja, Jojadas son, var överbefälhavare; Sadok och Ebjatar voro präster;
Asarja, Natans son, var överfogde; Sabud, Natans son, en präst, var konungens vän;
Ahisar var överhovmästare; Adoniram, Abdas son, hade uppsikten över de allmänna arbetena.
Och Salomo hade satt över hela Israel tolv fogdar, som skulle sörja för vad konungen och hans hus behövde; var och en hade årligen sin månad, då han skulle sörja för dessa behov.
Och följande voro deras namn: Ben-Hur i Efraims bergsbygd;
Ben-Deker i Makas, Saalbim, Bet-Semes, Elon, Bet-Hanan;
Ben-Hesed i Arubbot, vilken hade Soko och hela Heferlandet;
Ben-Abinadab i hela Nafat-Dor -- denne fick Salomos dotter Tafat till hustru --;
Baana, Ahiluds son, i Taanak och Megiddo och i hela den del av Bet-Sean, som ligger på sidan om Saretan, nedanför Jisreel, från Bet-Sean ända till Abel-Mehola och bortom Jokmeam;
Ben-Geber i Ramot i Gilead; han hade Manasses son Jairs byar, som ligga i Gilead; han hade ock landsträckan Argob, som ligger i Basan, sextio stora städer med murar och kopparbommar;
Ahinadab, Iddos son, i Mahanaim;
Ahimaas i Naftali; också han hade tagit en dotter av Salomo, Basemat, till hustru;
Baana, Husais son, i Aser och Alot;
Josafat, Paruas son, i Isaskar;
Simei, Elas son, i Benjamin;
Geber, Uris son, i Gileads land, det land som hade tillhört Sihon, amoréernas konung, och Og, konungen i Basan; ty allenast en enda fogde fanns i det landet.
Juda och Israel voro då talrika, så talrika som sanden vid havet; och man åt och drack och var glad.
Så var nu Salomo herre över alla riken ifrån floden till filistéernas land och ända ned till Egyptens gräns; de förde skänker till Salomo och voro honom underdåniga, så länge han levde.
Och vad Salomo för var dag behövde av livsmedel var: trettio korer fint mjöl och sextio korer vanligt mjöl,
tio gödda oxar, tjugu valloxar och hundra far, förutom hjortar, gaseller, dovhjortar och gödda fåglar.
Ty han rådde över hela landet på andra sidan floden, ifrån Tifsa ända till Gasa, över alla konungar på andra sidan floden; och han hade fred på alla sidor, runt omkring,
Så att Juda och Israel sutto i trygghet, var och en under sitt vinträd och sitt fikonträd, ifrån Dan ända till Beer-Seba, så länge Salomo levde.
Och Salomo hade fyrtio tusen spann vagnshästar och tolv tusen ridhästar.
Och de nämnda fogdarna sörjde var sin månad för konung Salomos behov, och för allas som hade tillträde till konung Salomos bord; de läto intet fattas.
Och kornet och halmen för hästarna och travarna förde de, var och en i sin ordning, till det ställe där han uppehöll sig.
Och Gud gav Salomo vishet och förstånd i mycket rikt mått och så mycken insikt, att den kunde liknas vid sanden på havets strand,
så att Salomos vishet var större än alla österlänningars vishet och all Egyptens vishet.
Han var visare än alla andra människor, visare än esraiten Etan och Heman och Kalkol och Darda, Mahols söner; och ryktet om honom gick ut bland alla folk runt omkring.
Han diktade tre tusen ordspråk, och hans sånger voro ett tusen fem.
Han talade om träden, från cedern på Libanon ända till isopen, som växer fram ur väggen.
Han talade ock om fyrfotadjuren, om fåglarna, om kräldjuren och om fiskarna.
Och från alla folk kom man för att höra Salomos visdom, från alla konungar på jorden, som hade hört talas om hans visdom.
Och Hiram, konungen i Tyrus, sände sina tjänare till Salomo, sedan han hade fått höra att denne hade blivit smord till konung efter sin fader; ty Hiram hade alltid varit Davids vän.
Och Salomo sände till Hiram och lät säga:
»Du vet själv att min fader David icke kunde bygga något hus åt HERRENS, sin Guds, namn, för de krigs skull med vilka fienderna runt omkring ansatte honom, till dess att HERREN lade dem under hans fötter
Men nu har HERREN, min Gud, låtit mig få ro på alla sidor; ingen motståndare finnes, och ingen olycka är på färde.
Därför tänker jag nu på att bygga ett hus åt HERRENS, min Guds, namn, såsom HERREN talade till min fader David, i det han sade: 'Din son, den som jag skall sätta på din tron efter dig, han skall bygga huset åt mitt namn.'
Så bjud nu att man hugger åt mig cedrar på Libanon.
Härvid skola mina tjänare vara dina tjänare behjälpliga; och jag vill giva dig betalning för dina tjänares arbete, alldeles såsom du själv begär.
Ty du vet själv att bland oss icke finnes någon som är så skicklig att hugga virke som sidonierna.»
Då nu Hiram hörde Salomos ord, blev han mycket glad; och han sade: »Lovad vare HERREN i dag, han som har givit David en så vis son till att regera över detta talrika folk!»
Och Hiram sände till Salomo och lät säga: »Jag har hört det budskap du har sänt till mig.
Jag vill göra allt vad du begär i fråga om cederträ och cypressträ.
Mina tjänare skola föra virket från Libanon ned till havet, och jag skall låta lägga det i flottar på havet och föra det till det ställe som du anvisar mig, och lossa det där; men du må själv avhämta det.
Du åter skall göra vad jag begär, nämligen förse mitt hus med livsmedel.»
Så gav då Hirom åt Salomo cederträ och cypressträ, så mycket han begärde.
Men Salomo gav åt Hiram tjugu tusen korer vete, till föda för hans hus, och tjugu korer olja av stötta oliver.
Detta gav Salomo åt Hiram för vart år.
Och HERREN hade givit Salomo vishet, såsom han hade lovat honom.
Och vänskap rådde mellan Hiram och Salomo; och de slöto förbund med varandra.
Och konung Salomo bådade upp arbetsfolk ur hela Israel, och arbetsfolket utgjorde trettio tusen man.
Dessa sände han till Libanon, tio tusen i vår månad, skiftevis, så att de voro en månad på Libanon och två månader hemma; och Adoniram hade uppsikten över de allmänna arbetena.
Och Salomo hade sjuttio tusen män som buro bördor, och åttio tusen som höggo sten i bergen,
förutom de överfogdar som av Salomo voro anställda över arbetet, tre tusen tre hundra, vilka hade befälet över folket som utförde arbetet.
Och på konungens befallning bröto de stora och dyrbara stenar, för att husets grund skulle kunna läggas med huggen sten,
Och Salomos byggningsmän och Hiroms byggningsmän och männen från Gebal höggo och tillredde både det trävirke och de stenar som behövdes till att bygga huset.
I det fyra hundra åttionde året efter Israels barns uttåg ur Egyptens land, i det fjärde året av Salomos regering över Israel, i månaden Siv, det är den andra månaden, begynte han bygga huset åt HERREN.
Huset som konung Salomo byggde åt HERREN var sextio alnar långt, tjugu alnar brett och trettio alnar högt.
Förhuset framför tempelsalen var tjugu alnar långt, framför husets kortsida, och tio alnar brett, där det låg framför huset.
Och han gjorde fönster på huset, slutna fönster, med bjälkramar.
Och runt omkring huset, utmed dess vägg, uppförde han en ytterbyggnad, som gick runt omkring husets väggar, både utmed tempelsalen och utmed koret; och han gjorde däri sidokamrar runt omkring.
Den nedersta våningen i ytterbyggnaden var fem alnar bred, den mellersta sex alnar bred och den tredje sju alnar bred; ty han hade gjort avsatser på huset runt omkring utvändigt, för att icke behöva göra fästhål i husets väggar.
Och när huset uppfördes, byggdes det av sten som hade blivit färdighuggen vid stenbrottet; alltså hördes varken hammare eller yxa eller andra järnverktyg vid huset, när det byggdes.
Dörren till mellersta sidokammaren hade sin plats på husets södra sida, och genom en trappgång kom man upp till den mellersta våningen, och från den mellersta våningen upp till den tredje.
Så byggde han huset och fullbordade det.
Och han panelade huset med inläggningar och med cederplankor i rader.
Och i ytterbyggnaden utmed hela huset byggde han våningarna fem alnar höga; och den var fäst vid huset med cederbjälkar.
Och HERRENS ord kom till Salomo; han sade:
»Med detta hus som du nu bygger skall så ske: om du vandrar efter mina stadgar och gör efter mina rätter och håller alla mina bud och vandrar efter dem, så skall jag på dig uppfylla mitt ord, det som jag talade till din fader David:
jag skall bo mitt ibland Israels barn och skall icke övergiva mitt folk Israel.»
Så byggde nu Salomo huset och fullbordade det.
Han täckte husets väggar invändigt med bräder av cederträ.
Från husets golv ända upp till takbjälkarna överklädde han det med trä invändigt; husets golv överklädde han med bräder av cypressträ.
Och han täckte de tjugu alnarna i det innersta av huset med bräder av cederträ, från golvet ända upp till bjälkarna; så inrättade han rummet därinne åt sig till ett kor: det allraheligaste.
Och fyrtio alnar mätte den del av huset, som utgjorde tempelsalen därframför.
Och innantill hade huset en beläggning av cederträ med utsirningar i form av gurkfrukter och blomsterband; alltsammans var där av cederträ, ingen sten syntes.
Och ett kor inredde han i det inre av huset för att där ställa HERRENS förbundsark.
Och framför koret, som var tjugu alnar långt, tjugu alnar brett och tjugu alnar högt, och som han överdrog med fint guld, satte han ett altare, överklätt med cederträ.
Och Salomo överdrog det inre av huset med fint guld.
Och med kedjor av guld stängde han för koret; och jämväl detta överdrog han med guld.
Alltså överdrog han hela huset med guld, till dess att hela huset var helt och hållet överdraget med guld.
Han överdrog ock med guld hela det altare som hörde till koret.
Och till koret gjorde han två keruber av olivträ.
Den ena av dem var tio alnar hög;
och den kerubens ena vinge var fem alnar, och kerubens andra vinge var ock fem alnar, så att det var tio alnar från den ena vingspetsen till den andra.
Den andra keruben var ock tio alnar.
Båda keruberna hade samma mått och samma form:
den ena keruben var tio alnar hög och likaså den andra keruben.
Och han ställde keruberna i de innersta av huset, och keruberna bredde ut sina vingar, så att den enas ena vinge rörde vid den ena väggen och den andra kerubens ena vinge rörde vid den andra väggen; och mitt i huset rörde deras båda andra vingar vid varandra.
Och han överdrog keruberna med guld.
Och alla husets väggar runt omkring utsirade han med snidverk i form av keruber, palmer och blomsterband; så både i det inre rummet och i det yttre.
Och husets golv överdrog han med guld; så både i det inre rummet och i det yttre.
För ingången till koret gjorde han dörrar av olivträ.
Dörrinfattningen hade formen av en femkant.
Och de båda dörrarna av olivträ prydde han med utsirningar i form av keruber, palmer och blomsterband, och överdrog dem med guld; han lade ut guldet över keruberna och palmerna.
Likaså gjorde han för ingången till tempelsalen dörrposter av olivträ, i fyrkant,
och två dörrar av cypressträ, var dörr bestående av två dörrhalvor som kunde vridas.
Och han utsirade dem med keruber, palmer och blomsterband, och överdrog dem med guld, som lades jämnt över snidverken.
Vidare byggde han den inre förgårdsmuren av tre varv huggna stenar och ett varv huggna bjälkar av cederträ.
I det fjärde året blev grunden lagd till HERRENS hus, i månaden Siv.
Och i det elfte året, månaden Bul, det är den åttonde månaden, var huset färdigt till alla sina delar alldeles såsom det skulle vara.
Han byggde alltså därpå i sju år.
Men på sitt eget hus byggde Salomo i tretton år, innan han fick hela sitt hus färdigt.
Han byggde Libanonskogshuset, hundra alnar långt, femtio alnar brett och trettio alnar högt, med fyra rader pelare av cederträ och med huggna bjälkar av cederträ ovanpå pelarna.
Det hade ock ett tak av cederträ över sidokamrarna, vilka vilade på pelarna, som tillsammans voro fyrtiofem, femton i var rad.
Och det hade bjälklag i tre rader; och fönsteröppningarna sutto mitt emot varandra i tre omgångar.
Alla dörröppningar och dörrposter voro fyrkantiga, av bjälkar; och fönsteröppningarna sutto alldeles mitt emot varandra i tre omgångar.
Vidare gjorde han pelarförhuset, femtio alnar långt och trettio alnar brett, och framför detta också ett förhus med pelare, och med ett trapphus framför dessa.
Och han gjorde tronförhuset, där han skulle skipa rätt, domsförhuset; det var belagt med cederträ från golv till tak.
Och hans eget hus, där han själv skulle bo, på den andra gården, innanför förhuset, var byggt på samma sätt.
Salomo byggde ock ett hus, likadant som detta förhus, åt Faraos dotter, som han hade tagit till hustru.
Allt detta var av dyrbara stenar, avmätta såsom byggnadsblock och sågade med såg invändigt och utvändigt, alltsammans, ända ifrån grunden upp till taklisterna; och likaså allt därutanför, ända till den stora förgårdsmuren.
Och grunden var lagd med dyrbara och stora stenar, stenar av tio alnars längd och av åtta alnars längd.
Därovanpå lågo dyrbara stenar, avmätta såsom byggnadsblock, ävensom cederbjälkar.
Och den stora förgårdsmuren där runt omkring var uppförd av tre varv huggna stenar och ett varv huggna bjälkar av cederträ.
Så var det ock med den inre förgårdsmuren till HERRENS hus, så jämväl med husets förhus.
Och konung Salomo sände och lät hämta Hiram från Tyrus.
Denne var son till en änka av Naftali stam, och hans fader var en tyrisk man, en kopparsmed; han hade konstskicklighet och förstånd och kunskap i fullt mått till att utföra alla slags arbeten av koppar.
Han kom nu till konung Salomo och utförde alla hans arbeten.
Han förfärdigade de båda pelarna av koppar.
Aderton alnar hög var den ena pelaren, och en tolv alnar lång tråd mätte omfånget av den andra pelaren.
Han gjorde ock två pelarhuvuden, gjutna av koppar, till att sätta ovanpå pelarna; vart pelarhuvud var fem alnar högt.
Nätlika utsirningar, som bildade ett nätverk, hängprydnader i form av kedjor funnos på pelarhuvudena som sutto ovanpå pelarna, sju på vart pelarhuvud.
Och han gjorde pelarna så, att två rader gingo runt omkring över det ena av de nätverk som tjänade till att betäcka pelarhuvudena, vilka höjde sig över granatäpplena; och likadant gjorde han på det andra pelarhuvudet.
Och pelarhuvudena som sutto ovanpå pelarna inne i förhuset voro utformade till liljor, och mätte fyra alnar.
På båda pelarna funnos pelarhuvuden, också ovantill invid den bukformiga delen inemot nätverket.
Och granatäpplena voro två hundra, i rader runt omkring, över det andra pelarhuvudet.
Pelarna ställde han upp vid förhuset till tempelsalen.
Åt den pelare han ställde upp på högra sidan gav han namnet Jakin, och åt den han ställde upp på vänstra sidan gav han namnet Boas.
Överst voro pelarna utformade till liljor.
Så blev då arbetet med pelarna fullbordat.
Han gjorde ock havet, i gjutet arbete.
Det var tio alnar från den ena kanten till den andra, runt allt omkring, och fem alnar högt; och ett trettio alnar långt snöre mätte dess omfång.
Och under kanten voro gurklika sirater, som omgåvo det runt omkring -- tio alnar brett som det var -- så att de gingo runt omkring havet.
De gurklika siraterna sutto i två rader, och de voro gjutna i ett stycke med det övriga.
Det stod på tolv oxar, tre vända mot norr, tre vända mot väster, tre vända mot söder och tre vända mot öster; havet stod ovanpå dessa, och deras bakdelar voro alla vända inåt.
Dess tjocklek var en handsbredd; och dess kant var gjord såsom kanten på en bägare, i form av en utslagen lilja.
Det rymde två tusen bat.
Vidare gjorde han de tio bäckenställen, av koppar.
Vart ställ var fyra alnar långt, fyra alnar brett och tre alnar högt.
Och på följande sätt voro dessa ställ gjorda.
De voro försedda med sidolister, vilka sidolister hade sin plats mellan hörnlisterna.
På dessa sidolister mellan hörnlisterna funnos avbildade lejon, tjurar och keruber, och likaså på hörnlisterna upptill.
Under lejonen och tjurarna sutto nedhängande blomsterslingor.
Vart ställ hade fyra hjul av koppar med axlar av koppar; och dess fyra fötter voro försedda med bärarmar.
Dessa bärarmar voro gjutna till att sitta under bäckenet, och mitt för var och en sutto blomsterslingor.
Sin öppning hade det inom kransstycket, som höjde sig en aln uppåt. öppningen i detta var rund; det var så gjort, att det kunde tjäna såsom underlag, och det mätte en och en halv aln.
Också på dess öppning funnos utsirningar.
Men sidolisterna därtill voro fyrkantiga, icke runda.
De fyra hjulen sutto under sidolisterna, och hjulens hållare voro fästa vid bäckenstället.
Vart hjul mätte en och en halv aln.
Hjulen voro gjorda såsom vagnshjul; och deras hållare, deras ringar, deras ekrar och deras navar voro allasammans gjutna.
Fyra bärarmar funnos på vart ställ, i de fyra hörnen; bärarmarna voro gjorda i ett stycke med sitt ställ.
Överst på vart ställ var en helt och hållet rund uppsats, en halv aln hög; och ovantill på vart ställ sutto dess hållare, så ock dess sidolister gjorda i ett stycke därmed.
Och på hållarnas ytor och på sidolisterna inristade han keruber, lejon och palmer, alltefter som utrymme fanns på var och en, så ock blomsterslingor runt omkring.
På detta sätt gjorde han de tio bäckenställen; de voro alla gjutna på samma sätt och hade samma mått och samma form
Han gjorde ock tio bäcken, av koppar.
Fyrtio bat rymde vart bäcken, och vart bäcken mätte fyra alnar; till vart och ett av de tio bäckenställen gjordes ett bäcken.
Och han ställde fem av bäckenställen på högra sidan om huset och fem på vänstra sidan om huset.
Och havet ställde han på högra sidan om huset, åt sydost.
Hirom gjorde dessa bäcken, så ock skovlarna och skålarna.
Så förde Hiram allt det arbete till slut, som han fick utföra åt konung Salomo för HERRENS hus:
nämligen två pelare, och de två klotformiga pelarhuvuden som sutto ovanpå pelarna, och de två nätverk som skulle betäcka de båda klotformiga pelarhuvuden som sutto ovanpå pelarna,
därjämte de fyra hundra granatäpplena till de båda nätverken, två rader granatäpplen till vart nätverk, för att de båda klotformiga pelarhuvuden som sutto uppe på pelarna så skulle bliva betäckta,
Vidare de tio bäckenställen och de tio bäckenen på bäckenställen,
så ock havet, som var allenast ett, och de tolv oxarna under havet,
vidare askkärlen, skovlarna och skålarna, korteligen, alla redan nämnda föremål som Hiram gjorde åt konung Salomo för HERRENS hus.
Allt var av polerad koppar.
På Jordanslätten lät konungen gjuta det i lerformar, mellan Suckot och Saretan.
Och för den övermåttan stora myckenhetens skull lämnade Salomo alla föremålen ovägda, så att kopparens vikt icke blev utrönt.
Salomo gjorde ock alla övriga föremål som skulle finnas i HERRENS hus: det gyllene altaret, det gyllene bordet som skådebröden skulle ligga på,
så ock ljusstakarna, fem på högra sidan och fem på vänstra framför koret, av fint guld, med blomverket, lamporna och lamptängerna av guld,
vidare faten, knivarna, de båda slagen av skålar och fyrfaten, av fint guld, äntligen de gyllene gångjärnen till de dörrar som ledde till det innersta av huset, det allraheligaste, och till de dörrar i huset, som ledde till tempelsalen.
Sedan allt det arbete som konung Salomo lät utföra på HERRENS hus var färdigt, förde Salomo ditin vad hans fader David hade helgat åt HERREN: silvret, guldet och kärlen; detta lade han in i skattkamrarna i HERRENS hus.
Därefter församlade Salomo de äldste i Israel, alla huvudmännen för stammarna, Israels barns familjehövdingar, till konung Salomo i Jerusalem, för att hämta HERRENS förbundsark upp från Davids stad, det är Sion.
Så församlade sig då till konung Salomo alla Israels män under högtiden i månaden Etanim, det är den sjunde månaden.
När då alla de äldste i Israel hade kommit tillstädes, lyfte prästerna upp arken.
Och de hämtade HERRENS ark och uppenbarelsetältet ditupp, jämte alla heliga föremål som funnos i tältet; prästerna och leviterna hämtade det ditupp.
Och konung Salomo stod framför arken jämte Israels hela menighet, som hade församlats till honom; och de offrade därvid småboskap och fäkreatur i sådan myckenhet, att de icke kunde täljas eller räknas.
Och prästerna buro in HERRENS förbundsark till dess plats i husets kor, i det allraheligaste, till platsen under kerubernas vingar.
Ty keruberna bredde ut sina vingar fram över den plats där arken stod, så att arken och dess stänger ovantill betäcktes av keruberna.
Och stängerna voro så långa, att deras ändar väl kunde ses från helgedomen framför koret, men däremot icke voro synliga längre ute.
Och de hava blivit kvar där ända till denna dag.
I arken fanns intet annat än de två stentavlor som Mose hade lagt ned däri vid Horeb, när HERREN slöt förbund med Israels barn, sedan de hade dragit ut ur Egyptens land.
Men när prästerna gingo ut ur helgedomen, uppfyllde molnskyn HERRENS hus,
så att prästerna för molnskyns skull icke kunde stå där och göra tjänst; ty HERRENS härlighet uppfyllde HERRENS hus.
Då sade Salomo: »HERREN har sagt att han vill bo i töcknet.
Jag har nu byggt ett hus till boning åt dig, berett en plats där du må förbliva till evig tid.»
Sedan vände konungen sig om och välsignade Israels hela församling, under det att Israels hela församling förblev stående.
Han sade: »Lovad vare HERREN, Israels Gud, som med sin hand har fullbordat vad han med sin mun lovade min fader David, i det han sade:
'Från den dag då jag förde mitt folk Israel ut ur Egypten har jag icke i någon av Israels stammar utvalt en stad, till att i den bygga ett hus där mitt namn skulle vara; men David har jag utvalt till att råda över mitt folk Israel.'
Och min fader David hade väl i sinnet att bygga ett hus åt HERRENS, Israels Guds, namn;
men HERREN sade till min fader David: 'Då du nu har i sinnet att bygga ett hus åt mitt namn, så gör du visserligen väl däri att du har detta i sinnet;
dock skall icke du få bygga detta hus, utan din son, den som har utgått från din länd, han skall bygga huset åt mitt namn.'
Och HERREN har uppfyllt det löfte han gav; ty jag har kommit upp min fader Davids ställe och sitter nu på Israels tron, såsom HERREN lovade, och jag har byggt huset åt HERRENS, Israels Guds, namn.
Och där har jag tillrett ett rum för arken, i vilken förvaras det förbund som HERREN slöt med våra fäder, när han förde dem ut ur Egyptens land.»
Därefter trädde Salomo fram för HERRENS altare inför Israels hela församling, och uträckte sina händer mot himmelen
och sade: »HERRE, Israels Gud, ingen gud är dig lik, uppe i himmelen eller nere på jorden, du som håller förbund och bevarar nåd mot dina tjänare, när de vandra inför dig av allt sitt hjärta,
du som har hållit vad du lovade din tjänare David, min fader; ty vad du med din mun lovade, det fullbordade du med din hand, såsom nu har skett.
Så håll nu ock, HERRE, Israels Gud, vad du lovade din tjänare David, min fader, i det att du sade: 'Aldrig skall den tid komma, då på Israels tron icke inför mig sitter en avkomling av dig, om allenast dina barn hava akt på sin väg, så att de vandra inför mig, såsom du har vandrat inför mig.'
Så låt nu, o Israels Gud, de ord som du har talat till din tjänare David, min fader, bliva sanna.
Men kan då Gud verkligen bo på jorden?
Himlarna och himlarnas himmel rymma dig ju icke; huru mycket mindre då detta hus som jag har byggt!
Men vänd dig ändå till din tjänares bön och åkallan, HERRE, min Gud, så att du hör på det rop och den bön som din tjänare nu uppsänder till dig,
och låter dina ögon natt och dag vara öppna och vända mot detta hus -- den plats varom du har sagt: 'Mitt namn skall vara där' -- så att du ock hör den bön som din tjänare beder, vänd mot denna plats.
Ja, hör på den åkallan som din tjänare och ditt folk Israel uppsända, vända mot denna plats.
Må du höra den och låta den komma upp till himmelen, där du bor; och när du hör, så må du förlåta.
Om någon försyndar sig mot sin nästa och man ålägger honom en ed och låter honom svärja, och han så kommer och svär inför ditt altare i detta hus,
må du då höra det i himmelen och utföra ditt verk och skaffa dina tjänare rätt, i det att du dömer den skyldige skyldig och låter hans gärningar komma över hans huvud, men skaffar rätt åt den som har rätt och låter honom få efter hans rättfärdighet.
Om ditt folk Israel bliver slaget av en fiende, därför att de hava syndat mot dig, men de omvända sig till dig och prisa ditt namn och bedja och åkalla dig i detta hus,
må du då höra det i himmelen och förlåta ditt folk Israels synd och låta dem komma tillbaka till det land som du har givit åt deras fäder.
Om himmelen bliver tillsluten, så att regn icke faller, därför att de hava syndat mot dig, men de då bedja, vända mot denna plats, och prisa ditt namn och omvända sig från sin synd, när du bönhör dem,
må du då höra det i himmelen och förlåta dina tjänares och ditt folk Israels synd, i det att du lär dem den goda väg som de skola vandra; och må du låta det regna över ditt land, det som du har givit åt ditt folk till arvedel.
Om hungersnöd uppstår i landet, om pest uppstår, om sot eller rost, om gräshoppor eller gräsmaskar komma, om fienden tränger folket i det land där deras städer stå, eller om någon annan plåga eller sjukdom kommer, vilken det vara må,
och om då någon bön och åkallan höjes från någon människa, vilken det vara må, eller från hela ditt folk Israel, när de var för sig känna plågan därav i sitt hjärta och så uträcka sina händer mot detta hus,
må du då höra det i himmelen, där du bor, och förlåta och utföra ditt verk, i det att du giver var och en efter alla hans gärningar, eftersom du känner hans hjärta -- ty du allena känner alla människors hjärtan --
på det att de alltid må frukta dig, så länge de leva i det land som du har givit åt våra fäder.
Också om en främling, en som icke är av ditt folk Israel, kommer ifrån fjärran land för ditt namns skull
-- ty man skall ock där höra talas om ditt stora namn och din starka hand och din uträckta arm -- om någon sådan kommer och beder, vänd mot detta hus,
må du då i himmelen, där du bor, höra det och göra allt varom främlingen ropar till dig, på det att alla jordens folk må känna ditt namn och frukta dig, likasom ditt folk Israel gör, och förnimma att detta hus som jag har byggt är uppkallat efter ditt namn.
Om ditt folk drager ut i strid mot sin fiende, på den väg du sänder dem, och de då bedja till HERREN, vända i riktning mot den stad som du har utvalt, och mot det hus som jag har byggt åt ditt namn,
må du då i himmelen höra deras bön och åkallan och skaffa dem rätt.
Om de synda mot dig -- eftersom ingen människa finnes, som icke syndar -- och du bliver vred på dem och giver dem i fiendens våld, så att man tager dem till fånga och för dem bort till fiendens land, fjärran eller nära,
men de då besinna sig i det land där de äro i fångenskap, och omvända sig och åkalla dig i landet där man håller dem fångna och säga: 'Vi hava syndat och gjort illa, vi hava varit ogudaktiga',
om de så omvända sig till dig av allt sitt hjärta och av all sin själ, i sina fienders land -- deras som hava fört dem i fångenskap -- och bedja till dig, vända i riktning mot sitt land, det som du har givit åt deras fäder, och mot den stad som du har utvalt, och mot det hus som jag har byggt åt ditt namn,
må du då i himmelen, där du bor, höra deras bön och åkallan och skaffa dem rätt
och förlåta ditt folk vad de hava syndat mot dig, och alla de överträdelser som de hava begått mot dig, och låta dem finna barmhärtighet inför dem som hålla dem fångna, så att dessa förbarma sig över dem.
Ty de äro ju ditt folk och din arvedel, som du har fört ut ur Egypten, den smältugnen.
Ja, låt dina ögon vara öppna och vända till din tjänares och ditt folk Israels åkallan, så att du hör på dem, så ofta de ropa till dig.
Ty du har själv avskilt dem åt dig till arvedel bland alla folk på Jorden, såsom du talade genom din tjänare Mose, när du förde våra fäder ut ur Egypten, o Herre, HERRE.»
När Salomo hade slutat att med dessa ord bedja och åkalla HERREN, stod han upp från HERRENS altare, där han hade legat på sina knän med händerna uträckta mot himmelen,
och trädde fram och välsignade Israels hela församling med hög röst och sade:
»Lovad vare HERREN, som har givit sitt folk Israel ro, alldeles såsom han har sagt!
Alls intet har uteblivit av allt det goda som han lovade genom sin tjänare Mose.
Så vare då HERREN, vår Gud, med oss, såsom han har varit med våra fäder.
Han må icke övergiva oss och förskjuta oss,
utan böja våra hjärtan till sig, så att vi alltid vandra på hans vägar och hålla hans bud och stadgar och rätter, dem som han har givit våra fäder.
Och må dessa mina ord, med vilka jag har bönfallit inför HERRENS ansikte, vara nära HERREN, vår Gud, dag och natt, så att han skaffar rätt åt sin tjänare och rätt åt sitt folk Israel, efter var dags behov;
på det att alla folk på jorden må förnimma att HERREN är Gud, och ingen annan.
Och må edra hjärtan vara hängivna åt HERREN, vår Gud, så att I alltjämt vandren efter hans stadgar och hållen hans bud, såsom I nu gören.»
Och konungen jämte hela Israel offrade slaktoffer inför HERRENS ansikte.
Till det tackoffer som Salomo offrade åt HERREN tog han tjugutvå tusen tjurar och ett hundra tjugu tusen av småboskapen.
Så invigdes HERRENS hus av konungen och alla Israels barn.
På samma dag helgade konungen den mellersta delen av förgården framför HERRENS hus, ty där offrade han brännoffret, spisoffret och fettstyckena av tackoffret, eftersom kopparaltaret, som stod inför HERRENS ansikte, var för litet för att brännoffret, spisoffret och fettstyckena av tackoffret skulle kunna rymmas där.
Vid detta tillfälle firade Salomo högtiden, och med honom hela Israel -- en stor församling ifrån hela landet, allt ifrån det ställe där vägen går till Hamat ända till Egyptens bäck -- inför HERRENS, vår Guds, ansikte i sju dagar och åter sju dagar, tillsammans fjorton dagar.
På åttonde dagen lät han folket gå, och de togo avsked av konungen.
Sedan gingo de till sina hyddor, fulla av glädje och fröjd över allt det goda som HERREN hade gjort mot sin tjänare David och sitt folk Israel.
Då nu Salomo hade byggt HERRENS hus färdigt, så ock konungshuset, ävensom allt annat som han hade känt åstundan och lust att utföra,
uppenbarade sig HERREN för andra gången för Salomo, likasom han förut hade uppenbarat sig för honom i Gibeon.
Och HERREN sade till honom »Jag har hört den bön och åkallan som du har uppsänt till mig; detta hus som du har byggt har jag helgat, till att där fästa mitt namn för evig tid.
Och mina ögon och mitt hjärta skola vara där alltid.
Om du nu vandrar inför mig, såsom din fader David vandrade, med ostraffligt hjärta och i redlighet, så att du gör allt vad jag har bjudit dig och håller mina stadgar och rätter
då skall jag upprätthålla din konungatron över Israel evinnerligen, såsom jag lovade angående din fader David, när jag sade: 'Aldrig skall på Israels tron saknas en avkomling av dig.'
Men om I och edra barn vänden om och övergiven mig, och icke hållen de bud och stadgar som jag har förelagt eder, utan gån bort och tjänen andra gudar och tillbedjen dem,
då skall jag utrota Israel ur det land som jag har givit dem; och det hus som jag har helgat åt mitt namn skall jag förkasta ifrån mitt ansikte; och Israel skall bliva ett ordspråk och en visa bland alla folk.
Och huru upphöjt detta hus nu än må vara, skall då var och en som går därförbi bliva häpen och vissla.
Och när man frågar: 'Varför har HERREN gjort så mot detta land och detta hus?',
då skall man svara: 'Därför att de övergåvo HERREN, sin Gud, som hade fört deras fäder ut ur Egyptens land, och höllo sig till andra gudar och tillbådo dem och tjänade dem, därför har HERREN låtit allt detta onda komma över dem.'»
När de tjugu år voro förlidna, under vilka Salomo byggde på de två husen, HERRENS hus och konungshuset,
gav konung Salomo tjugu städer i Galileen åt Hiram, konungen i Tyrus, som hade försett honom med cederträ, cypressträ och guld, så mycket han begärde.
Men när Hiram från Tyrus begav sig ut för att bese de städer som Salomo hade givit honom, behagade de honom icke,
utan han sade: »Vad är detta för städer som du har givit mig, min broder?»
Och han kallade dem Kabuls land, såsom de heta ännu i dag.
Men Hiram sände till konungen ett hundra tjugu talenter guld.
Och på följande sätt förhöll det sig med det arbetsfolk som konung Salomo bådade upp för att bygga HERRENS hus och hans eget hus och Millo, ävensom Jerusalems murar, så ock Hasor, Megiddo och Geser.
(Farao, konungen i Egypten, hade nämligen dragit upp och intagit Geser och bränt upp det i eld och dräpt de kananéer som bodde i staden, varefter han hade givit den till hemgift åt sin dotter, Salomos hustru.
Men Salomo byggde upp Geser, ävensom Nedre Bet-Horon,
så ock Baalat och Tamar i öknen där i landet,
vidare alla Salomos förrådsstäder, vagnsstäderna och häststäderna, och vad annat Salomo kände åstundan att bygga i Jerusalem, på Libanon och eljest i hela det land som lydde under hans välde.)
Allt det folk som fanns kvar av amoréerna, hetiterna, perisséerna hivéerna och jebuséerna, korteligen, alla de som icke voro av Israels barn --
deras avkomlingar, så många som funnos kvar i landet efter dem, i det Israels barn icke hade förmått giva dem till spillo, dessa pålade Salomo att vara arbetspliktiga tjänare, såsom de äro ännu i dag.
Men av Israels barn gjorde Salomo ingen till träl, utan de blevo krigare och blevo hans tjänare och hövitsman och kämpar, eller uppsyningsmän över hans vagnar och ridhästar.
Överfogdarna över Salomos arbeten voro fem hundra femtio; dessa hade befälet över folket som utförde arbetet.
Men så snart Faraos dotter hade flyttat upp från Davids stad till det hus som han hade byggt åt henne, byggde han ock Millo.
Och Salomo offrade tre gånger om året brännoffer och tackoffer på det altare som han hade byggt åt HERREN, och tände därjämte rökelsen inför HERRENS ansikte.
Så hade han då gjort huset färdigt.
Konung Salomo byggde ock en flotta i Esjon-Geber, som ligger vid Elot, på stranden av Röda havet, i Edoms land.
På denna flotta sände Hiram av sitt folk sjökunnigt skeppsmanskap, som åtföljde Salomos folk.
De foro till Ofir och hämtade därifrån guld, fyra hundra tjugu talenter, som de förde till konung Salomo.
När drottningen av Saba fick höra ryktet om Salomo och vad han hade gjort för HERRENS namn, kom hon för att sätta honom på prov med svåra frågor.
Hon kom till Jerusalem med ett mycket stort följe, med kameler, som buro välluktande kryddor och guld i stor myckenhet, så ock ädla stenar.
Och när hon kom inför Salomo, förelade hon honom allt vad hon hade i tankarna.
Men Salomo gav henne svar på alla hennes frågor; intet var förborgat för konungen, utan han kunde giva henne svar på allt.
När nu drottningen av Saba såg all Salomos vishet, och såg huset som han hade byggt,
och såg rätterna på hans bord, och såg huru hans tjänare sutto där, och huru de som betjänade honom utförde sina åligganden, och huru de voro klädda, och vidare såg hans munskänkar, och när hon såg brännoffren som han offrade i HERRENS hus, då blev hon utom sig av förundran.
Och hon sade till konungen: »Sant var det tal som jag hörde i mitt land om dig och om din vishet.
Jag ville icke tro vad man sade, förrän jag själv kom och med egna ögon fick se det; men nu finner jag att det icke ens till hälften har blivit omtalat för mig.
Du har långt mer vishet och rikedom, än jag genom ryktet hade hört.
Sälla äro dina män, sälla äro dessa dina tjänare, som beständigt få stå inför dig och höra din visdom.
Lovad vare HERREN, din Gud, som har funnit sådant behag i dig, att han har satt dig på Israels tron!
Ja, därför att HERREN älskar Israel evinnerligen, därför har han satt dig till konung, för att du skall skipa lag och rätt.»
Och hon gav åt konungen ett hundra tjugu talenter guld, så ock välluktande kryddor i stor myckenhet, därtill ädla stenar; en så stor myckenhet av välluktande kryddor, som drottningen av Saba gav åt konung Salomo, har aldrig mer blivit införd.
När Hirams flotta hämtade guld från Ofir, hemförde också den från Ofir almugträ i stor myckenhet, ävensom ädla stenar.
Av almugträet lät konungen göra tillbehör till HERRENS hus och till konungshuset, så ock harpor och psaltare för sångarna.
Så mycket almugträ har sedan intill denna dag icke införts eller blivit sett i landet.
Konung Salomo åter gav åt drottningen av Saba allt vad hon åstundade och begärde, och skänkte henne i sin konungsliga frikostighet också annat därutöver.
Sedan vände hon om och for till sitt land igen med sina tjänare.
Det guld som årligen inkom till Salomo vägde sex hundra sextiosex talenter,
förutom det som inkom genom kringresande handelsmän och genom krämares köpenskap, så ock från Erebs alla konungar och från ståthållarna i landet.
Och konung Salomo lät göra två hundra stora sköldar av uthamrat guld och använde till var sådan sköld sex hundra siklar guld;
likaledes tre hundra mindre sköldar av uthamrat guld och använde till var sådan sköld tre minor guld; och konungen satte upp dem i Libanonskogshuset.
Vidare lät konungen göra en stor tron av elfenben och överdrog den med fint guld.
Tronen hade sex trappsteg, och tronens ryggstycke var ovantill avrundat; på båda sidor om sitsen voro armstöd, och två lejon stodo utmed armstöden;
och tolv lejon stodo där på de sex trappstegen, på båda sidor.
Något sådant har aldrig blivit förfärdigat i något annat rike.
Och alla konung Salomos dryckeskärl voro av guld, och alla kärl i Libanonskogshuset voro av fint guld; av silver fanns intet, det aktades icke för något i Salomos tid.
Ty konungen hade en egen Tarsisflotta på havet jämte Hirams flotta; en gång vart tredje år kom Tarsisflottan hem och förde med sig guld och silver, elfenben, apor och påfåglar.
Och konung Salomo blev större än någon annan konung på jorden, både i rikedom och i vishet.
Från alla länder kom man för att besöka Salomo och höra den vishet som Gud hade nedlagt i hans hjärta.
Och var och en förde med sig skänker: föremål av silver och av guld, kläder, vapen, välluktande kryddor, hästar och mulåsnor.
Så skedde år efter år.
Salomo samlade ock vagnar och ridhästar, så att han hade ett tusen fyra hundra vagnar och tolv tusen ridhästar; dem förlade han dels i vagnsstäderna, dels i Jerusalem, hos konungen själv.
Och konungen styrde så, att silver blev lika vanligt i Jerusalem som stenar, och cederträ lika vanligt som mullbärsfikonträ i Låglandet.
Och hästarna som Salomo lät anskaffa infördes från Egypten; ett antal kungliga uppköpare hämtade ett visst antal av dem till bestämt pris.
Var vagn som hämtades upp från Egypten och infördes kostade sex hundra siklar silver, och var häst ett hundra femtio.
Sammalunda infördes ock genom deras försorg sådana till hetiternas alla konungar och till konungarna i Aram.
Men konung Salomo hade utom Faraos dotter många andra utländska kvinnor som han älskade: moabitiskor, ammonitiskor, edomeiskor, sidoniskor och hetitiskor,
kvinnor av de folk om vilka HERREN hade lagt till Israels barn: »I skolen icke inlåta eder med dem, och de få icke inlåta sig med eder; de skola förvisso eljest förleda edra hjärtan att avfalla till deras gudar.»
Till dessa höll sig Salomo och älskade dem.
Han hade sju hundra furstliga gemåler och tre hundra bihustrur.
Dessa kvinnor förledde hans hjärta till avfall.
Ja, när Salomo blev gammal, förledde kvinnorna hans hjärta att avfalla till andra gudar, så att hans hjärta icke förblev hängivet åt HERREN, hans Gud, såsom hans fader Davids hjärta hade varit.
Så kom Salomo att följa efter Astarte, sidoniernas gudinna, och Milkom, ammoniternas styggelse.
Och Salomo gjorde vad ont var i HERRENS ögon och följde icke i allt efter HERREN, såsom hans fader David hade gjort.
Salomo byggde nämligen då en offerhöjd åt Kemos, moabiternas styggelse, på berget öster om Jerusalem, och likaså en åt Molok, Ammons barns styggelse.
På samma sätt gjorde han för alla sina utländska kvinnor, så att de fingo tända offereld och frambära offer åt sina gudar.
Och HERREN blev vred på Salomo, därför att hans hjärta hade avfallit från HERREN, Israels Gud, som dock två gånger hade uppenbarat sig för honom,
och som hade givit honom ett särskilt bud angående denna sak, att han icke skulle följa efter andra gudar, ett HERRENS bud som han icke hade hållit.
Därför sade HERREN till Salomo: »Eftersom det är så med dig, och eftersom du icke har hållit det förbund och de stadgar som jag har givit dig, skall jag rycka riket ifrån dig och giva det åt din tjänare.
Men för din fader Davids skull vill jag icke göra detta i din tid; först ur din sons hand skall jag rycka det.
Dock skall jag icke rycka hela riket ifrån honom, utan en stam skall jag giva åt din son, för min tjänare Davids skull och för Jerusalems skull, som jag har utvalt.»
Och HERREN lät en motståndare till Salomo uppstå i edoméen Hadad.
Denne var av konungasläkten i Edom.
Ty när David var i strid med Edom, och härhövitsmannen Joab drog upp för att begrava de slagna och därvid förgjorde allt mankön i Edom
-- ty Joab och hela Israel stannade där i sex månader, till dess att han hade utrotat allt mankön i Edom --
då flydde Adad jämte några edomeiska män som hade varit i hans faders tjänst, och de togo vägen till Egypten; Hadad var då en ung gosse.
De begav sig åstad från Midjan och kommo till Paran; och de togo folk med sig från Paran och kommo så till Egypten, till Farao, konungen i Egypten.
Denne gav honom ett hus och anslog ett underhåll åt honom och gav honom land.
Och Hadad fann mycken nåd för Faraos ögon, så att denne gav honom till hustru en syster till sin gemål, en syster till drottning Tapenes.
Denna syster till Tapenes födde åt honom sonen Genubat, och Tapenes lät avvänja honom i Faraos hus; sedan vistades Genubat i Faraos hus bland Faraos söner.
Då nu Hadad i Egypten hörde att David hade gått till vila hos sina fäder, och att härhövitsmannen Joab var död, sade han till Farao: »Låt mig fara hem till mitt land.»
Men Farao sade till honom: »Vad fattas dig här hos mig, eftersom du vill fara till ditt land?»
Han svarade: »Hindra mig icke, utan låt mig gå.
Och Gud lät ännu en motståndare till honom uppstå i Reson, Eljadas son, som hade flytt ifrån sin herre, Hadadeser, konungen i Soba.
När David sedan anställde blodbadet ibland dem, samlade denne folk omkring sig och blev hövitsman för en strövskara; dessa drogo därefter till Damaskus och slogo sig ned där och gjorde sig till herrar i Damaskus.
Denne var nu under Salomos hela livstid Israels motståndare och gjorde det skada, han såväl som Hadad.
Han avskydde Israel; och han blev konung över Aram.
Och en av Salomos tjänare hette Jerobeam; han var son till Nebat, en efraimit, från Sereda, och hans moder hette Seruga och var änka.
Denne reste sig upp mot konungen.
Orsaken varför han reste sig upp mot konungen var följande.
Salomo byggde då på Millo; han ville befästa det blottade stället på sin fader Davids stad.
Nu var Jerobeam en dugande man; och då Salomo såg att den unge mannen var driftig i sitt arbete, satte han honom över allt det arbete som ålåg Josefs hus.
Vid den tiden hände sig en gång att Jerobeam hade begivit sig ut ur Jerusalem; då kom profeten Ahia från Silo emot honom på vägen, där han gick klädd i en ny mantel; och de båda voro ensamma på fältet.
Och Ahia fattade i den nya manteln som han hade på sig och ryckte sönder den i tolv stycken.
Därefter sade han till Jerobeam: »Tag här tio stycken för dig.
Ty så säger HERREN, Israels Gud: Se, jag vill rycka riket ur Salomos hand och giva tio av stammarna åt dig;
den ena stammen skall han få behålla för min tjänare Davids skull och för Jerusalems skull, den stads som jag har utvalt ur alla Israels stammar.
Så skall ske, därför att de hava övergivit mig och tillbett Astarte, sidoniernas gudinna, och Kemos, Moabs gud, och Milkom, Ammons barns gud, och icke vandrat på mina vägar och icke gjort vad rätt är i mina ögon, efter mina stadgar och rätter, såsom hans fader David gjorde.
Dock skall jag icke taga ifrån honom själv det samlade riket, utan jag vill låta honom förbliva furste, så länge han lever, för min tjänare Davids skull, som jag utvalde, därför att han höll mina bud och stadgar.
Men från hans son skall jag taga konungadömet och giva det åt dig, nämligen de tio stammarna.
En stam skall jag giva åt hans son, så att min tjänare David alltid har en lampa inför mitt ansikte i Jerusalem, den stad som jag har utvalt åt mig, till att där fästa mitt namn.
Dig vill jag alltså taga och vill låta dig regera över allt vad dig lyster; du skall bliva konung över Israel.
Om du nu hörsammar allt vad jag bjuder dig och vandrar på mina vägar och gör vad rätt är i mina ögon, så att du håller mina stadgar och bud, såsom min tjänare David gjorde, så skall jag vara med dig och bygga åt dig ett hus som bliver beståndande, såsom jag byggde ett hus åt David, och jag skall giva Israel åt dig. --
Ja, för den sakens skull skall jag ödmjuka Davids säd, dock icke för alltid.»
Och Salomo sökte tillfälle att döda Jerobeam; men Jerobeam stod upp och flydde till Egypten, till Sisak, konungen i Egypten.
Och han stannade i Egypten till Salomos död.
Vad nu mer är att säga om Salomo, om allt vad han gjorde och om hans vishet, det finnes upptecknat i Salomos krönika.
Den tid Salomo regerade i Jerusalem över hela Israel var fyrtio år.
Och Salomo gick till vila hos sina fäder och blev begraven i sin fader Davids stad.
Och hans son Rehabeam blev konung efter honom.
Och Rehabeam drog till Sikem, ty hela Israel hade kommit till Sikem för att göra honom till konung.
När Jerobeam, Nebats son, hörde detta -- han var då ännu kvar i Egypten, dit han hade flytt för konung Salomo; Jerobeam bodde alltså i Egypten,
men de sände ditbort och läto kalla honom åter -- då kom han tillstädes jämte Israels hela församling och talade till Rehabeam och sade:
»Din fader gjorde vårt ok för svårt; men lätta nu du det svåra arbete och det tunga ok som din fader lade på oss, så vilja vi tjäna dig.»
Han svarade dem: »Gån bort och vänten ännu tre dagar, och kommen så tillbaka till mig.»
Och folket gick.
Då rådförde sig konung Rehabeam med de gamle som hade varit i tjänst hos hans fader Salomo, medan denne ännu levde; han sade: »Vilket svar råden I mig att giva detta folk?»
De svarade honom och sade: »Om du i dag underkastar dig detta folk och bliver dem till tjänst, om du lyssnar till deras bön och talar goda ord till dem, så skola de för alltid bliva dina tjänare.»
Men han aktade icke på det råd som de gamle hade givit honom, utan rådförde sig med de unga män som hade vuxit upp med honom, och som nu voro i hans tjänst.
Han sade till dem: »Vilket svar råden I oss att giva detta folk som har talat till mig och sagt: 'Lätta det ok som din fader har lagt på oss'?»
De unga männen som hade vuxit upp med honom svarade honom då och sade: »Så bör du säga till detta folk som har talat till dig och sagt: 'Din fader gjorde vårt ok tungt, men lätta du det för oss' -- så bör du tala till dem: 'Mitt minsta finger är tjockare än min faders länd.
Så veten nu, att om min fader har belastat eder med ett tungt ok, så skall jag göra edert ok ännu tyngre; har min fader tuktat eder med ris, så skall jag tukta eder med skorpiongissel.'»
Så kom nu Jerobeam med allt folket till Rehabeam på tredje dagen, såsom konungen hade befallt, i det han sade: »Kommen tillbaka till mig på tredje dagen.»
Då gav konungen folket ett hårt svar; ty han aktade icke på det råd som de gamle hade givit honom.
Han talade till dem efter de unga männens råd och sade: »Har min fader gjort edert ok tungt, så skall jag göra edert ok ännu tyngre; har min fader tuktat eder med ris, så skall jag tukta eder med skorpiongissel.»
Alltså hörde konungen icke på folket; ty det var så skickat av HERREN, för att hans ord skulle uppfyllas, det som HERREN hade talat till Jerobeam, Nebats son, genom Ahia från Silo.
Då nu hela Israel förnam att konungen icke ville höra på dem, gav folket konungen detta svar: »Vad del hava vi i David?
Ingen arvslott hava vi i Isais son.
Drag hem till dina hyddor, Israel.
Se nu själv om ditt hus, du David.»
Därefter drog Israel hem till sina hyddor.
Allenast över de israeliter som bodde i Juda städer förblev Rehabeam konung.
Och när konung Rehabeam sände åstad Adoram, som hade uppsikten över de allmänna arbetena, stenade hela Israel denne till döds; och konung Rehabeam själv måste med hast stiga upp i sin vagn och fly till Jerusalem.
Så avföll Israel från Davids hus och har varit skilt därifrån ända till denna dag.
Men när hela Israel hörde att Jerobeam hade kommit tillbaka, sände de och läto kalla honom till folkförsamlingen och gjorde honom till konung över hela Israel; ingen höll sig till Davids hus, utom Juda stam allena.
Och när Rehabeam kom till Jerusalem, församlade han hela Juda hus och Benjamins stam, ett hundra åttio tusen utvalda krigare, för att de skulle strida mot Israels hus och återvinna konungadömet åt Rehabeam, Salomos son.
Men Guds ord kom till gudsmannen Semaja;
han sade: »Säg till Rehabeam, Salomos son, Juda konung, och till hela Juda hus och Benjamin och till det övriga folket:
Så säger HERREN: I skolen icke draga upp och strida mot edra bröder, Israels barn.
Vänden tillbaka hem, var och en till sitt, ty vad som har skett har kommit från mig.»
Och de lyssnade till HERRENS ord och vände om och gingo sin väg, såsom HERREN hade befallt.
Men Jerobeam befäste Sikem i Efraims bergsbygd och bosatte sig där.
Därifrån drog han åstad och befäste Penuel.
Och Jerobeam sade vid sig själv: »Såsom nu är, kan riket komma tillbaka till Davids hus.
Ty om folket här får draga upp och anställa slaktoffer i HERRENS hus i Jerusalem, så kan folkets hjärta vända tillbaka till deras herre Rehabeam, Juda konung; ja, då kunna de dräpa mig och vända tillbaka till Rehabeam, Juda konung.»
Sedan nu konungen hade överlagt härom, lät han göra två kalvar av guld.
Därefter sade han till folket: »Nu må det vara nog med edra färder upp till Jerusalem.
Se, här är din Gud, Israel, han som har fört dig upp ur Egyptens land.»
Och han ställde upp den ena i Betel, och den andra satte han upp i Dan.
Detta blev en orsak till synd; folket gick ända till Dan för att träda fram inför den ena av dem.
Han byggde också upp offerhöjdshus och gjorde till präster allahanda män ur folket, sådana som icke voro av Levi barn.
Och Jerobeam anordnade en högtid i åttonde månaden, på femtonde dagen i månaden, lik högtiden Juda, och steg då upp till altaret; så gjorde han i Betel för att offra åt de kalvar som han hade låtit göra.
Och de män som han hade gjort till offerhöjdspräster lät han göra tjänst i Betel.
Till det altare som han hade gjort i Betel steg han alltså upp på femtonde dagen i åttonde månaden, den månad som han av eget påfund hade valt.
Han anordnade nämligen då en högtid för Israels barn och steg upp till altaret för att där tända offereld.
Men då kom på HERRENS befallning en gudsman från Juda till Betel, just när Jerobeam stod vid altaret för att där tända offereld.
Och mannen ropade mot altaret på HERRENS befallning och sade: »Altare!
Altare!
Så säger HERREN: Se, åt Davids hus skall födas en son vid namn Josia, han skall på dig slakta offerhöjdsprästerna som antända offereld på dig, och människoben skall man då bränna upp på dig.»
På samma gång angav han ett tecken, i det han sade: »Detta är tecknet på att det är HERREN som har talat: se, altaret skall rämna, och askan därpå skall spillas ut.»
När konung Jerobeam hörde dessa ord, som gudsmannen ropade mot altaret i Betel, räckte han ut sin hand från altaret och sade: »Gripen honom.»
Men handen som han hade räckt ut mot honom förvissnade, och han kunde icke draga den tillbaka till sig igen.
Och altaret rämnade, och askan på altaret spilldes ut; det var det tecken som gudsmannen på HERRENS befallning hade angivit.
Då tog konungen till orda och sade till gudsmannen: »Bönfall inför HERREN, din Gud, och bed för mig att jag må kunna draga min hand tillbaka till mig igen.»
Och gudsmannen bönföll inför HERREN; och konungen kunde då draga sin hand tillbaka till sig igen, och den var likadan som förut.
Då talade konungen till gudsmannen: »Kom hem med mig och vederkvick dig; sedan vill jag giva dig en gåva.»
Men gudsmannen svarade konungen: »Om du än vill giva mig hälften av vad som finnes i ditt hus, så kommer jag dock icke med dig; här på orten vill jag varken äta eller dricka.
Ty så har HERREN genom sitt ord bjudit mig och sagt: Du skall varken äta eller dricka, och ej heller vända tillbaka samma väg du har gått hit.»
Därefter gick han sina färde en annan väg och vände icke tillbaka samma väg han hade kommit till Betel.
Men i Betel bodde en gammal profet.
Dennes son kom och förtäljde för honom allt vad gudsmannen den dagen hade gjort i Betel, huru han hade talat till konungen.
När de hade förtäljt detta för sin fader,
frågade deras fader dem vilken väg han hade gått.
Och hans söner visste vilken väg gudsmannen som kom från Juda hade gått.
Då sade han till sina söner: »Sadlen åsnan åt mig.»
När de då hade sadlat åsnan åt honom, satte han sig på den
och begav dig åstad efter gudsmannen och fann honom sittande under terebinten; och han frågade honom: »Är du den gudsman som har kommit från Juda?»
Han svarade: »Ja.»
Då sade han till honom: »Kom med mig hem och ät med mig.»
Men han svarade: »Jag kan icke vända om med dig och följa dig, och jag vill icke äta eller dricka med dig här på orten;
ty så har blivit mig sagt genom HERRENS ord: Du skall varken äta eller dricka där; du skall icke heller gå tillbaka samma väg du har gått dit.»
Han sade till honom: »Jag är ock en profet såsom du, och en ängel har talat till mig på HERRENS befallning och sagt: 'För honom tillbaka med dig hem och giv honom att äta och dricka.'»
Men häri ljög han för honom.
Då vände han tillbaka med honom och åt i hans hus och drack.
Men under det att de sutto till bords, kom HERRENS ord till profeten som hade fört honom tillbaka.
Och han ropade till gudsmannen som hade kommit från Juda och sade: »Så säger HERREN: Därför att du har varit gensträvig mot HERRENS ord och icke hållit det bud som HERREN, din Gud, har givit dig,
utan vänt tillbaka och ätit och druckit på den ort där han hade förbjudit, dig att äta och dricka, därför skall din döda kropp icke komma i dina fäders grav.
Sedan han nu hade ätit och druckit, sadlade han åsnan åt honom, åt profeten som han hade fört tillbaka.
Och denne begav sig åstad; men ett lejon kom emot honom på vägen och dödade honom.
Sedan låg hans döda kropp utsträckt där på vägen, under det att åsnan stod bredvid den; och lejonet stod också bredvid den döda kroppen.
Då nu folk som gick därförbi fick se den döda kroppen ligga utsträckt på vägen och lejonet stå bredvid den döda kroppen, gingo de in i staden där den gamle profeten bodde och omtalade det där.
När profeten, som hade fört honom tillbaka från hans väg, hörde det, sade han: »Det är gudsmannen, han som var gensträvig mot HERRENS ord; därför har HERREN givit honom i lejonets våld, och det har krossat och dödat honom, i enlighet med det ord som HERREN hade talat till honom.»
Därefter tillsade han sina söner att de skulle sadla åsnan åt honom; och de sadlade den.
Så begav han sig åstad och fann den döda kroppen liggande utsträckt på vägen och åsnan och lejonet stående bredvid den döda kroppen; lejonet hade icke ätit av den döda kroppen och ej heller krossat åsnan.
Då tog profeten upp gudsmannens döda kropp och lade den på åsnan och förde den tillbaka; och den gamle profeten begav sig in i sin stad för att hålla dödsklagan och begrava honom.
Och han lade hans döda kropp i sin egen grav; och de höllo dödsklagan efter honom och ropade: »Ack ve, min broder!»
Då han nu hade begravit honom, sade han till sina söner: »När jag dör, så begraven mig i den grav där gudsmannen ligger begraven; läggen mina ben vid sidan av hans ben.
Ty förvisso skall det ord gå i fullbordan, som han på HERRENS befallning ropade mot altaret i Betel och mot alla offerhöjdshus i Samariens städer.»
Dock vände Jerobeam efter detta icke om från sin onda väg, utan gjorde åter allahanda man ur folket till offerhöjdspräster; vem som hade lust därtill fick av honom mottaga handfyllning till att vara offerhöjdspräst.
På detta sätt blev han för Jerobeams hus en orsak till synd, och en orsak till att det blev utplånat och utrotat från jorden.
Vid den tiden blev Abia, Jerobeams son, sjuk.
Då sade Jerobeam till sin hustru: »Stå upp och förkläd dig, så att ingen kan märka att du är Jerobeams hustru, och gå till Silo, ty där bor profeten Ahia, han som förkunnade om mig att jag skulle bliva konung över detta folk.
Och tag med dig tio bröd, därtill smått bakverk och en kruka honung, och gå in till honom; han skall då förkunna för dig huru det skall gå med gossen.»
Jerobeams hustru gjorde så; hon stod upp och gick till Silo och kom till Ahias hus.
Och Ahia kunde icke se, ty hans ögon voro starrblinda av ålderdom.
Men HERREN hade sagt till Ahia: »Just nu kommer Jerobeams hustru för att förfråga sig hos dig om sin son, ty han är sjuk; så och så skall du tala till henne.
Men när hon kommer, skall hon ställa sig främmande.
Då nu Ahia hörde ljudet av hennes steg, när hon kom i dörren, sade han: »Kom in, du Jerobeams hustru.
Varför ställer du dig främmande?
Jag har ju fått uppdrag att giva dig ett hårt budskap.
Gå och säg Jerobeam: Så säger HERREN, Israels Gud: Se, jag har upphöjt dig ur folket och satt dig till furste över mitt folk Israel
och har ryckt riket från Davids hus och givit det åt dig.
Men du har icke varit sådan som min tjänare David, som höll mina bud och följde efter mig av allt sitt hjärta, så att han gjorde allenast vad rätt var i mina ögon;
utan du har gjort mer ont än alla som hava varit före dig och har gått bort och gjort dig andra gudar, nämligen gjutna beläten, för att förtörna mig, och har kastat mig bakom din rygg.
Därför skall jag låta olycka komma över Jerobeams hus och utrota allt mankön av Jerobeams hus, både små och stora i Israel; och jag skall bortsopa Jerobeams hus, såsom man sopar bort orenlighet, till dess det bliver en ände därpå.
Den av Jerobeams hus, som dör i staden, skola hundarna äta upp, och den som dör ute på marken, skola himmelens fåglar äta upp.
Ty så har HERREN talat.
Så stå du nu upp och gå hem igen.
När din fot träder in i staden, skall barnet dö.
Och hela Israel skall hålla dödsklagan efter honom, och man skall begrava honom; ty av Jerobeams hus skall allenast han komma i en grav, därför att i Jerobeams hus dock hos honom blev funnet något som var gott inför HERREN, Israels Gud.
Men HERREN skall låta en konung över Israel uppstå åt sig, en konung som skall utrota Jerobeams hus.
Detta är den dagen; och vad skall icke nu ske!
HERREN skall slå Israel, så att det bliver likt vassen, som vaggar hit och dit i vattnet.
Och han skall rycka upp Israel ur detta goda land, som han har givit åt deras fäder, och skall förströ dem på andra sidan floden, därför att de hava gjort sig Aseror och därmed förtörnat HERREN.
Och han skall prisgiva Israel för de synders skull som Jerobeam har begått, och genom vilka han har kommit Israel att synda.»
Då stod Jerobeams hustru upp och gick sin väg och kom till Tirsa; och just som hon beträdde husets tröskel, gav gossen upp andan.
Och man begrov honom, och hela Israel höll dödsklagan efter honom, i enlighet med det ord som HERREN hade talat genom sin tjänare, profeten Ahia.
Vad nu mer är att säga om Jerobeam, om hans krig och om hans regering, det finnes upptecknat i Israels konungars krönika.
Den tid Jerobeam regerade var tjugutvå år.
Så gick han till vila hos sina fäder; och hans son Nadab blev konung efter honom.
Men Rehabeam, Salomos son, var konung i Juda.
Fyrtioett år gammal var Rehabeam, när han blev konung, och han regerade sjutton år i Jerusalem, den stad som HERREN hade utvalt ur alla Israels stammar, till att där fästa sitt namn.
Hans moder hette Naama, ammonitiskan.
Och Juda gjorde vad ont var i HERRENS ögon; med de synder som de begingo retade de honom långt mer, än deras fäder hade gjort.
Ty också de byggde sig offerhöjder och reste stoder och Aseror på alla höga kullar och under alla gröna träd;
ja, också tempelbolare funnos i landet.
De gjorde efter alla styggelser hos de folk som HERREN hade fördrivit för Israels barn.
Men i konung Rehabeams femte regeringsår drog Sosak, konungen i Egypten, upp mot Jerusalem.
Och han tog skatterna i HERRENS hus och skatterna i konungshuset; alltsammans tog han.
Han tog ock alla de gyllene sköldar som Salomo hade låtit göra.
I deras ställe lät konung Rehabeam göra sköldar av koppar, och dessa lämnade han i förvar åt hövitsmännen för drabanterna som höllo vakt vid ingången till konungshuset.
Och så ofta konungen gick till HERRENS hus, buro drabanterna dem; sedan förde de dem tillbaka till drabantsalen.
Vad nu mer är att säga om Rehabeam och om allt vad han gjorde, det finnes upptecknat i Juda konungars krönika.
Men Rehabeam och Jerobeam lågo i krig med varandra, så länge de levde.
Och Rehabeam gick till vila hos sina fäder och blev begraven hos sina fäder i Davids stad.
Hans moder hette Naama, ammonitiskan.
Och hans son Abiam blev konung efter honom.
I konung Jerobeams, Nebats sons, adertonde regeringsår blev Abiam konung över Juda.
Han regerade tre år i Jerusalem.
Hans moder hette Maaka, Abisaloms dotter.
Och han vandrade i alla de synder som hans fader hade begått före honom, och hans hjärta var icke hängivet åt HERREN, hans Gud, såsom hans fader Davids hjärta hade varit.
Allenast för Davids skull lät HERREN, hans Gud, honom få en lampa i Jerusalem, i det att han uppsatte hans son efter honom och lät Jerusalem hava bestånd --
detta därför att David gjorde vad rätt var i HERRENS ögon och icke vek ifrån något som han bjöd honom, så länge han levde, utom i saken med hetiten Uria.
Men Rehabeam och Jerobeam lågo i krig med varandra, så länge den förre levde.
Vad nu mer är att säga om Abiam och om allt vad han gjorde, det finnes upptecknat i Juda konungars krönika.
Men Abiam och Jerobeam lågo i krig med varandra.
Och Abiam gick till vila hos sina fäder, och man begrov honom i Davids stad.
Och hans son Asa blev konung efter honom.
I Jerobeams, Israels konungs, tjugonde regeringsår blev Asa konung över Juda.
Han regerade fyrtioett år i Jerusalem.
Hans moder hette Maaka, Abisaloms dotter.
Och Asa gjorde vad rätt var i HERRENS ögon, såsom hans fader David hade gjort
Han drev ut tempelbolarna ur landet och skaffade bort alla de eländiga avgudabeläten som hans fader hade låtit göra.
Ja, sin moder Maaka avsatte han från hennes drottningsvärdighet, därför att hon hade satt upp en styggelse åt Aseran; Asa högg nu ned styggelsen och brände upp den i Kidrons dal.
Men offerhöjderna blevo icke avskaffade; dock var Asas hjärta hängivet åt HERREN, så länge han levde.
Och han förde in i HERRENS hus både vad hans fader och vad han själv hade helgat åt HERREN: silver, guld och kärl.
Men Asa och Baesa, Israels konung, lågo i krig med varandra, så länge de levde.
Baesa, Israels konung, drog upp mot Juda och begynte befästa Rama, för att hindra att någon komme vare sig till eller ifrån Asa, Juda konung.
Då tog Asa allt silver och guld som fanns kvar i skattkamrarna i HERRENS hus, ävensom skatterna i konungshuset, och lämnade detta åt sina tjänare; därefter sände konung Asa dem till Ben-Hadad, son till Tabrimmon, son till Hesjon, konungen i Aram, som bodde i Damaskus, och lät säga:
»Ett förbund består ju mellan mig och dig, såsom det var mellan min fader och din fader.
Se, här sänder jag dig skänker av silver och guld, så bryt då nu ditt förbund med Baesa, Israels konung, för att han må lämna mig i fred.»
Och Ben-Hadad lyssnade till konung Asa och sände sina krigshövitsmän mot Israels städer och förhärjade Ijon, Dan, Abel-Bet-Maaka och hela Kinarot jämte hela Naftali land.
När Baesa hörde detta, avstod han från att befästa Rama och höll sig sedan stilla i Tirsa.
Men konung Asa bådade upp hela Juda, ingen fritagen; och de förde bort stenar och trävirke som Baesa använde till att befästa Rama.
Därmed befäste nu konung Asa Geba i Benjamin, så ock Mispa.
Allt vad mer är att säga om Asa, om alla hans bedrifter, om allt vad han gjorde och om de städer han byggde, det finnes upptecknat i Juda konungars krönika.
Men på sin ålderdom fick han en sjukdom i sina fötter.
Och Asa gick till vila hos sina fäder och blev begraven hos sina fäder i sin fader Davids stad.
Och hans son Josafat blev konung efter honom.
Men Nadab, Jerobeams son, blev konung över Israel i Asas, Juda konungs, andra regeringsår, och han regerade över Israel i två år.
Han gjorde vad ont var i HERRENS ögon och vandrade på sin faders väg och i den synd genom vilken denne hade kommit Israel att synda.
Men Baesa, Ahias son, av Isaskar hus, anstiftade en sammansvärjning mot honom, och Baesa dräpte honom vid Gibbeton, som tillhörde filistéerna; Nadab med hela Israel höll nämligen på med att belägra Gibbeton.
I Asas, Juda konungs, tredje regeringsår var det som Baesa dödade honom, och han blev så själv konung i hans ställe.
Och när han hade blivit konung förgjorde han hela Jerobeams hus; han lät intet som anda hade bliva kvar av Jerobeams hus, utan utrotade det, i enighet med det ord som HERREN hade talat genom sin tjänare Ahia från Silo --
detta för de synders skull som Jerobeam hade begått, och genom vilka han kom Israel att synda, så att han därmed förtörnade HERREN, Israels Gud.
Vad nu mer är att säga om Nadab och om allt vad han gjorde det finnes upptecknat i Israels konungars krönika.
Men Asa och Baesa, Israels konung, lågo i krig med varandra, länge de levde.
I Asas, Juda konungs, tredje regeringsår blev Baesa, Ahias son, konung över hela Israel i Tirsa och regerade i tjugufyra år.
Han gjorde vad ont var i HERRENS ögon och vandrade på Jerobeams väg och i den synd genom vilken denne hade kommit Israel att synda.
Och HERRENS ord kom till Jehu, Hananis son, mot Baesa; han sade:
»Se, jag har lyft dig upp ur stoftet och satt dig till furste över mitt folk Israel.
Men du har vandrat på Jerobeams väg och kommit mitt folk Israel att synda, så att de hava förtörnat mig genom sina synder.
Därför vill jag bortsopa Baesa och hans hus; ja, jag vill göra med ditt hus såsom jag gjorde med Jerobeams, Nebats sons, hus.
Den av Baesas hus, som dör i staden, skola hundarna äta upp, och den av hans hus, som dör ute på marken, skola himmelens fåglar äta upp.»
Vad nu mer är att säga om Baesa, om vad han gjorde och om hans bedrifter, det finnes upptecknat i Israels konungars krönika.
Och Baesa gick till vila hos sina fäder och blev begraven i Tirsa.
Och hans son Ela blev konung efter honom.
Men genom profeten Jehu, Hananis son, hade HERRENS ord kommit till Baesa och hans hus, icke allenast för allt det onda som han hade gjort i HERRENS ögon, då han förtörnade honom genom sina händers verk, så att det måste gå honom såsom det gick Jerobeams hus, utan ock därför att han hade förgjort detta.
I Asas, Juda konungs, tjugusjätte regeringsår blev Ela, Baesas son, konung över Israel i Tirsa och regerade i två år.
Men hans tjänare Simri, som var hövitsman för den ena hälften av stridsvagnarna, anstiftade en sammansvärjning mot honom.
Och en gång, då han i Tirsa hade druckit sig drucken i Arsas hus, överhovmästarens i Tirsa,
kom Simri dit och slog honom till döds -- det var i Asas, Juda konungs, tjugusjunde regeringsår -- och han själv blev så konung i hans ställe.
Och när han hade blivit konung och intagit sin tron, förgjorde han hela Baesas hus, utan att låta någon av mankön bliva kvar, varken hans blodsförvanter eller hans vänner.
Så utrotade Simri hela Baesas hus, i enlighet med det ord som HERREN hade talat till Baesa genom profeten Jehu --
detta för alla de synders skull som Baesa och hans son Ela hade begått, och genom vilka de hade kommit Israel att synda, så att de förtörnade HERREN, Israels Gud, med de fåfängliga avgudar som de dyrkade.
Vad nu mer är att säga om Ela och om allt vad han gjorde, det finnes upptecknat i Israels konungars krönika.
I Asas, Juda konungs, tjugusjunde regeringsår blev Simri konung och regerade i sju dagar, i Tirsa.
Folket höll då på att belägra Gibbeton, som tillhörde filistéerna.
Medan nu folket höll på med belägringen, fingo de höra sägas »Simri har anstiftat en sammansvärjning; han har ock dräpt konungen.»
Då gjorde hela Israel samma dag Omri, den israelitiske härhövitsmannen, till konung, i lägret.
Därefter drog Omri med hela Israel upp från Gibbeton, och de angrepo Tirsa.
Men när Simri såg att staden var intagen, gick han in i konungshusets palatsbyggnad och brände upp konungshuset jämte sig själv i eld och omkom så --
detta för de synders skull som han hade begått, i det att han gjorde vad ont var i HERRENS ögon och vandrade på Jerobeams väg och i den synd som denne hade gjort, och genom vilken han hade kommit Israel att synda.
Vad nu mer är att säga om Simri och om den sammansvärjning som han anstiftade, det finnes upptecknat i Israels konungars krönika.
Nu delade sig Israels folk i två hälfter; den ena hälften av folket höll sig till Tibni, Ginats son, och ville göra honom till konung, och den andra hälften höll sig till Omri.
Men den del av folket som höll sig till Omri, fick överhanden över den del som höll sig till Tibni, Ginats son.
Och när Tibni var död, blev Omri konung.
I Asas, Juda konungs, trettioförsta regeringsår blev Omri konung över Israel och regerade i tolv år; i Tirsa regerade han i sex år.
Han köpte berget Samaria av Semer för två talenter silver; och han bebyggde berget och kallade staden som han byggde där Samaria, efter Semer, den man som hade varit bergets ägare.
Men Omri gjorde vad ont var i HERRENS ögon; han gjorde mer ont än någon av dem som hade varit före honom.
Han vandrade i allt på Jerobeams, Nebats sons, väg och i de synder genom vilka denne hade kommit Israel att synda, så att de förtörnade HERREN, Israels Gud, med de fåfängliga avgudar de dyrkade.
Vad nu mer är att säga om Omri, om vad han gjorde och om de bedrifter han utförde, det finnes upptecknat i Israels konungars krönika.
Och Omri gick till vila hos sina fäder och blev begraven i Samaria.
Och hans son Ahab blev konung efter honom.
Ahab, Omris son, blev konung över Israel i Asas, Juda konungs, trettioåttonde regeringsår; sedan regerade Ahab, Omris son, i tjugutvå år över Israel i Samaria.
Men Ahab, Omris son, gjorde vad ont var i HERRENS ögon, mer än någon av dem som hade varit före honom.
Det var honom icke nog att vandra i Jerobeams, Nebats sons, synder; han tog ock till hustru Isebel, dotter till Etbaal, sidoniernas konung, och gick så åstad och tjänade Baal och tillbad honom.
Och han reste ett altare åt Baal i Baalstemplet som han hade byggt i Samaria.
Därtill lät Ahab göra Aseran.
Så gjorde Ahab mer till att förtörna HERREN, Israels Gud, än någon av de Israels konungar som hade varit före honom.
Under hans tid byggde beteliten Hiel åter upp Jeriko.
Men när han lade dess grund, kostade det honom hans äldste son Abiram, och när han satte upp dess portar, kostade det honom hans yngste son Segib -- i enlighet med det ord som HERREN hade talat genom Josua, Nuns son.
Och tisbiten Elia, en man som förut hade uppehållit sig i Gilead, sade till Ahab: »Så sant HERREN, Israels Gud, lever, han vilkens tjänare jag är, under dessa år skall varken dagg eller regn falla, med mindre jag säger det.»
Och HERRENS ord kom till honom; han sade:
»Gå bort härifrån och begiv dig österut, och göm dig vid bäcken Kerit, som österifrån rinner ut i Jordan.
Din dryck skall du få ur bäcken, och korparna har jag bjudit att där förse dig med föda.»
Då gick han bort och gjorde såsom HERREN hade befallt; han gick bort och uppehöll sig vid bäcken Kerit, som österifrån rinner ut i Jordan.
Och korparna förde till honom bröd och kött om morgonen, och bröd och kött om aftonen, och sin dryck fick han ur bäcken.
Men efter någon tid torkade bäcken ut, därför att det icke regnade i landet.
Då kom HERRENS ord till honom; han sade:
»Stå upp och gå till Sarefat, som hör till Sidon, och uppehåll dig där.
Se, jag har där bjudit en änka att förse dig med föda.»
Han stod upp och gick till Sarefat.
Och när han kom till stadsporten, fick han där se en änka som samlade ved.
Då ropade han till henne och sade: »Hämta litet vatten åt mig i kärlet, så att jag får dricka.»
När hon nu gick för att hämta det, ropade han efter henne och sade: »Tag ock med dig ett stycke bröd åt mig.»
Men hon svarade: »Så sant HERREN, din Gud, lever, jag äger icke en kaka bröd, utan allenast en hand full mjöl i krukan och litet olja i kruset.
Och se, här har jag samlat ihop ett par vedpinnar, och jag går nu hem och tillreder det åt mig och min son, för att vi må äta det och sedan dö.»
Då sade Elia till henne: »Frukta icke; gå och gör såsom du har sagt.
Men red först till en liten kaka därav åt mig, och bär ut den till mig; red sedan till åt dig och din son.
Ty så säger HERREN, Israels Gud: Mjölet i krukan skall icke taga slut, och oljan i kruset skall icke tryta, intill den dag då HERREN låter det regna på jorden.»
Då gick hon åstad och gjorde såsom Elia hade sagt.
Och hon hade sedan att äta, hon själv och han och hennes husfolk, en lång tid.
Mjölet i krukan tog icke slut, och oljan i kruset tröt icke, i enlighet med det ord som HERREN hade talat genom Elia.
Men härefter hände sig, att kvinnans, hans värdinnas, son blev sjuk; hans sjukdom blev mycket svår, så att han till slut icke mer andades.
Då sade hon till Elia: »Vad har du med mig att göra, du gudsman?
Du har kommit till mig, för att min missgärning skulle bliva ihågkommen, så att min son måste dö.»
Men han sade till henne: »Giv mig din son.»
Och han tog honom ur hennes famn och bar honom upp i salen där han bodde och lade honom på sin säng.
Och han ropade till HERREN och sade: »HERRE, min Gud, har du väl kunnat göra så illa mot denna änka, vilkens gäst jag är, att du har dödat hennes son?»
Därefter sträckte han sig ut över gossen tre gånger och ropade till HERREN och sade: »HERRE, min Gud, låt denna gosses själ komma tillbaka in i honom.»
Och HERREN hörde Elias röst, och gossens själ kom tillbaka in i honom, och han fick liv igen.
Och Elia tog gossen och bar honom från salen ned i huset och gav honom åt hans moder.
Och Elia sade: »Se, din son lever.»
Då sade kvinnan till Elia: »Nu vet jag att du är en gudsman, och att HERRENS ord i din mun är sanning.»
En lång tid härefter, på tredje året, kom HERRENS ord till Elia; han sade: »Gå åstad och träd fram för Ahab, så skall jag sedan låta det regna på jorden.»
Då gick Elia åstad för att träda fram för Ahab.
Men hungersnöden var då stor i Samaria.
Och Ahab kallade till sig Obadja, sin överhovmästare; men Obadja dyrkade HERREN med stor iver.
Och när Isebel utrotade HERRENS profeter, hade Obadja tagit ett hundra profeter och gömt dem, femtio man åt gången, i en grotta och försett dem med mat och dryck.
Ahab sade nu till Obadja: »Far igenom landet till alla vattenkällor och alla bäckar.
Kanhända skola vi finna gräs, så att vi kunna behålla hästar och mulåsnor vid liv och slippa att slakta ned någon boskap.»
Och de fördelade mellan sig landet som de skulle draga i genom.
Ahab for en väg för sig, och Obadja for en annan väg för sig.
När nu Obadja färdades sin väg fram, fick han se Elia komma emot sig.
Och han kände igen denne och föll ned på Sitt ansikte och sade: »Är du här, min herre Elia?»
Han svarade honom: »Ja.
Gå och säg till din herre: 'Elia är här.'»
Då sade han: »Varmed har jag försyndat mig, eftersom du vill giva din tjänare i Ahabs hand och låta honom döda mig?
Så sant HERREN, din Gud, lever, det finnes icke något folk eller något rike dit min herre icke har sänt för att söka efter dig; och om man har svarat: 'Han är icke här', så har han av det riket eller det folket tagit en ed, att man icke har funnit dig.
Och nu säger du: 'Gå och säg till din herre: Elia är här!'
Om nu, när jag går ifrån dig, HERRENS Ande skulle rycka bort dig, jag vet icke vart, och jag likväl komme med ditt budskap till Ahab, så skulle han dräpa mig, när han icke funne dig.
Och dock har ju jag, din tjänare, fruktat HERREN allt ifrån min ungdom.
Har det icke blivit berättat för min herre vad jag gjorde, när Isebel dräpte HERRENS profeter, huru jag gömde ett hundra av HERRENS profeter, femtio man och åter femtio, i en grotta och försåg dem med mat och dryck?
Och nu säger du: 'Gå och säg till din herre: Elia är här!' -- för att han skall dräpa mig.»
Men Elia svarade: »Så sant HERREN Sebaot lever, han vilkens tjänare jag är, redan i dag skall jag träda fram för honom.»
Då gick Obadja Ahab till mötes och förkunnade detta för honom; och Ahab begav sig åstad för att möta Elia.
Och när Ahab fick se Elia, sade Ahab till honom: »Är du här, du som drager olycka över Israel?»
Han svarade: »Det är icke jag, som drager olycka över Israel, utan du och din faders hus, därmed att I övergiven HERRENS bud, och därmed att du följer efter Baalerna.
Men sänd nu bort och församla hela Israel till mig på berget Karmel, jämte Baals fyra hundra femtio profeter och Aserans fyra hundra profeter, som äta vid Isebels bord.»
Då sände Ahab omkring bland Israels barn och lät församla profeterna på berget Karmel.
Och Elia trädde fram för allt folket och sade: »Huru länge viljen I halta på båda sidor?
Är det HERREN som är Gud, så följen efter honom; men om Baal är det, så följen efter honom.»
Och folket svarade honom icke ett ord.
Då sade Elia till folket: »Jag allena är kvar såsom HERRENS Profet, och Baals profeter äro fyra hundra femtio man.
Må man nu giva oss två tjurar, och må de välja ut åt sig den ena tjuren och stycka den och lägga den på veden, utan att tända eld därpå, så vill jag reda till den andra tjuren och lägga den på veden, utan att tända eld därpå.
Därefter mån I åkalla eder guds namn, men själv vill jag åkalla HERRENS namn. »Den gud som då svarar med eld, han vare Gud.»
Allt folket svarade och sade. »Ditt förslag är gott.»
Då sade Elia till Baals profeter: »Väljen ut åt eder den ena tjuren och reden till den, I först, ty I ären flertalet; åkallen därefter eder guds namn, men eld fån I icke tända.»
Då togo de den tjur som han gav dem och redde till den; sedan åkallade de Baals namn från morgonen ända till middagen och ropade: »Baal, svara oss.»
Men icke ett ljud hördes, och ingen svarade.
Och alltjämt haltade de åstad kring altaret som man hade gjort.
När det så blev middag, gäckades Elia med dem och sade: »Ropen ännu högre, ty visserligen är han en gud, men han har väl något att begrunda, eller ock har han gått avsides, eller är han på resa; kanhända sover han, men då skall han väl vakna.»
Då ropade de ännu högre och ristade sig, såsom deras sed var, med svärd och spjut, så att blodet kom ut på dem.
När det sedan hade blivit eftermiddag, fattades de av profetiskt raseri, och höllo så på ända till den tid då spisoffret frambäres.
Men icke ett ljud hördes, ingen svarade, och ingen tycktes heller akta på dem.
Och Elia sade till allt folket: »Träden hitfram till mig.»
Så trädde nu allt folket fram till honom.
Då satte han åter i stånd HERRENS altare, som hade blivit nedrivet.
Elia tog tolv stenar, lika många som Jakobs söners stammar -- den mans, till vilken detta HERRENS ord hade kommit: »Israel skall vara ditt namn.»
Och han byggde av stenarna ett altare i HERRENS namn och gjorde omkring altaret en grav, stor nog för ett utsäde av två sea-mått.
Därefter lade han upp veden, styckade tjuren och lade den på veden.
Sedan sade han: »Fyllen fyra krukor med vatten, och gjuten ut vattnet över brännoffret och veden.»
Han sade ytterligare: »Gören så ännu en gång.»
Och de gjorde så för andra gången.
Därefter sade han: »Gören så för tredje gången.»
Och de gjorde så för tredje gången.
Och vattnet flöt runt omkring altaret; och han lät fylla också graven med vatten.
Då nu tiden var inne att frambära spisoffret, trädde profeten Elia fram och sade: »HERRE, Abrahams, Isaks och Israels Gud, låt det i dag bliva kunnigt att du är Gud i Israel, och att jag är din tjänare, och att det är på din befallning jag har gjort allt detta.»
Svara mig, HERRE, svara mig, så att detta folk förnimmer att det är du, HERRE, som är Gud, i det att du vänder om deras hjärtan.»
»Då föll HERRENS ed ned och förtärde brännoffret, veden, stenarna och jorden, och uppslickade vattnet som var i graven.
När allt folket såg detta, föllo de ned på sina ansikten och sade: »HERREN är det som är Gud!
HERREN är det som är Gud!»
Men Elia sade till dem: »Gripen Baals profeter; låten ingen av dem komma undan.»
Och de grepo dem.
Och Elia lät föra dem ned till bäcken Kison och slakta dem där.
Och Elia sade till Ahab: »Begiv dig ditupp, ät och drick, ty jag hör bruset av regn.»
Då begav sig Ahab ditupp för att äta och dricka.
Men Elia steg upp på Karmels topp, hukade sig ned mot jorden och sänkte sitt ansikte mellan sina knän.
Och han sade till sin tjänare »Gå upp och skåda ut åt havet.»
Denne gick då upp och skådade ut, men sade: »Jag ser ingenting.»
Så tillsade han honom sju gånger att gå tillbaka.
När han då kom dit sjunde gången sade han: »Nu ser jag ett litet moln, icke större än en mans hand, stiga upp ur havet.»
Då sade han: »Gå upp och säg till Ahab: Spänn för och far ned, så att regnet icke håller dig kvar.»
Och i ett ögonblick förmörkades himmelen av moln och storm, och ett starkt regn föll.
Och Ahab steg upp i sin vagn och for till Jisreel.
Men HERRENS hand hade kommit över Elia, så att han omgjorde sina länder och sprang framför Ahab ända inemot Jisreel.
Men när Ahab berättade för Isebel allt vad Elia hade gjort, och huru han hade dräpt alla profeterna med svärd,
Sände Isebel en budbärare till Elia och lät säga: »Gudarna straffe mig nu och framgent om jag icke i morgon vid denna tid låter det gå med ditt liv såsom det gick med alla dessas liv.»
När han förnam detta, stod han upp och begav sig i väg för att rädda sitt liv, och han kom så till Beer-Seba, som hör till Juda; där lämnade han kvar sin tjänare.
Men själv gick han ut i öknen en dagsresa.
Där satte han sig under en ginstbuske; och han önskade sig döden och sade: »Det är nog; tag nu mitt liv, HERRE, ty jag är icke förmer än mina fäder.»
Därefter lade han sig att sova under en ginstbuske.
Men se, då rörde en ängel vid honom och sade till honom: »Stå upp och ät.»
När han då såg upp, fick han vid sin huvudgärd se ett bröd, sådant som bakas på glödande stenar, och ett krus med vatten.
Och han åt och drack och lade sig åter ned.
Men HERRENS ängel rörde åter vid honom, för andra gången, och sade: »Stå upp och ät, ty eljest bliver vägen dig för lång.»
Då stod han upp och åt och drack, och gick så, styrkt av den maten, i fyrtio dagar och fyrtio nätter, ända till Guds berg Horeb.
Där gick han in i en grotta, och i den stannade han över natten.
Då kom HERRENS ord till honom; han sade till honom: »Vad vill du här, Elia?»
Han svarade: »Jag har nitälskat för HERREN, härskarornas Gud.
Ty Israels barn hava övergivit ditt förbund, rivit ned dina altaren och dräpt dina profeter med svärd; jag allena är kvar, och de stå efter att taga mitt liv.»
Han sade: »Gå ut och ställ dig på berget inför HERREN.»
Då gick HERREN fram där, och en stor och stark storm, som ryckte loss berg och bröt sönder klippor, gick före HERREN; men icke var HERREN i stormen.
Efter stormen kom en jordbävning; men icke var HERREN i jordbävningen.
Efter jordbävningen kom en eld; men icke var HERREN i elden.
Efter elden kom ljudet av en sakta susning.
Så snart Elia hörde detta, skylde han sitt ansikte med manteln och gick ut och ställde sig vid ingången till grottan.
Då kom en röst till honom och sade: »Vad vill du här, Elia?»
Han svarade: »Jag har nitälskat för HERREN, härskarornas Gud.
Ty Israels barn hava övergivit ditt förbund, rivit ned dina altaren och dräpt dina profeter med svärd; jag allena är kvar, och de stå efter att taga mitt liv.»
HERREN sade till honom: »Gå nu tillbaka igen, och tag vägen till Damaskus' öken, och gå in och smörj Hasael till konung över Aram.
Och Jehu, Nimsis son, skall du smörja till konung över Israel.
Och till profet i ditt ställe skall du smörja Elisa, Safats son, från Abel-Mehola.
Och så skall ske: den som kommer undan Hasaels svärd, honom skall Jehu döda, och den som kommer undan Jehus svärd, honom skall Elisa döda.
Men jag skall låta sju tusen män bliva kvar i Israel, alla de knän som icke hava böjt sig för Baal, och var mun som icke har givit honom hyllningskyss.»
När han sedan gick därifrån, träffade han på Elisa, Safats son, som höll på att plöja; tolv par oxar gingo framför honom, och själv körde han det tolfte paret.
Och Elia gick fram till honom och kastade sin mantel över honom.
Då släppte han oxarna och skyndade efter Elia och sade: »Låt mig först få kyssa min fader och min moder, så vill jag sedan följa dig.»
Han sade till honom: »Välan, du må gå tillbaka igen; du vet ju vad jag har gjort med dig.»
Då lämnade han honom och gick tillbaka och tog sina båda oxar och slaktade dem, och med oxarnas ok kokade han deras kött; detta gav han åt folket, och de åto.
Därefter stod han upp och följde Elia och blev hans tjänare.
Och Ben-Hadad, konungen i Aram, samlade hela sin här; han hade med sig trettiotvå konungar jämte hästar och vagnar.
Han drog upp och belägrade Samaria och ansatte det.
Och han skickade sändebud in i staden till Ahab, Israels konung,
och lät säga honom: »Så säger Ben-Hadad: Ditt silver och ditt guld tillhör mig, och det bästa du har av kvinnor och barn tillhör mig ock.»
Israels konung svarade och sade: »Såsom du har sagt, min herre konung: jag själv och allt vad jag har tillhör dig.»
Men sändebuden kommo tillbaka och sade: »Så säger Ben-Hadad: Jag har ju sänt till dig och låtit säga: 'Ditt silver och ditt guld, dina kvinnor och dina barn skall du giva mig.'
Och nu skall jag sannerligen i morgon vid denna tid sända mina tjänare till dig, för att de må genomsöka ditt hus och dina tjänares hus; och allt som är dina ögons lust skola de taga med sig och föra bort.»
Då kallade Israels konung till sig alla de äldste i landet och sade: »Märken och sen huru denne står efter vårt fördärv.
Ty när han sände till mig och begärde mina kvinnor och mina barn, mitt silver och mitt guld, vägrade jag ju icke att giva honom det.»
Alla de äldste och allt folket sade till honom: »Hör icke på honom och gör honom icke till viljes.»
Så svarade han då Ben-Hadads sändebud: »Sägen till min herre konungen: Allt, varom du förra gången sände bud till din tjänare, det vill jag foga mig i; men detta kan jag icke foga mig i.»
Och sändebuden vände tillbaka med detta svar.
Då sände Ben-Hadad till honom och lät säga: »Gudarna straffe mig nu och framgent, om Samarias grus skall räcka till att fylla händerna på allt det folk som följer mig.»
Men Israels konung svarade och sade: »Sägen så: Icke må den som omgjordar sig med svärdet berömma sig likt den som spänner det av sig.»
Så snart Ben-Hadad hörde detta svar, där han satt och drack med konungarna i lägerhyddorna, sade han till sina tjänare: »Gören eder redo.»
Och de gjorde sig redo till att angripa staden.
Då trädde en profet fram till Ahab, Israels konung, och sade: »Så säger HERREN: Ser du hela denna stor hop?
Se, jag vill i dag giva den i din hand, på det att du må förnimma att jag är HERREN.»
Då frågade Ahab: »Genom vem?
Han svarade: »Så säger HERREN: Genom landshövdingarnas män.»
Han frågade ytterligare: »Vem skall begynna striden?»
Han svarade: »Du själv.»
Så mönstrade han då landshövdingarnas män, och de voro två hundra trettiotvå, därefter mönstrade han allt folket, alla Israels barn, sju tusen man.
Och vid middagstiden gjorde de ett utfall, just när Ben-Hadad höll på att dricka sig drucken i lägerhyddorna, tillsammans med de trettiotvå konungar som sade kommit honom till hjälp.
Landshövdingarnas män drogo först ut.
Och de kunskapare som Ben-Hadad sände ut underrättade honom om att folk kom ut från Samaria.
Då sade han: »Om de hava dragit ut i fredlig avsikt, så gripen dem levande; och om de hava dragit ut till strid, så gripen dem ock levande.»
Men när dessa -- landshövdingarnas män och hären som följde dem -- hade kommit ut ur staden,
höggo de ned var och en sin man, och araméerna flydde, och Israel förföljde dem.
Och Ben-Hadad, konungen i Aram, kom undan på en häst, jämte några ryttare.
Och Israels konung drog ut och slog både ryttarhären och vagnshären och tillfogade araméerna ett stort nederlag.
Men profeten trädde fram till Israels konung och sade till honom: »Grip dig nu an; och betänk och se till, vad du bör göra, ty nästa år kommer konungen i Aram att åter draga upp mot dig.»
Men den arameiske konungens tjänare sade till honom: »Deras gud är en bergsgud; därför hava de blivit oss övermäktiga.
Låt oss nu strida mot dem på slätten, så skola vi förvisso bliva dem övermäktiga.
Och vidare måste du göra så: avsätt var och en av konungarna från hans plats, och insätt ståthållare i deras ställe.
Skaffa dig sedan själv en här, lika stor som den du har förlorat, med lika många hästar och lika många vagnar, och låt oss sedan strida mot dem på slätten, så skola vi förvisso bliva dem övermäktiga.»
Och han lyssnade till deras ord och gjorde så.
Följande år mönstrade Ben-Hadad araméerna och drog så upp till Afek för att strida mot Israel.
Israels barn hade ock blivit mönstrade och försedda med livsmedel och tågade därefter emot dem.
Och Israels barn lägrade sig gent emot dem, lika två små gethjordar, under det att araméerna uppfyllde landet.
Då trädde gudsmannen fram och sade till Israels konung: »Så säger HERREN: Därför att araméerna hava sagt: 'HERREN är en bergsgud och icke en dalgud', därför giver jag hela denna stora hop i din hand, på det att I mån förnimma att jag är HERREN.»
Och de voro lägrade mitt emot varandra i sju dagar.
På sjunde dagen kom det till strid, och Israels barn slogo då av araméerna hundra tusen man fotfolk, detta på en enda dag.
De återstående flydde in i staden Afek; men stadsmuren föll ned över tjugusju tusen man, dem som återstodo.
Ben-Hadad flydde också och kom in i staden och sprang från kammare till kammare.
Då sade hans tjänare till honom: »Vi hava hört att konungarna av Israels hus äro nådiga konungar.
Låt oss därför sätta säcktyg om våra länder och rep om våra huvuden och giva oss åt Israels konung; kanhända låter han dig då få leva.»
Och de bundo säcktyg omkring sina länder och rep omkring sina huvuden och kommo så till Israels konung och sade: »Din tjänare Ben-Hadad beder: 'Låt mig få leva.'»
Han svarade: »Är han ännu vid liv, han min broder?»
Männen, som i detta hans ord sågo ett gott varsel, skyndade att taga fasta därpå och sade: »Ja, din broder är Ben-Hadad.»
Han sade: »Gån och hämten honom hit.»
Då gav sig Ben-Hadad åt honom, och han lät honom stiga upp i sin vagn.
Och Ben-Hadad sade till honom: »De städer som min fader tog från din fader vill jag giva tillbaka, och du skall för din räkning få inrätta handelskvarter i Damaskus, såsom min fader fick göra i Samaria.» »Välan», sade Ahab, »på sådana villkor vill jag giva dig fri.»
Och han slöt ett fördrag med honom och gav honom fri.
Och en av profetlärjungarna sade på HERRENS befallning till en annan: »Slå till mig.»
Men mannen vägrade att slå honom.
Då sade han till honom: »Eftersom du icke har lyssnat till HERRENS röst, därför skall ett lejon slå ned dig, när du går ifrån mig.»
Och när han gick sin väg ifrån honom, kom ett lejon emot honom och slog ned honom.
Sedan träffade han en annan man och sade: »Slå till mig.»
Och mannen slog honom så hårt, att sår uppstod därav.
Därefter gick profeten och ställde sig i konungens väg, sedan han hade gjort sig oigenkännlig genom att sätta en bindel över ögonen.
När nu konungen kom därfram, ropade han till konungen och sade: »Din tjänare hade givit sig ut i striden, då i detsamma en man kom därifrån och förde till mig en annan man och sade: 'Vakta denne man; om han kommer bort, skall det gå dig såsom det skulle hava gått honom, eller ock måste du betala en talent silver.'
Nu hände sig, under det din tjänare hade att syssla än här än där, att mannen kom undan.»
Israels konung sade till honom: »Din dom är given; du har ju själv avkunnat den.»
Då tog han skyndsamt bort bindeln från sina ögon, och Israels konung kände igen honom och såg att han var en av profeterna.
Och han sade till konungen: »Så säger HERREN: Därför att du har släppt ur din hand den man som av mig var given till spillo, skall det gå dig såsom det skulle hava gått honom, och ditt folk såsom det har gått hans folk.»
Och Israels konung begav sig hem, missmodig och vred, och kom till Samaria.
Därefter hände sig följande.
Jisreeliten Nabot hade en vingård i Jisreel bredvid Ahabs palats, konungens i Samaria.
Och Ahab talade till Nabot och sade: »Låt mig få din vingård för att därav göra mig en köksträdgård, eftersom den ligger så nära intill mitt hus; jag vill giva dig en bättre vingård i stället, eller om dig så behagar, vill jag giva dig penningar såsom betalning för den.»
Men Nabot svarade Ahab: »HERREN låte det vara fjärran ifrån mig att jag skulle låta dig få mina fäders arvedel.»
Då gick Ahab hem till sitt, missmodig och vred för det svars skull som jisreeliten Nabot hade givit honom, när denne sade: »Jag vill icke låta dig få mina fäders arvedel.»
Och han lade sig på sin säng och vände bort sitt ansikte och åt intet.
Då kom hans hustru Isebel in till honom och frågade honom: »Varför är du så missmodig, och varför äter du intet?»
Han svarade henne: »Därför att när jag talade till jisreeliten Nabot och sade till honom: 'Låt mig få din vingård för penningar, eller om du så önskar, vill jag giva dig en annan vingård i stället', då svarade han: 'Jag vill icke låta dig få min vingård.'
Då sade hans hustru Isebel honom: »Är det du som nu regerar över Israel?
Stå upp och ät och var vid gott mod; jag skall skaffa dig jisreeliten Nabot vingård.
Därefter skrev hon ett brev i Ahabs namn och satte sigill under det med hans signetring, och sände så brevet till de äldste och förnämsta i Nabots stad, de som bodde där jämte honom.
Och hon skrev i brevet så: »Lysen ut en fasta, och låten Nabot sitta längst fram bland folket.
Och låten så två onda män sätta sig mitt emot honom, och låten dem vittna emot honom och säga: 'Du har talat förgripligt mot Gud och konungen.'
Fören så ut honom och stenen honom till döds.»
Och de äldsta och förnämsta männen i staden, de som bodde där i hans stad, handlade i enlighet med det bud som Isebel hade sänt dem, och såsom det var skrivet i brevet som hon hade sänt till dem.
De lyste ut en fasta och läto Nabot sitta längst fram bland folket.
Och de två onda männen kommo och satte sig mitt emot honom; och de onda männen vittnade mot Nabot inför folket och sade: Nabot har talat förgripligt mot Gud och konungen.»
Då förde man honom utanför staden och stenade honom till döds.
Därefter sände de bud till Isebel och läto säga: »Nabot har blivit stenad till döds.»
Så snart Isebel hörde att Nabot var stenad till döds, sade hon till Ahab: »Stå upp och tag jisreeliten Nabots vingård i besittning, den som han vägrade att låta dig få för penningar; ty Nabot är icke längre vid liv, utan han är död.»
Så snart Ahab hörde att Nabot var död, stod han upp och begav sig åstad ned till jisreeliten Nabots vingård för att taga den i besittning.
Men HERRENS ord kom till tisbiten Elia; han sade:
»Stå upp, gå åstad och möt Ahab, Israels konung, som bor i Samaria.
Du träffar honom i Nabots vingård, dit han har gått ned för att taga den i besittning.
Och du skall tala till honom och säga: 'Så säger HERREN: Har du till redan hunnit att både dräpa och tillträda arvet?'
Därefter skall du tala till honom och säga: 'Så säger HERREN: På samma ställe där hundarna hava slickat Nabots blod skola hundarna slicka också ditt blod.'»
Ahab sade till Elia: »Har du äntligen funnit mig, du min fiende?»
Han svarade: »Ja, jag har funnit dig.
Eftersom du har sålt dig till att göra vad ont är i HERRENS ögon,
därför skall jag ock låta vad ont är komma över dig och skall bortsopa dig, och av Ahabs hus skall jag utrota allt mankön, både små och stora i Israel.
Och jag skall göra med ditt hus såsom jag gjorde med Jerobeams, Nebats sons, hus, och såsom jag gjorde med Baesas, Ahias sons, hus, därför att du har förtörnat mig och kommit Israel att synda.
Också om Isebel har HERREN talat och sagt: Hundarna skola äta upp Isebel invid Jisreels murar.
Ja, den av Ahabs hus, som dör i staden, skola hundarna äta upp, och den som dör ute på marken skola himmelens fåglar äta upp.»
(Också har ingen varit såsom Ahab, han som sålde sig till att göra vad ont var i HERRENS ögon, när hans hustru Isebel uppeggade honom därtill.
Mycken styggelse förövade han, i det han följde efter de eländiga avgudarna, alldeles såsom amoréerna hade gjort, vilka HERREN fördrev för Israels barn.)
Men när Ahab hörde de orden, rev han sönder sina kläder och svepte säcktyg om sin kropp och fastade; och han låg höljd i säcktyg och gick tyst omkring.
Då kom HERRENS ord till tisbiten Elia; han sade:
»Har du sett huru Ahab ödmjukar sig inför mig?
Därför att han så ödmjukar sig inför mig, skall jag icke låta olyckan komma i hans tid; först i hans sons tid skall jag låta olyckan komma över hans hus.»
Och de sutto i ro i tre år, under vilka intet krig var mellan Aram och Israel.
Men i det tredje året for Josafat, Juda konung, ned till Israels konung.
Och Israels konung sade till sina tjänare: »I veten ju att Ramot i Gilead tillhör oss.
Och likväl sitta vi stilla och taga det icke ifrån konungen i Aram.»
Och han frågade Josafat: Vill du draga med mig för att belägra Ramot i Gilead?»
Josafat svarade Israels konung: »Jag såsom du, mitt folk såsom ditt folk, mina hästar såsom dina hästar!»
Men Josafat sade ytterligare till Israels konung: »Fråga dock först HERREN härom.»
Då församlade Israels konung profeterna, vid pass fyra hundra män, och frågade dem: »Skall jag draga åstad mot Ramot i Gilead för att belägra det, eller skall jag avstå därifrån?»
De svarade: »Drag ditupp; Herren skall giva det i konungens hand.»
Men Josafat sade: »Finnes här ingen annan HERRENS profet, så att vi kunna fråga genom honom?»
Israels konung svarade Josafat: »Här finnes ännu en man, Mika, Jimlas son, genom vilken vi kunna fråga HERREN; men han är mig förhatlig, ty han profeterar aldrig lycka åt mig, utan allenast olycka.»
Josafat sade: »Konungen säge icke så.»
Då kallade Israels konung till sig en hovman och sade: »Skaffa skyndsamt hit Mika, Jimlas son.»
Israels konung och Josafat, Juda konung, sutto nu var och en på sin tron, iklädda sina skrudar, på en tröskplats vid Samarias port, under det att alla profeterna profeterade inför dem.
Då gjorde sig Sidkia, Kenaanas son, horn av järn och sade: »Så säger HERREN: Med dessa skall du stånga araméerna, så att de förgöras.»
Och alla profeterna profeterade på samma sätt och sade: »Drag upp mot Ramot i Gilead, så skall du bliva lyckosam; HERREN skall giva det i konungens hand.»
Och budet som hade gått för att tillkalla Mika talade till honom och sade: »Det är så, att profeterna med en mun lova konungen lycka; låt nu dina ord stämma överens med vad de hava talat, och lova också du lycka.»
Men Mika svarade: »Så sant HERREN lever, jag skall allenast tala det som HERREN säger till mig.»
När han sedan kom till konungen, frågade konungen honom: »Mika, skola vi draga åstad till Ramot i Gilead för att belägra det, eller skola vi avstå därifrån?»
Han svarade honom: »Drag ditupp, så skall du bliva lyckosam; HERREN skall giva det i konungens hand.»
Men konungen sade till honom: »Huru många gånger skall jag besvärja dig att icke tala till mig annat än sanning i HERRENS namn?»
Då sade han: »Jag såg hela Israel förskingrat på bergen, likt får som icke hava någon herde.
Och HERREN sade: 'Dessa hava icke någon herre; må de vända tillbaka hem i frid, var och en till sitt.'»
Då sade Israels konung till Josafat: »Sade jag dig icke att denne aldrig profeterar lycka åt mig, utan allenast olycka?»
Men han sade: »Hör alltså HERRENS ord.
Jag såg HERREN sitta på sin tron och himmelens hela härskara stå där hos honom, på hans högra sida och på hans vänstra.
Och HERREN sade: 'Vem vill locka Ahab att draga upp mot Ramot i Gilead, för att han må falla där?'
Då sade den ene så och den andre så.
Slutligen kom anden fram och ställde sig inför HERREN och sade: 'Jag vill locka honom därtill.'
HERREN frågade honom: 'På vad sätt?'
Han svarade: 'Jag vill gå ut och bliva en lögnens ande i alla hans profeters mun.'
Då sade han: 'Du må försöka att locka honom därtill, och du skall också lyckas; gå ut och gör så.'
Och se, nu har HERREN lagt en lögnens ande i alla dessa dina profeters mun, medan HERREN ändå har beslutit att olycka skall komma över dig.»
Då trädde Sidkia, Kenaanas son, fram och gav Mika ett slag på kinden och sade: »På vilken väg har då HERRENS Ande gått bort ifrån mig för att tala med dig?»
Mika svarade: »Du skall få se det på den dag då du nödgas springa från kammare till kammare för att gömma dig.»
Men Israels konung sade: »Tag Mika och för honom tillbaka till Amon, hövitsmannen i staden, och till Joas, konungasonen.
Och säg: Så säger konungen: Sätten denne i fängelse och bespisen honom med fångkost, till dess jag kommer välbehållen hem.»
Mika svarade: »Om du kommer välbehållen tillbaka, så har HERREN icke talat genom mig.»
Och han sade ytterligare: »Hören detta, I folk, allasammans.»
Så drog nu Israels konung jämte Josafat, Juda konung, upp till Ramot i Gilead.
Och Israels konung sade till Josafat: »Jag vill förkläda mig, när jag drager ut i striden, men du må vara klädd i dina egna kläder.»
Så förklädde sig Israels konung, när han drog ut i striden.
Men konungen i Aram hade bjudit och sagt till sina trettiotvå vagnshövitsmän: »I skolen icke giva eder i strid med någon, vare sig liten eller stor, utom med Israels konung allena.»
När då hövitsmännen över vagnarna fingo se Josafat, tänkte de: »Förvisso är detta Israels konung», och vände sig därför till anfall mot honom.
Då gav Josafat upp ett rop.
Så snart nu hövitsmännen över vagnarna märkte att det icke var Israels konung, vände de om och läto honom vara.
Men en man som spände sin båge och sköt på måfå träffade Israels konung i en fog på rustningen.
Då sade denne till sin körsven: »Sväng om vagnen och för mig ut ur hären, ty jag är sårad.»
Och striden blev på den dagen allt häftigare, och konungen stod upprätt i sin vagn, vänd mot araméerna; men om aftonen gav han upp andan.
Och blodet från såret hade runnit ned i vagnen.
Och vid solnedgången gick ett rop genom hären: »Var och en till sin stad igen!
Var och en till sitt land igen!»
Så dödades då konungen och blev förd till Samaria; och man begrov konungen där i Samaria.
Och när man sköljde vagnen i dammen i Samaria, slickade hundarna hans blod, och skökorna badade sig däri -- såsom HERREN hade sagt.
Vad nu mer är att säga om Ahab och om allt vad han gjorde, om elfenbenshuset som han byggde, och om alla de städer som han byggde, det finnes upptecknat i Israels konungars krönika.
Och Ahab gick till vila hos sina fäder.
Och hans son Ahasja blev konung efter honom.
Men Josafat, Asas sons blev konung över Juda i Ahabs, Israels konungs, fjärde regeringsår.
Trettiofem år gammal var Josafat, när han blev konung, och han regerade tjugufem år i Jerusalem.
Hans moder hette Asuba, Silhis dotter.
Och han vandrade i allt på sin fader Asas väg, utan att vika av ifrån den; han gjorde nämligen vad rätt var i HERRENS ögon.
Dock blevo offerhöjderna icke avskaffade, utan folket fortfor att frambära offer och tända offereld på höjderna.
Och Josafat höll fred med Israels konung.
Vad nu mer är att säga om Josafat och om de bedrifter han utförde och om hans krig, det finnes upptecknat i Juda konungars krönika.
Han utrotade ock ur landet de tempelbolare som ännu funnos där, vilka hade lämnats kvar i hans fader Asas tid.
I Edom fanns då ingen konung, utan en ståthållare regerade där.
Och Josafat hade låtit bygga Tarsis-skepp, som skulle gå till Ofir för att hämta guld; men de kommo aldrig åstad, ty de ledo skeppsbrott vid Esjon-Geber.
Då sade Ahasja, Ahabs son, till Josafat: »Låt mitt folk fara med ditt folk på skeppen.»
Men Josafat ville icke.
Och Josafat gick till vila hos sina fäder och blev begraven hos sina fäder i sin fader Davids stad.
Och hans son Joram blev konung efter honom.
Ahasja, Ahabs son, blev konung över Israel i Samaria i Josafats, Juda konungs, sjuttonde regeringsår, och han regerade över Israel i två år.
Han gjorde vad ont var i HERRENS ögon och vandrade på sin faders och sin moders väg och på Jerobeams, Nebats sons, väg, hans som hade kommit Israel att synda.
Och han tjänade Baal och tillbad honom och förtörnade HERREN, Israels Gud, alldeles såsom hans fader hade gjort.
Efter Ahabs död avföll Moab från Israel.
Och Ahasja störtade ned genom gallret i sin Övre sal i Samaria och skadade sig, så att han blev sjuk.
Då skickade han åstad sändebud och sade till dem: »Gån och frågen Baal-Sebub, guden i Ekron, om jag skall tillfriskna från denna sjukdom.»
Men HERRENS ängel hade talat så till tisbiten Elia: »Stå upp och gå emot konungens i Samaria sändebud och tala så till dem: 'Är det därför att ingen Gud finnes i Israel som I gån åstad och frågen Baal-Sebub, guden i Ekron?
Därför att I gören detta, säger HERREN så: Du skall icke komma upp ur den säng i vilken du har lagt dig, ty du skall döden dö.'»
Och Elia gick.
När sedan sändebuden kommo tillbaka till konungen, frågade han dem: »Varför kommen I tillbaka?»
De svarade honom: »En man kom emot oss och sade till oss: 'Gån tillbaka till konungen, som har sänt eder, och talen så till honom: Så säger HERREN: Är det därför att ingen Gud finnes i Israel som du sänder bud för att fråga Baal-Sebub, guden i Ekron?
Därför att du så gör skall du icke komma upp ur den säng i vilken du har lagt dig, ty du skall döden dö.'»
Då frågade han dem: »Huru såg den mannen ut, som kom emot eder och talade till eder på detta sätt?»
De svarade honom: »Mannen bar en hårmantel och var omgjordad med en lädergördel om sina länder.»
Då sade han: »Det var tisbiten Elia.»
Och han sände till honom en underhövitsman med femtio man.
Och när denne kom upp till honom, där han satt på toppen av berget, sade han till honom: »Du gudsman, konungen befaller dig att komma ned.»
Men Elia svarade och sade till underhövitsmannen: »Om jag är en gudsman, så komme eld ned från himmelen och förtäre dig och dina femtio.»
Då kom eld ned från himmelen och förtärde honom och hans femtio.
Och han sände åter till honom en annan underhövitsman med femtio man.
Denne tog till orda och sade till honom: »Du gudsman, så säger konungen: Kom strax ned.»
Men Elia svarade och sade till dem: »Om jag är en gudsman, så komme eld ned från himmelen och förtäre dig och dina femtio.»
Då kom Guds eld ned från himmelen och förtärde honom och hans femtio.
Åter sände han åstad en tredje underhövitsman med femtio man Och denne tredje underhövitsman drog ditupp, och när han kom fram, föll han ned på sina knän för Elia och bad honom och sade till honom: »Du gudsman, låt mitt liv och dessa dina femtio tjänares liv vara något aktat i dina ögon.
Se, eld har kommit ned från himmelen och förtärt de första två underhövitsmännen med deras femtio man; men låt nu mitt liv vara något aktat i dina ögon.
Och HERRENS ängel sade till Elia: »Gå ned med honom, frukta icke för honom.»
Då stod han upp och gick med honom ned till konungen
Och han sade till denne: »Så säger HERREN: Eftersom du skickade sändebud för att fråga Baal-Sebub, guden i Ekron -- likasom om i Israel icke funnes någon Gud, som du kunde fråga härom -- fördenskull skall du icke få komma upp ur den säng i vilken du har lagt dig, ty du skall döden dö.»
Och han dog, i enlighet med det HERRENS ord som Elia hade talat; och Joram blev konung efter honom, i Jorams, Josafats sons, Juda konungs, andra regeringsår.
Han hade nämligen ingen son.
Vad nu mer är att säga om Ahasja, om vad han gjorde, det finnes upptecknat i Israels konungars krönika.
Vid den tid då HERREN ville upptaga Elia till himmelen i en stormvind gingo Elia och Elisa från Gilgal.
Och Elia sade till Elisa: »Stanna här, ty HERREN har sänt mig till Betel.»
Men Elisa svarade: »Så sant HERREN lever, och så sant du själv lever, jag lämnar dig icke.
Och de gingo ned till Betel.
Då kommo profetlärjungarna i Betel ut till Elisa och sade till honom: »Vet du att HERREN i dag vill taga din herre ifrån dig, upp över ditt huvud?»
Han svarade: »Ja, jag vet det; tigen stilla.»
Och Elia sade till honom: »Elisa, stanna här, ty HERREN har sänt mig till Jeriko.»
Men han svarade: »Så sant HERREN lever, och så sant du själv lever, jag lämnar dig icke.»
Och de kommo till Jeriko.
Då gingo profetlärjungarna i Jeriko fram till Elisa och sade till honom: »Vet du att HERREN i dag vill taga din herre ifrån dig, upp över ditt huvud?»
Han svarade: »Ja, jag vet det; tigen stilla.»
Och Elia sade till honom: »Stanna här, ty HERREN har sänt mig till Jordan.»
Men han svarade: »Så sant HERREN lever, och så sant du själv lever, jag lämnar dig icke.»
Och de gingo båda åstad.
Men femtio män av profetlärjungarna gingo ock åstad och ställde sig på något avstånd, längre bort, under det att de båda stodo vid Jordan.
Och Elia tog sin mantel och vek ihop den och slog på vattnet; då delade sig detta åt två sidor.
Och de gingo så båda på torr mark därigenom.
När de hade kommit över, sade Elia till Elisa: »Bed mig om vad jag skall göra för dig, innan jag bliver tagen ifrån dig.»
Elisa sade »Må en dubbel arvslott av din ande falla mig till.»
Han svarade: »Du har bett om något svårt.
Men om du ser mig, när jag bliver tagen ifrån dig, då kommer det dock att så ske dig; varom icke, så sker det ej.»
Under det att de nu gingo och talade, syntes plötsligt en vagn eld, med hästar av eld, och skilde de båda från varandra; och Elia for i stormvinden upp till himmelen.
Och Elisa såg det och ropade: »Min fader, min fader!
Du som för Israel är både vagnar och ryttare!»
Sedan såg han honom icke mer.
Och han fattade i sina kläder och rev sönder dem i två stycken.
Därefter tog han upp Elias mantel, som hade fallit av denne, och vände så om och ställde sig vid Jordans strand.
Och han tog Elias mantel, som hade fallit av denne, och slog på vattnet och sade: »Var är HERREN, Elias Gud?»
Då nu också Elisa slog på vattnet, delade det sig åt två sidor, och han gick över.
När profetlärjungarna, som voro vid Jeriko på något avstånd, sågo detta, sade de: »Elias ande vilar på Elisa.»
Och de kommo honom till mötes och bugade sig ned till jorden för honom.
Och de sade till honom: »Se, bland dina tjänare finnas femtio raska män; låt dessa gå och söka efter din herre.
Kanhända har HERRENS Ande lyft upp honom och kastat honom på något berg eller i någon dal.»
Men han svarade: »Sänden ingen åstad.
Men när de länge och väl enträget hade bett honom därom, sade han: »Så sänden då åstad.»
Då sände de åstad femtio män; och dessa sökte efter honom i tre dagar, men funno honom icke.
När de sedan kommo tillbaka till honom, medan han ännu vistades i Jeriko, sade han till dem: »Sade jag icke till eder att I icke skullen gå?»
Och männen i staden sade till Elisa: »Stadens läge är ju gott, såsom min herre ser, men vattnet är dåligt, och därav komma missfall i landet.»
Han sade: »Hämten hit åt mig en ny skål och läggen salt däri.»
Och de hämtade en åt honom.
Därefter gick han ut till vattenkällan och kastade salt däri och sade: »Så säger HERREN: Jag har nu gjort detta vatten sunt; död och missfall skola icke mer komma därav.
Och vattnet blev sunt, och har förblivit så ända till denna dag, i enlighet med det ord Elisa talade.
Därifrån begav han sig upp till Betel.
Och under det han var på väg ditupp, kom en skara gossar ut ur staden; och de begynte driva gäck med honom och ropade till honom: »Upp med dig, du flintskalle!
Upp med dig, du flintskalle!»
När han då vände sig om och fick se dem, uttalade han en förbannelse över dem i HERRENS namn.
Då kommo två björninnor ut ur skogen och sleto sönder fyrtiotvå av barnen.
Därifrån gick han till berget Karmel och vände sedan därifrån tillbaka till Samaria.
Joram, Ahabs son, blev konung över Israel i Samaria i Josafats, Juda konungs, adertonde regeringsår, och han regerade i tolv år.
Han gjorde vad ont var i HERRENS ögon; dock icke såsom hans fader och moder, ty han skaffade bort den Baalsstod som hans fader hade låtit göra.
Dock höll han fast vid de Jerobeams, Nebats sons, synder genom vilka denne hade kommit Israel att synda; från dessa avstod han icke.
Mesa, konungen i Moab, som ägde mycken boskap, hade i skatt till konungen i Israel erlagt hundra tusen lamm och ull av hundra tusen vädurar.
Men när Ahab var död, avföll konungen i Moab från konungen i Israel.
Då drog konung Joram ut från Samaria och mönstrade hela Israel.
Därefter sände han åstad bud till Josafat, konungen i Juda, och lät säga honom: »Konungen i Moab har avfallit från mig.
Vill du draga med mig för att strida mot Moab?»
Han svarade: »Ja, jag vill draga ditupp -- jag såsom du, mitt folk såsom ditt folk, mina hästar såsom dina hästar!»
Och han frågade: »Vilken väg skola vi draga ditupp?»
Han svarade »Vägen genom Edoms öken.»
Så drogo då konungen i Israel konungen i Juda och konungen i Edom åstad; men när de hade färdats sju dagsresor, fanns intet vatten för hären och för djuren som de hade med sig.
Då sade Israels konung: »Ack att HERREN skulle kalla tillhopa dessa tre konungar för att giva dem i Moabs hand!»
Men Josafat sade: »Finnes här ingen HERRENS profet, så att vi kunna fråga HERREN genom honom?»
Då svarade en av Israels konungs tjänare och sade: »Elisa, Safats son, finnes här, han som plägade gjuta vatten på Elias händer.»
Josafat sade: »Hos honom är HERRENS ord.»
Israels konung och Josafat och Edoms konung gingo då ned till honom.
Men Elisa sade till Israels konung: »Vad har du med mig att göra?
Gå du till din faders profeter och till din moders profeter.»
Israels konung svarade honom: »Bort det, att HERREN skulle hava kallat tillhopa dessa tre konungar för att giva dem i Moabs hand!»
Då sade Elisa: »Så sant HERREN Sebaot lever, han vilkens tjänare jag är: om jag icke hade undseende för Josafat, Juda konung, så skulle jag icke akta på dig eller se till dig.
Men hämten nu hit åt mig en harpospelare.»
Så ofta harpospelaren spelade, kom nämligen HERRENS hand över honom.
Och han sade: »Så säger HERREN: Gräven i denna dal grop vid grop.
Ty så säger HERREN: I skolen icke märka någon vind, ej heller se något regn, men likväl skall denna dal bliva full med vatten, så att både I själva skolen hava att dricka och eder boskap och edra övriga djur.
Dock anser HERREN icke ens detta vara nog, utan han vill ock giva Moab i eder hand.
Och I skolen intaga alla befästa städer och alla andra ansenliga städer, I skolen fälla alla nyttiga träd och kasta igen alla vattenkällor, och alla bördiga åkerstycken skolen I fördärva med stenar.»
Och se, om morgonen, vid den tid då spisoffret frambäres, strömmade vatten till från Edomssidan, så att landet fylldes med vatten.
Moabiterna hade nu allasammans hört att konungarna hade dragit upp för att strida mot dem, och alla de som voro vid vapenför ålder eller därutöver blevo uppbådade och stodo nu vid gränsen.
Men bittida om morgonen, när solen gick upp och lyste på vattnet, sågo moabiterna vattnet framför sig rött såsom blod.
Då sade de: »Det är blod!
Konungarna hava helt visst råkat i strid och därvid dräpt varandra.
Nu till plundring, Moab!»
Men när de kommo till Israels läger, bröto israeliterna fram och slogo moabiterna, så att de flydde för dem.
Och de drogo in i landet och slogo ytterligare moabiterna.
Och städerna förstörde de, och på alla bördiga åkerstycken kastade de var och en sin sten, till dess de hade överhöljt dem, och alla vattenkällor täppte de till, och alla nyttiga träd fällde de, så att de till slut lämnade kvar allenast stenarna av Kir-Hareset.
Men när slungkastarna omringade staden och besköto den
och Moabs konung såg att han icke kunde hålla stånd i striden, tog han med sig sju hundra svärdbeväpnade män för att slå sig igenom till Edoms konung; men de kunde det icke.
Då tog han sin förstfödde son, den som skulle bliva konung efter honom, och offrade denne på muren till ett brännoffer.
Då drabbades Israel av svår hemsökelse, så att de måste bryta upp och lämna honom i fred och vända tillbaka till sitt land igen.
Och en kvinna som var hustru till en av profetlärjungarna ropade till Elisa och sade: »Min man, din tjänare, har dött, och du vet att din tjänare fruktade HERREN; nu kommer hans fordringsägare och vill taga mina båda söner till trälar.
Elisa sade till henne: »Vad kan jag göra för dig?
Säg mig, vad har du i huset?»
Hon svarade: »Din tjänarinna har intet annat i huset än en flaska smörjelseolja.»
Då sade han: »Gå och låna dig kärl utifrån av alla dina grannar, tomma kärl, men icke för få.
Gå så in, och stäng igen dörren om dig och dina söner, och gjut i alla dessa kärl; och när ett kärl är fullt, så flytta undan det.»
Då gick hon ifrån honom.
Och sedan hon hade stängt igen dörren om sig och sina söner, buro de fram kärlen till henne, och hon göt i.
Och när kärlen voro fulla, sade hon till sin son: »Bär fram åt mig ännu ett kärl.»
Men han svarade henne: »Här finnes intet kärl mer.
Då stannade oljan av.
Och hon kom och berättade detta för gudsmannen.
Då sade han: »Gå och sälj oljan, och betala din skuld.
Sedan må du med dina söner leva av det som bliver över.»
En dag kom Elisa över till Sunem.
Där bodde en rik kvinna, som nödgade honom att äta hos sig; och så ofta han sedan kom ditöver, tog han in där och åt.
Då sade hon en gång till sin man: »Se, jag har förnummit att han som beständigt kommer hitöver är en helig gudsman.
Så låt oss nu mura upp ett litet rum på taket och där sätta in åt honom en säng, ett bord, en stol och en ljusstake, så att han kan få taga in där, när han kommer till oss.»
Så kom han dit en dag och fick då taga in i rummet och ligga där.
Och han sade till sin tjänare Gehasi: »Kalla hit sunemitiskan.»
Då kallade han dit henne, och hon infann sig där hos tjänaren.
Ytterligare tillsade han honom: »Säg till henne: 'Se, du har haft allt detta besvär för oss.
Vad kan nu jag göra för dig?
Har du något att andraga hos konungen eller hos härhövitsmannen?'»
Men hon svarade: »Nej; jag bor ju här mitt ibland mitt folk.»
Sedan frågade han: »Vad kan jag då göra för henne?»
Gehasi svarade: »Jo, hon har ingen son, och hennes man är gammal.»
Så sade han då: »Kalla henne hitin.»
Då kallade han dit henne, och hon stannade i dörren.
Och han sade: »Nästa år vid just denna tid skall du hava en son i famnen.»
Hon svarade: »Nej, min herre, du gudsman, inbilla icke din tjänarinna något sådant.»
Men kvinnan blev havande och födde en son följande år, just vid den tid som Elisa hade sagt henne.
Och när gossen blev större, hände sig en dag att han gick ut till sin fader hos skördemännen.
Då begynte han klaga för sin fader: »Mitt huvud!
Mitt huvud!»
Denne sade till sin tjänare: »Tag honom och bär honom till hans moder.
Han tog honom då och förde honom till hans moder.
Och han satt i hennes knä till middagstiden; då gav han upp andan.
Men hon gick upp och lade honom på gudsmannens säng och stängde igen om honom och gick ut.
Därefter kallade hon på sin man och sade: »Sänd till mig en av tjänarna med en åsninna, så vill jag skynda till gudsmannen; sedan kommer jag strax tillbaka.»
Han sade: »Varför vill du i dag fara till honom?
Det är ju varken nymånad eller sabbat.»
Hon svarade: »Oroa dig icke!»
Sedan lät hon sadla åsninnan och sade till sin tjänare: »Driv på framåt, och gör icke något uppehåll i min färd, förrän jag säger dig till.»
Så begav hon sig åstad och kom till gudsmannen på berget Karmel.
Då nu gudsmannen fick se henne på något avstånd, sade han till sin tjänare Gehasi: »Se, där är sunemitiskan.
Skynda nu emot henne och fråga henne: 'Allt står väl rätt till med dig och med din man och med gossen?'»
Hon svarade: »Ja.»
Men när hon kom upp till gudsmannen på berget, fattade hon om hans fötter.
Då gick Gehasi fram och ville driva henne undan; men gudsmannen sade: »Låt henne vara, ty hennes själ är bedrövad; men HERREN hade fördolt detta för mig och icke låtit mig få veta det.»
Och hon sade: »Hade jag väl bett min herre om en son?
Sade jag icke fastmer att du icke skulle inbilla mig något?»
Då sade han till Gehasi: »Omgjorda dina länder och tag min stav i din hand och gå åstad; om du möter någon, så hälsa icke på honom, och om någon hälsar på dig, så besvara icke hans hälsning.
Och lägg sedan min stav på gossens ansikte.»
Men gossens moder sade: »Så sant HERREN lever, och så sant du själv lever, jag släpper dig icke.»
Då stod han upp och följde med henne.
Men Gehasi hade redan gått före dem och lagt staven på gossens ansikte; dock hördes icke ett ljud, och intet spår av förnimmelse kunde märkas.
Då vände han om och gick honom till mötes och berättade det för honom och sade: »Gossen har icke vaknat upp.»
Och när Elisa kom in i huset, fick han se att gossen låg död på hans säng.
Då gick han in och stängde igen dörren om dem båda och bad till HERREN.
Och han steg upp i sängen och lade sig över gossen, så att han hade sin mun på hans mun, sina ögon på hans ögon och sina händer på hans händer.
När han så lutade sig ned över gossen, blev kroppen varm.
Därefter gick han åter fram och tillbaka i rummet och steg så åter upp i sängen och lutade sig ned över honom.
Då nös gossen, ända till sju gånger.
Och därpå slog gossen upp ögonen.
Sedan ropade han på Gehasi och sade: »Kalla hit sunemitiskan.»
Då kallade han in henne, och när hon kom in till honom, sade han: »Tag din son.»
Då kom hon fram och föll ned för hans fötter och bugade sig mot jorden.
Därefter tog hon sin son och gick ut.
Och Elisa kom åter till Gilgal, medan hungersnöden var i landet.
När då profetlärjungarna sutto där inför honom, sade han till sin tjänare »Sätt på den stora grytan och koka något till soppa åt profetlärjungarna.»
Och en av dem gick ut på marken för att plocka något grönt; då fick han se en vild slingerväxt, och av den plockade han något som liknade gurkor, sin mantel full.
När han sedan kom in, skar han sönder dem och lade dem i soppgrytan; ty de kände icke till dem.
Och de öste upp åt männen, för att de skulle äta.
Men så snart de hade begynt äta av soppan, gåvo de upp ett rop och sade: »Döden är i grytan, du gudsman!»
Och de kunde icke äta.
Då sade han: »Skaffen hit mjöl.»
Detta kastade han i grytan.
Därefter sade han: »Ös upp åt folket och låt dem äta.»
Och intet skadligt fanns nu mer i grytan.
Och en man kom från Baal-Salisa och förde med sig åt gudsmannen förstlingsbröd; tjugu kornbröd, och ax av grönskuren säd i sin påse.
Då sade han: »Giv det åt folket att äta.»
Men hans tjänare sade: »Huru skall jag kunna sätta fram detta för hundra män?»
Han sade: »Giv det åt folket att äta; ty så säger HERREN: De skola äta och få över.
Då satte han fram det för dem.
Och de åto och fingo över, såsom HERREN hade sagt.
Naaman, den arameiske konungens härhövitsman, hade stort anseende hos sin herre och var högt aktad, ty genom honom hade HERREN givit seger åt Aram; och han var en tapper stridsman, men spetälsk.
Nu hade araméerna, en gång då de drogo ut på strövtåg, fört med sig såsom fånge ur Israels land en ung flicka, som kom i tjänst hos Naamans hustru.
Denna sade till sin fru: »Ack att min herre vore hos profeten i Samaria, så skulle denne nog befria honom från hans spetälska!»
Då gick hon åstad och berättade detta för sin herre och sade: »Så och så har flickan ifrån Israels land sagt.
Konungen i Aram svarade: »Far dit, så skall jag sända brev till konungen i Israel.»
Så for han då och tog med sig tio talenter silver och sex tusen siklar guld, så ock tio högtidsdräkter.
Och han överlämnade brevet till Israels konung, och däri stod det: »Nu, när detta brev kommer dig till handa, må du veta att jag har sänt till dig min tjänare Naaman, för att du må befria honom från hans spetälska.»
När Israels konung hade läst brevet, rev han sönder sina kläder och sade: »Är jag då Gud, så att jag skulle kunna döda och göra levande, eftersom denne sänder bud till mig att jag skall befria en man från hans spetälska?
Märken nu och sen huru han söker sak med mig.»
Men när gudsmannen Elisa hörde att Israels konung hade rivit sönder sina kläder, sände han till konungen och lät säga: »Varför har du rivit sönder dina kläder?
Låt honom komma till mig, så skall han förnimma att en profet finnes i Israel.»
Så kom då Naaman med sina hästar och vagnar och stannade vid dörren till Elisas hus.
Då sände Elisa ett bud ut till honom och lät säga: »Gå bort och bada dig sju gånger i Jordan, så skall ditt kött åter bliva sig likt, och du skall bliva ren.»
Men Naaman blev vred och for sin väg, i det han sade: »Jag tänkte att han skulle gå ut till mig och träda fram och åkalla HERRENS, sin Guds, namn och föra sin hand fram och åter över stället och så taga bort spetälskan.
Äro icke Damaskus' floder, Abana och Parpar, bättre än alla vatten Israel?
Då kunde jag ju lika gärna bada mig i dem för att bliva ren.»
Så vände han om och for sin väg i vrede.
Men hans tjänare gingo fram och talade till honom och sade: »Min fader, om profeten hade förelagt dig något svårt, skulle du då icke hava gjort det?
Huru mycket mer nu, då han allenast har sagt till dig: 'Bada dig, så bliver du ren'!
Då for han ned och doppade sig i Jordan sju gånger, såsom gudsmannen hade sagt; och hans kött blev då åter sig likt, friskt såsom en ung gosses kött, och han blev ren.
Därefter vände han tillbaka till gudsmannen med hela sin skara och gick in och trädde fram för honom och sade: »Se, nu vet jag att ingen Gud finnes på hela jorden utom i Israel.
Så tag nu emot en tacksamhetsskänk av din tjänare.»
Men han svarade: »Så sant HERREN lever, han vilkens tjänare jag är, jag vill icke taga emot den.»
Och fastän han enträget bad honom att taga emot den, ville han icke.
Då sade Naaman: »Om du icke vill detta, så låt då din tjänare få så mycket jord som ett par mulåsnor kunna bära.
Ty din tjänare vill icke mer offra brännoffer och slaktoffer åt andra gudar, utan allenast åt HERREN.
Detta må dock HERREN förlåta din tjänare: när min herre går in i Rimmons tempel för att där böja knä, och han då stöder sig vid min hand, och jag också böjer knä där i Rimmons tempel, må då HERREN förlåta din tjänare, när jag så böjer knä i Rimmons tempel.
Han sade till honom: »Far i frid.»
Men när hän hade lämnat honom och farit ett stycke väg framåt,
tänkte Gehasi, gudsmannen Elisas tjänare: »Se, min herre har släppt denne Naaman från Aram, utan att taga emot av honom vad han hade fört med sig.
Så sant HERREN lever, jag vill skynda efter honom och söka få något av honom.»
Så gav sig då Gehasi åstad efter Naaman.
Men när Naaman såg någon skynda efter sig, steg han med hast ned från vagnen och gick emot honom och sade: »Allt står väl rätt till?»
Han svarade: »Ja; men min herre har sänt mig och låter säga: 'Just nu hava två unga män, profetlärjungar, kommit till mig från Efraims bergsbygd; giv dem en talent silver och två högtidsdräkter.'»
Naaman svarade: »Värdes taga två talenter.»
Och han bad honom enträget och knöt så in två talenter silver i två pungar och tog fram två högtidsdräkter, och lämnade detta åt två av sina tjänare, och dessa buro det framför honom.
Men när han kom till kullen, tog han det ur deras hand och lade det i förvar i huset; sedan lät han männen gå sin väg.
Därefter gick han in och trädde fram för sin herre.
Då frågade Elisa honom: »Varifrån kommer du, Gehasi?»
Han svarade: »Din tjänare har ingenstädes varit.»
Då sade han till honom: »Menar du att jag icke i min ande var med, när en man vände om från sin vagn och gick emot dig?
Är det nu tid att du skaffar dig silver och skaffar dig kläder, så ock olivplanteringar, vingårdar, får och fäkreatur, tjänare och tjänarinnor,
nu då Naamans spetälska kommer att låda vid dig och vid dina efterkommande för evigt?»
Så gick denne ut ifrån honom, vit såsom snö av spetälska.
Profetlärjungarna sade till Elisa: »Se, rummet där vi sitta inför dig är för trångt för oss.»
Låt oss därför gå till Jordan och därifrån hämta var sin timmerstock, så att vi där kunna bygga oss ett annat hus att sitta i.»
Han svarade: »Gån åstad.»
Men en av dem sade: »Värdes själv gå med dina tjänaren.»
Han varade: »Ja, jag skall gå med.»
Så gick han med dem.
Och när de kommo till Jordan, begynte de hugga ned träd.
Men under det att en av dem höll på att fälla en stock, föll yxjärnet i vattnet.
Då gav han upp ett rop och sade: »Ack, min herre, yxan var ju lånad.»
Gudsmannen frågade: »Var föll den i?»
Och han visade honom stället.
Då högg han av ett stycke trä och kastade det i där och fick så järnet att flyta upp.
Sedan sade han: »Tag nu upp det.»
Då räckte mannen ut sin hand och tog det.
Och konungen i Aram låg i krig med Israel.
Men när han rådförde sig med sina tjänare och sade: »På det och det stället vill jag lägra mig»,
då sände gudsmannen bud till Israels konung och lät säga: »Tag dig till vara för att tåga fram vid det stället, ty araméerna ligga där.»
Då sände Israels konung till det ställe som gudsmannen hade angivit för honom och varnat honom för; och han tog sig till vara där.
Detta skedde icke allenast en gång eller två gånger.
Häröver blev konungen i Aram mycket orolig; och han kallade till sig sina tjänare och sade till dem: »Kunnen I icke säga mig vem av de våra det är som håller med Israels konung?»
Då svarade en av hans tjänare: »Icke så, min herre konung; men Elisa, profeten i Israel, kungör för Israels konung vart ord som du talar i din sovkammare.»
Han sade: »Gån och sen till, var han finnes, så att jag kan sända åstad och gripa honom.»
Och man berättade för honom att han var i Dotan.
Då sände han dit hästar och vagnar och en stor här; och de kommo dit om natten och omringade staden.
När nu gudsmannens tjänare bittida om morgonen stod upp och gick ut, fick han se att en här hade lägrat sig runt omkring staden med hästar och vagnar.
Då sade tjänaren till honom: »Ack, min herre, huru skola vi nu göra?»
Han svarade: »Frukta icke; ty de som äro med oss äro flera än de som äro med dem.»
Och Elisa bad och sade: »HERRE, öppna hans ögon, så att han ser.»
Då öppnade HERREN tjänarens ögon, och han fick se att berget var fullt med hästar och vagnar av eld, runt omkring Elisa.
När de nu drogo ned mot honom, bad Elisa till HERREN och sade: »Slå detta folk med blindhet.»
Då slog han dem med blindhet, såsom Elisa bad.
Och Elisa sade till dem: »Detta är icke den rätta vägen eller den rätta staden.
Följen mig, så skall jag föra eder till den man som I söken.»
Därefter förde han dem till Samaria.
Men när de kommo till Samaria, sade Elisa: »HERRE, öppna dessas ögon, så att de se.»
Då öppnade HERREN deras ögon, och de fingo se att de voro mitt i Samaria.
När då Israels konung såg dem, sade han till Elisa: »Skall jag hugga ned dem, min fader, skall jag hugga ned dem?»
Han svarade: »Du skall icke hugga ned dem.
Du plägar ju icke ens hugga ned dem som du har tagit till fånga med svärd och båge.
Sätt fram för dem mat och dryck och låt dem äta och dricka, och låt dem sedan gå till sin herre igen»
Då tillredde han åt dem en stor måltid, och när de hade ätit och druckit, lät han dem gå; och de gingo till sin herre igen.
Sedan kommo icke vidare några arameiska strövskaror in i Israels land.
Därefter hände sig att Ben-Hadad, konungen i Aram, samlade hela sin här och drog upp och belägrade Samaria.
Och medan de belägrade Samaria, uppstod där en så stor hungersnöd, att man betalade åttio siklar silver för ett åsnehuvud och fem siklar silver för en fjärdedels kab duvoträck.
Och en gång då Israels konung gick omkring på muren ropade en kvinna till honom och sade: »Hjälp, min herre konung!»
Han svarade: »Hjälper icke HERREN dig, varifrån skall då jag kunna skaffa hjälp åt dig?
Från logen eller från vinpressen?»
Och konungen frågade henne: »Vad fattas dig?»
Hon svarade: »Kvinnan där sade till mig: 'Giv hit din son, så att vi få äta honom i dag, så skola vi äta min son i morgon.'
Så kokade vi min son och åto upp honom.
Nästa dag sade jag till henne: 'Giv nu hit din son, så att vi få äta honom.'
Men då gömde hon undan sin son.»
När konungen hörde kvinnans ord, rev han sönder sina kläder, där han gick på muren.
Då fick folket se att han hade säcktyg inunder, närmast kroppen.
Och han sade: »Gud straffe mig nu och framgent, om Elisas, Safats sons, huvud i dag får sitta kvar på honom.»
Så sände han då dit en man före sig, under det att Elisa satt i sitt hus och de äldste sutto där hos honom.
Men innan den utskickade hann fram till honom, sade han till de äldste: »Sen I huru denne mördarson sänder hit en man för att taga mitt huvud?
Men sen nu till, att I stängen igen dörren, när den utskickade kommer; och spärren så vägen för honom med den.
Jag hör nu ock ljudet av hans herres steg efter honom.»
Medan han ännu talade med dem, kom den utskickade ned till honom.
Och denne sade: »Se, detta är en olycka som kommer från HERREN; huru skall jag då längre kunna hoppas på HERREN?»
Men Elisa svarade: »Hören HERRENS ord.
Så säger HERREN: I morgon vid denna tid skall man få ett sea-mått fint mjöl för en sikel, så ock två sea-mått korn för en sikel, i Samarias port.»
Den kämpe vid vilkens hand konungen stödde sig svarade då gudsmannen och sade: »Om HERREN också gjorde fönster på himmelen, huru skulle väl detta kunna ske?»
Han sade: »Du skall få se det med egna ögon, men du skall icke få äta därav.»
Utanför stadsporten uppehöllo sig då fyra spetälska män.
Dessa sade till varandra: »Varför skola vi stanna kvar här, till dess vi dö?»
Om vi besluta oss för att gå in i staden nu då hungersnöd är i staden, så skola vi dö där, och om vi stanna här, skola vi ock dö.
Välan då, låt oss gå över till araméernas läger; låta de oss leva, så få vi leva, och döda de oss, så må vi dö.»
Så stodo de då upp i skymningen för att gå in i araméernas läger.
Men när de kommo till utkanten av araméernas läger, se, då fanns ingen människa där.
Ty Herren hade låtit ett dån av vagnar och hästar höras i araméernas läger, ett dån såsom av en stor här, så att de hade sagt till varandra: »Förvisso har Israels konung lejt hjälp mot oss av hetiternas och egyptiernas konungar, för att dessa skola komma över oss.»
Därför hade de brutit upp och flytt i skymningen och hade övergivit sina tält, sina hästar och åsnor, lägret sådant det stod; de hade flytt för att rädda sina liv.
När de spetälska nu kommo till utkanten av lägret, gingo de in i ett tält och åto och drucko, och togo därur silver och guld och kläder, och gingo så bort och gömde det.
Sedan vände de tillbaka och gingo in i ett annat tält och togo vad där fanns, och gingo så bort och gömde det.
Men därefter sade de till varandra: »Vi bete oss icke rätt.
I dag kunna vi frambära ett glädjebudskap.
Men om vi nu tiga och vänta till i morgon, när det bliver dager, så skall det tillräknas oss såsom missgärning.
Välan då, låt oss gå och berätta detta i konungens hus.
Så gingo de åstad och ropade an vakten vid stadsporten och berättade för dem och sade: »Vi kommo till araméernas läger, men där fanns ingen människa, och icke ett ljud av någon människa hördes; där stodo allenast hästarna och åsnorna bundna och tälten såsom de pläga stå.»
Detta ropades sedan ut av dem som höllo vakt vid porten, och man förkunnade det också inne i konungens hus.
Konungen stod då upp om natten och sade till sina tjänare: »Jag vill säga eder vad araméerna hava för händer mot oss.
De veta att vi lida hungersnöd, därför hava de gått ut ur lägret och gömt sig ute på marken, i det de tänka att de skola gripa oss levande, när vi nu gå ut ur staden, och att de så skola komma in i staden.»
Men en av hans tjänare svarade och sade: »Låt oss taga fem av de återstående hästarna, dem som ännu finnas kvar härinne -- det skall ju eljest gå dem såsom det går hela hopen av israeliter som ännu äro kvar härinne, eller såsom det har gått hela hopen av israeliter som redan hava omkommit -- och låt oss sända åstad och se efter.»
Så tog man då två vagnar med hästar för, och konungen sände dem åstad efter araméernas här och sade: »Faren åstad och sen efter.»
Dessa foro nu efter dem ända till Jordan; och se, hela vägen var full med kläder och andra saker som araméerna hade kastat ifrån sig, när de hastade bort.
Och de utskickade kommo tillbaka och berättade detta för konungen.
Då drog folket ut och plundrade Araméernas läger; och nu fick man ett sea-mått fint mjöl för en sikel och likaså två sea-mått korn för en sikel, såsom HERREN hade sagt.
Och den kämpe vid vilkens hand konungen plägade stödja sig hade av honom blivit satt till att hålla ordning vid stadsporten; men folket trampade honom till döds i porten, detta i enlighet med gudsmannens ord, vad denne hade sagt, när konungen kom ned till honom.
Ty när gudsmannen sade till konungen: »I morgon vid denna tid skall man i Samarias port få två sea-mått korn för en sikel och likaså ett sea-mått fint mjöl för en sikel»,
då svarade kämpen gudsmannen och sade: »Om HERREN också gjorde fönster på himmelen, huru skulle väl något sådant kunna ske?»
Då sade han: »Du skall få se det med egna ögon, men du skall icke få äta därav.»
Så gick det honom ock, ty folket trampade honom till döds i porten.
Och Elisa talade till den kvinna vilkens son han hade gjort levande, han sade: »Stå upp och drag bort med ditt husfolk och vistas var du kan, ty HERREN har bjudit hungersnöden komma, och den har redan kommit in i landet och skall räcka i sju år.»
Då stod kvinnan upp och gjorde såsom gudsmannen sade; hon drog bort med sitt husfolk och vistades i filistéernas land i sju år.
Men när de sju åren voro förlidna, kom kvinnan tillbaka ifrån filistéernas land; och hon gick åstad för att anropa konungen om att återfå sitt hus och sin åker.
Och konungen höll då på att tala med Gehasi, gudsmannens tjänare, och sade: »Förtälj för mig alla de stora ting som Elisa har gjort.»
Och just som han förtäljde för konungen huru han hade gjort en död levande, då kom den kvinna vilkens son han hade gjort levande och anropade konungen om att återfå sitt hus och sin åker.
Då sade Gehasi: »Min herre konung, detta är kvinnan, och detta är hennes son, den som Elisa har gjort levande.»
Då frågade konungen kvinnan, och hon förtäljde allt för honom.
Sedan lät konungen henne få en hovman med sig och sade: »Skaffa tillbaka allt vad som tillhör henne, och därtill all avkastning av åkern, från den dag då hon lämnade landet ända till nu.»
Och Elisa kom till Damaskus, under det att Ben-Hadad, konungen i Aram, låg sjuk.
När man nu berättade för denne att gudsmannen hade kommit dit,
sade konungen till Hasael: »Tag skänker med dig och gå gudsmannen till mötes, och fråga HERREN genom honom om jag skall tillfriskna från denna sjukdom.
Så gick då Hasael honom till mötes och tog med sig skänker, allt det bästa som fanns i Damaskus, så mycket som fyrtio kameler kunde bära.
Och han kom och trädde fram för honom och sade: »Din son Ben-Hadad, konungen i Aram, har sänt mig till dig och låter fråga: 'Skall jag tillfriskna från denna sjukdom?'»
Elisa svarade honom: »Gå och säg till honom: 'Du skall tillfriskna.'
Men HERREN har uppenbarat för mig att han likväl skall dö.»
Och gudsmannen stirrade framför sig och betraktade honom länge och väl; därefter begynte han gråta.
Då sade Hasael: »Varför gråter min herre?»
Han svarade: »Därför att jag vet huru mycket ont du skall göra Israels barn: du skall sätta eld på deras fästen, deras unga män skall du dräpa med svärd, deras späda barn skall du krossa, och deras havande kvinnor skall du upprista.»
Hasael sade: »Vad är väl din tjänare, den hunden, eftersom han skulle kunna göra så stora ting?»
Elisa svarade: »HERREN har uppenbarat för mig att du skall bliva konung över Aram.»
Och han gick ifrån Elisa och kom till sin herre.
Då frågade denne honom: »Vad sade Elisa till dig?»
Han svarade: »Han sade till mig att du skall tillfriskna.»
Men dagen därefter tog han täcket och doppade det i vatten och bredde ut det över hans ansikte; detta blev hans död.
Och Hasael blev konung efter honom.
I Jorams, Ahabs sons, Israels konungs, femte regeringsår, medan Josafat var konung i Juda, blev Joram, Josafats son, konung i Juda.
Han var trettiotvå år gammal, när han blev konung, och han regerade åtta år i Jerusalem.
Men han vandrade på Israels konungars väg, såsom Ahabs hus hade gjort, ty en dotter till Ahab var hans hustru; han gjorde vad ont var i HERRENS ögon.
Dock ville HERREN icke fördärva Juda, för sin tjänare Davids skull, enligt sitt löfte till honom, att han skulle låta honom och hans söner hava en lampa för alltid.
I hans tid avföll Edom från Juda välde och satte en egen konung över sig.
Då drog Joram över till Sair med alla sina stridsvagnar.
Och om natten gjorde han ett anfall på edoméerna, som hade omringat honom, och slog dem och hövitsmannen över deras vagnar, men folket flydde till sina hyddor.
Så avföll Edom från Juda välde, och det har varit skilt därifrån ända till denna dag.
Vid just samma tid avföll ock Libna.
Vad nu mer är att säga om Joram och om allt vad han gjorde, det finnes upptecknat i Juda konungars krönika.
Och Joram gick till vila hos sina fäder och blev begraven hos sina fäder i Davids stad.
Och hans son Ahasja blev konung efter honom.
I Jorams, Ahabs sons, Israels konungs, tolfte regeringsår blev Ahasja, Jorams son, konung i Juda.
Tjugutvå år gammal var Ahasja, när han blev konung, och han regerade ett år i Jerusalem.
Hans moder hette Atalja, dotter till Omri, Israels konung.
Han vandrade på Ahabs hus' väg och gjorde vad ont var i HERRENS ögon likasom Ahabs hus; han var ju nära besläktad med Ahabs hus.
Och han drog åstad med Joram, Ahabs son, och stridde mot Hasael, konungen i Aram, vid Ramot Gilead.
Men Joram blev sårad av araméerna.
Då vände konung Joram tillbaka, för att i Jisreel låta hela sig från de sår som araméerna hade tillfogat honom vid Rama, i striden mot Hasael, konungen i Aram.
Och Ahasja, Jorams son, Juda konung, for ned för att besöka Joram, Ahabs son, i Jisreel, eftersom denne låg sjuk.
Profeten Elisa kallade till sig en av profetlärjungarna och sade till honom: »Omgjorda dina länder och tag denna oljeflaska med dig, och gå till Ramot i Gilead.
Och när du har kommit dit, så sök upp Jehu, son till Josafat, son till Nimsi, och gå in och bed honom stå upp, där han sitter bland sina bröder, och för honom in i den innersta kammaren.
Tag så oljeflaskan och gjut olja på hans huvud och säg: 'Så säger HERREN: Jag har smort dig till konung över Israel.'
Öppna sedan dörren och fly, utan att dröja.»
Så gick då den unge mannen, profetens tjänare, åstad till Ramot i Gilead.
Och när han kom dit, fick han se härens hövitsmän sitta där.
Då sade han: »Jag har ett ärende till dig, hövitsman.»
Jehu frågade: »Till vem av oss alla här?»
Han svarade: »Till dig själv, hövitsman.»
Då stod han upp och gick in i huset; och han göt oljan på hans huvud och sade till honom: »Så säger HERREN Israels Gud: Jag har smort dig till konung över HERRENS folk, över Israel.
Och du skall förgöra Ahabs, din herres, hus; ty jag vill på Isebel hämnas mina tjänare profeterna blod, ja, alla HERRENS tjänares blod.
Och Ahabs hela hus skall förgås jag skall utrota allt mankön av Ahab hus, både små och stora i Israel.
Och jag skall göra med Ahab hus såsom jag gjorde med Jerobeams, Nebats sons, hus, och såsom jag gjorde med Baesas, Ahias sons, hus.
Och hundarna skola äta upp Isebel på Jisreels åkerfält, och ingen skall begrava henne.»
Därefter öppnade han dörren och flydde.
När sedan Jehu åter kom ut till sin herres tjänare, frågade man honom: »Allt står väl rätt till?
Varför kom denne vanvetting till dig?»
Han svarade dem: »I kännen ju den mannen och hans tal.»
Men de sade: »Du vill bedraga oss; säg oss sanningen.»
Då sade han: »Så och så talade han till mig och sade: 'Så säger HERREN: Jag har smort dig till konung över Israel.'»
Strax tog då var och en av dem sin mantel och lade den under honom på själva trappan; och de stötte i basun och ropade: »Jehu har blivit konung.»
Och Jehu, son till Josafat, son till Nimsi, anstiftade nu en sammansvärjning mot Joram.
(Joram hade då med hela Israel legat vid Ramot i Gilead för att försvara det mot Hasael, konungen i Aram;
men själv hade konung Joram vänt tillbaka, för att i Jisreel låta hela sig från de sår som araméerna hade tillfogat honom under hans strid mot Hasael, konungen i Aram.)
Och Jehu sade: »Om I så viljen, så låten ingen slippa ut ur staden, som kan gå åstad och berätta detta i Jisreel.»
Och Jehu steg upp i sin vagn och for till Jisreel, ty Joram låg sjuk där; och Ahasja, Juda konung, hade farit ditned för att besöka Joram.
När nu väktaren som stod på tornet i Jisreel fick se Jehus skara, då han kom, sade han: »Jag ser en skara.»
Då bjöd Joram att man skulle taga en ryttare och sända honom dem till mötes och låta honom fråga om allt stode rätt till.
Ryttaren red honom då till mötes och sade: »Konungen låter fråga 'Allt står väl rätt till?'»
Då svarade Jehu: »Vad kommer den saken dig vid?
Vänd, och följ efter mig.»
Och väktaren berättade och sade: »Den utskickade har hunnit fram till dem, men han kommer icke tillbaka.»
Då sände han en annan ryttare. när denne hade hunnit fram till dem, sade han: »Konungen låter fråga: 'Allt står väl rätt till?'»
Jehu svarade: »Vad kommer den saken dig vid?
Vänd, och följ efter mig.»
Väktaren berättade åter och sade: »Han har hunnit fram till dem men han kommer icke tillbaka.
På deras sätt att fara fram ser det ut som vore det Jehu, Nimsis son, ty han far fram såsom en vanvetting.»
Då sade Joram: »Spänn för.»
Och man spände för hans vagn.
Och Joram, Israels konung, for nu ut med Ahasja, Juda konung, var och en i sin vagn; de foro ut för att möta Jehu.
Och de träffade tillsammans med honom på jisreeliten Nabots åkerstycke.
När Joram nu fick se Jehu, sade han: »Allt står väl rätt till, Jehu?»
Denne svarade: »Huru skulle det kunna stå rätt till, så länge som du tål din moder Isebels avgudiska väsen och hennes många trolldomskonster?»
Då svängde Joram om vagnen och flydde, i det han ropade till Ahasja: »Förräderi, Ahasja!»
Men Jehu hade fattat bågen i sin hand och sköt Joram i ryggen, att pilen gick ut genom hjärtat, och han sjönk ned i sin vagn.
Därefter sade han till sin livkämpe Bidkar: »Tag honom och kasta ut honom på jisreeliten Nabots åkerstycke; kom ihåg huru HERREN, när jag och du bredvid varandra redo bakom hans fader Ahab, om denne uttalade den utsagan:
'Sannerligen, så visst som jag i går såg Nabots och hans söners blod, säger HERREN, skall jag just på detta åkerstycke vedergälla dig, säger HERREN.'
Tag därför honom nu och kasta ut honom här på åkerstycket, i enlighet med HERRENS ord.»
När Ahasja, Juda konung, såg detta, flydde han åt Trädgårdshuset till.
Men Jehu jagade efter honom och ropade: »Skjuten ned också honom i vagnen.»
Så skedde ock på Gurhöjden vid Jibleam; men han flydde vidare till Megiddo och dog där.
Sedan förde hans tjänare honom i vagnen till Jerusalem; och man begrov honom i hans grav hos hans fäder, i Davids stad.
Ahasja hade blivit konung över Juda i Jorams, Ahabs sons, elfte regeringsår.
Så kom nu Jehu till Jisreel.
När Isebel fick höra detta, sminkade hon sig kring ögonen och smyckade sitt huvud och såg ut genom fönstret.
Och när Jehu kom in genom porten, ropade hon: »Allt står väl rätt till, du, Simri, som har dräpt din herre?»
Han lyfte sitt ansikte upp mot fönstret och sade: »Vem håller med mig?
Vem?»
Då sågo två eller tre hovmän ut, ned på honom.
Han sade: »Störten ned henne.»
Och de störtade ned henne, så att hennes blod stänkte på väggen och på hästarna; och han körde över henne.
Därefter gick han in och åt och drack.
Sedan sade han: »Tagen vara på henne, den förbannade, och begraven henne, ty hon är dock en konungadotter.»
Men när de då gingo åstad för att begrava henne, funno de av henne intet annat än huvudskålen, fötterna och händerna.
och de vände tillbaka och berättade detta för honom.
Då sade han: »Detta är vad HERREN talade genom sin tjänare tisbiten Elia, i det han sade: 'På Jisreels åkerfält skola hundarna äta upp Isebels kött;
och Isebels döda kropp skall ligga såsom gödsel på marken på Jisreels åkerfält, så att ingen skall kunna säga: Detta är Isebel.'»
Men Ahab hade sjuttio söner i Samaria.
Och Jehu skrev brev och sände till Samaria, till de överste i Jisreel, de äldste, och till de fostrare som Ahab hade utsett;
han skrev: »Nu, när detta brev kommer eder till handa, I som haven eder herres söner hos eder, och som haven vagnarna och hästarna hos eder, och därtill en befäst stad och vapen,
mån I utse den som är bäst och lämpligast av eder herres söner och sätta honom på hans faders tron och strida för eder herres hus.»
Men de blevo övermåttan förskräckta och sade: »De två konungarna hava ju icke kunnat hålla stånd mot honom; huru skulle då vi kunna hålla stånd!»
Och överhovmästaren och hövdingen över staden och de äldste och konungasönernas fostrare sände till Jehu och läto säga: »Vi äro dina tjänare; allt vad du säger oss villa vi göra.
Vi vilja icke göra någon till konung; gör vad dig täckes.»
Då skrev han ett annat brev till dem, vari det stod: »Om I hållen med mig och viljen lyssna till mina ord, så tagen huvudena av eder herres söner och kommen i morgon vid denna tid till mig i Jisreel.»
De sjuttio konungasönerna bodde nämligen hos de store i staden, vilka fostrade dem.
Då nu brevet kom dem till handa, togo de konungasönerna och slaktade dem, alla sjuttio, och lade deras huvuden i korgar och sände dem till honom i Jisreel.
När då ett bud kom och berättade för honom att de hade fört dit konungasönernas huvuden, sade han: »Läggen dem till i morgon i två högar vid ingången till porten.»
Och om morgonen gick han ut och ställde sig där och sade till allt folket: »I ären utan skuld.
Det är jag som har anstiftat sammansvärjningen mot min herre och dräpt honom; men vem har slagit ihjäl alla dessa?
Märken nu huru intet av HERRENS ord faller till jorden, intet som HERREN har talat mot Ahabs hus.
Ja, HERREN har gjort vad han har sagt genom sin tjänare Elia.»
Sedan, dräpte Jehu alla som voro kvar av Ahabs hus i Jisreel, så ock alla hans store och hans förtrogne och hans präster; han lät ingen slippa undan.
Därefter stod han upp och begav sig åstad till Samaria; men under vägen, när Jehu kom till Bet-Eked-Haroim,
träffade han på Ahasjas, Juda konungs, bröder.
Han frågade dem: »Vilka ären I?»
De svarade: »Vi äro Ahasjas bröder, och vi äro på väg ned för att hälsa på konungasönerna och konungamoderns söner.»
Han sade: »Gripen dem levande.»
Då grepo de dem levande och slaktade dem och kastade dem i Bet-Ekeds brunn, alla fyrtiotvå; han lät ingen av dem bliva kvar.
När han sedan begav sig därifrån, träffade han Jonadab, Rekabs son, som kom honom till mötes; och han hälsade på honom och sade till honom: »Är du lika redligt sinnad mot mig som jag är mot dig?»
Jonadab svarade: »Ja.» »Är det så», sade han, »så räck mig din hand.»
Då räckte han honom sin hand; och han lät honom stiga upp till sig i vagnen.
Och han sade: »Far med mig och se huru jag nitälskar för HERREN.»
Så körde man åstad med honom i hans vagn.
Och när han kom till Samaria, dräpte han alla som voro kvar av Ahabs hus i Samaria och förgjorde det så, i enlighet med det ord som HERREN hade talat till Elia.
Och Jehu församlade allt folket och sade till dem: »Ahab har tjänat Baal litet; Jehu skall tjäna honom mycket.
Så kallen nu hit till mig alla Baals profeter, alla hans tjänare och alla hans präster -- ingen får saknas -- ty jag har ett stort offer åt Baal i sinnet; var och en som saknas skall mista livet.»
Men Jehu gjorde så med led list, i avsikt att utrota Baals tjänare.
Därefter sade Jehu: »Pålysen en helig högtidsförsamling åt Baal.»
Då lyste man ut en sådan.
Och Jehu sände bud över hela Israel, och alla Baals tjänare kommo; Ingen underlät att komma.
Och de gingo in i Baals tempel, och Baals tempel blev fullt, ifrån den ena ändan till den andra.
Sedan sade han till föreståndaren för klädkammaren: »Tag fram kläder åt alla Baals tjänare.»
Och han tog fram kläderna åt dem.
Därefter gick Jehu in i Baals tempel med Jonadab, Rekabs son.
Och han sade till Baals tjänare: »Sen nu noga efter, att här bland eder icke finnes någon HERRENS tjänare, utan allenast sådana som tjäna Baal.
De gingo alltså in för att offra slaktoffer och brännoffer.
Men Jehu hade därutanför ställt åttio man och sagt: »Om någon slipper undan av de män som jag nu överlämnar i edra händer, så skall liv givas för liv.»
Och när man hade offrat brännoffret, sade Jehu till drabanterna och kämparna: »Gån in och slån ned dem; låten ingen komma ut.»
Och de slogo dem med svärdsegg, och drabanterna och kämparna kastade undan deras kroppar.
Därefter gingo de in i det inre av Baals tempel
och kastade ut stoderna ur Baals tempel och brände upp dem.
Och själva Baalsstoden bröto de ned; de bröto ock ned Baals tempel och gjorde därav avträden, som finnas kvar ännu i dag.
Så utrotade Jehu Baal ur Israel.
Men från de Jerobeams, Nebats sons, synder genom vilka denne hade kommit Israel att synda, från dem avstod icke Jehu, icke från guldkalvarna i Betel och Dan.
Och HERREN sade till Jehu: »Därför att du har väl utfört vad rätt var i mina ögon, och gjort mot Ahabs hus allt vad jag hade i sinnet, därför skola dina söner till fjärde led sitta på Israels tron.
Men Jehu tog dock icke i akt att vandra efter HERRENS, Israels Guds, lag av allt sitt hjärta; han avstod icke från de Jerobeams synder genom vilka denne hade kommit Israel att synda.
Vid denna tid begynte HERREN skära bort stycken från Israel, ty Hasael slog israeliterna utefter hela deras gräns
och intog östra sidan om Jordan hela landet Gilead, gaditernas, rubeniternas och manassiternas land, området från Aroer vid bäcken Arnon, både Gilead och Basan.
Vad nu mer är att säga om Jehu, om allt vad han gjorde och om alla hans bedrifter, det finnes upptecknat i Israels konungars krönika.
Och Jehu gick till vila hos sina fäder, och man begrov honom i Samaria.
Och hans son Joahas blev konung efter honom.
Den tid Jehu regerade över Israel Samaria var tjuguåtta år.
När Atalja, Ahasjas moder, förnam att hennes son var död, stod hon upp och förgjorde hela konungasläkten.
Men just när konungabarnen skulle dödas, tog Joseba, konung Jorams dotter, Ahasjas syster, Joas, Ahasjas son, och skaffade honom jämte hans amma hemligen undan, in i sovkammaren; där höll man honom dold för Atalja, så att han icke blev dödad.
Sedan var han hos henne i HERRENS hus, där han förblev gömd i sex år, medan Atalja regerade i landet.
Men i det sjunde året sände Jojada åstad och lät hämta karéernas och drabanternas underhövitsmän och förde dem in till sig i HERRENS hus; och sedan han hade gjort en överenskommelse med dem och tagit en ed av dem i HERRENS hus visade han dem konungens son.
Därefter bjöd han dem och sade: »Detta är vad I skolen göra: en tredjedel av eder, I som haven att inträda i vakthållningen på sabbaten, skall hålla vakt i konungshuset
och en tredjedel vid Surporten och en tredjedel vid porten bakom drabanterna; så skolen hålla vakt vid huset var i sin ordning.
Men de båda andra avdelningarna av eder, nämligen alla som hava att avgå från vakthållningen på sabbaten, de skola hålla vakt i HERRENS hus hos konungen.
I skolen ställa eder runt omkring; konungen, var och en med sina vapen i handen; och om någon vill tränga sig inom leden, skall han dödas.
Och I skolen följa konungen, vare sig han går ut eller in.
Underhövitsmännen gjorde allt vad prästen Jojada hade bjudit dem; var och en av dem tog sina män, både de som skulle inträda i vakthållningen på sabbaten och de som skulle avgå därifrån på sabbaten, och de kommo så till prästen Jojada.
Och prästen gav åt underhövitsmännen det spjut och de sköldar som hade tillhört konung David, och som funnos i HERRENS hus.
Och drabanterna ställde upp sig, var och en med sina vapen i handen, från husets södra sida till husets norra sida, mot altaret och mot huset, runt omkring konungen.
Därefter förde han ut konungasonen och satte på honom kronan och gav honom vittnesbördet; och de gjorde honom till konung och smorde honom.
Och de klappade i händerna och ropade: »Leve konungen!»
När Atalja nu hörde drabanternas och folkets rop, gick hon in i HERRENS hus till folket.
Där fick hon då se konungen stå vid pelaren, såsom övligt var, och hövitsmännen och trumpetblåsarna bredvid konungen, och fick höra huru hela folkmängden jublade och stötte i trumpeterna.
Då rev Atalja sönder sina kläder och utropade: »Sammansvärjning!
Sammansvärjning!»
Men prästen Jojada gav underhövitsmännen som anförde skaran denna befallning: »Fören henne ut mellan leden, och om någon följer henne, så må han dödas med svärd.»
Prästen ville nämligen förhindra att hon dödades i HERRENS hus.
Alltså grepo de henne, och när hon hade kommit till den plats där hästarna plägade föras in i konungshuset, dödades hon där.
Och Jojada slöt det förbundet mellan HERREN, konungen och folket, att de skulle vara ett HERRENS folk; han slöt ock ett förbund mellan konungen och folket.
Och hela folkmängden begav sig till Baals tempel och rev ned det och förstörde i grund dess altaren och dess bilder; och Mattan, Baals präst, dräpte de framför altarna.
Därefter ställde prästen ut vakter vid HERRENS hus.
Och han tog med sig underhövitsmännen jämte karéerna och drabanterna och hela folkmängden, och de förde konungen ned från HERRENS hus och gingo in i konungshuset genom Drabantporten; och han satte sig på konungatronen.
Och hela folkmängden gladde sig, och staden förblev lugn.
Men Atalja hade de dödat med svärd i konungshuset.
Joas var sju år gammal, när han blev konung.
I Jehus sjunde regeringsår blev Joas konung, och han regerade fyrtio år i Jerusalem.
Hans moder hette Sibja, från Beer-Seba.
Och Joas gjorde vad rätt var HERRENS ögon, så länge han levde, prästen Jojada hade varit hans lärare.
Dock blevo offerhöjderna icke avskaffade, utan folket fortfor att frambära offer och tända offereld på höjderna.
Och Joas sade till prästerna: »Alla penningar vilka såsom heliga gåvor inflyta till HERRENS hus, gångbara penningar, sådana som utgöra lösen för personer, efter det värde som för var och en bestämmes, och alla penningar som någon av sitt hjärta manas att bära till HERRENS hus,
dem skola prästerna taga emot, var och en av sina bekanta, och de skola därmed sätta i stånd vad som är förfallet på HERRENS hus, överallt där något förfallet finnes.»
Men i konung Joas' tjugutredje regeringsår hade prästerna ännu icke satt i stånd vad som var förfallet på huset.
Då kallade konung Joas till sig prästen Jojada och de övriga prästerna och sade till dem: »Varför sätten I icke i stånd vad som är förfallet på huset?
Nu fån I icke längre taga emot penningar av edra bekanta, utan I skolen lämna dem ifrån eder till det som är förfallet på huset.»
Och prästerna samtyckte till att icke taga emot penningar av folket, och ej heller befatta sig med att sätta i stånd vad som var förfallet på huset.
Då tog prästen Jojada en kista och borrade ett hål på locket och ställde den bredvid altaret, på högra sidan, när man går in i HERRENS hus.
Och prästerna som höllo vakt vid tröskeln lade dit alla penningar som inflöto till HERRENS hus.
Men så snart de då märkte att mycket penningar fanns i kistan, gick konungens sekreterare ditupp jämte översteprästen, och de knöto in och räknade sedan de penningar som funnos i HERRENS hus.
Därefter överlämnades de uppvägda penningarna åt de män som förrättade arbete såsom tillsyningsmän vid HERRENS hus, och dessa betalade ut dem åt de timmermän och byggningsmän som arbetade på HERRENS hus,
och åt murarna och stenhuggarna, så ock till inköp av trävirke och huggen sten för att sätta i stånd vad som var förfallet på HERRENS hus, korteligen, till alla utgifter för att sätta huset i stånd.
Men man gjorde inga silverfat för HERRENS hus, ej heller knivar, skålar, trumpeter eller andra föremål av guld eller av silver, för de penningar som inflöto till HERRENS hus,
utan man gav dem åt arbetarna, och dessa satte därför HERRENS hus i stånd.
Och man höll icke någon räkenskap med de män åt vilka penningarna överlämnades, för att de skulle giva dem åt arbetarna, utan de fingo handla på heder och tro.
Men skuldoffers- och syndofferspenningarna gingo icke till HERRENS hus utan tillföllo prästerna.
På den tiden drog Hasael, konungen i Aram, upp och belägrade Gat och intog det, därefter ställde Hasael sitt tåg upp mot Jerusalem.
Då tog Joas, Juda konung, allt vad hans fäder Josafat, Joram och Ahasja, Juda konungar, hade helgat åt HERREN, och vad han själv hade helgat åt HERREN, och allt guld som fanns i skattkamrarna i HERRENS hus och i konungshuset, och sände det till Hasael, konungen i Aram, och då lämnade denne Jerusalem i fred.
Vad nu mer är att säga om Joas och om allt vad han gjorde, det finnes upptecknat i Juda konungars krönika.
Och hans tjänare uppreste sig och sammansvuro sig och dräpte Joas i Millobyggnaden, som sträcker sig ned mot Silla.
Det var hans tjänare Josakar, Simeats son, och Josabad, Somers son, som slogo honom till döds.
Och man begrov honom hos hans fäder i Davids stad.
Och hans son Amasja blev konung efter honom
I Joas', Ahasjas sons, Juda konungs, tjugutredje regeringsår blev Joahas, Jehus son, konung över Israel i Samaria och regerade i sjutton år.
Han gjorde vad ont var i HERRENS ögon och följde efter de Jerobeams, Nebats sons, synder genom vilka denne hade kommit Israel att synda; från dem avstod han icke.
Då upptändes HERRENS vrede mot Israel, och han gav dem i Hasaels, den arameiske konungens, hand och i Ben-Hadads, Hasaels sons, hand hela denna tid.
(Men Joahas bönföll inför HERREN, och HERREN hörde honom, eftersom han såg Israels betryck, då nu konungen i Aram förtryckte dem.
Och HERREN gav åt Israel en frälsare, så att de blevo räddade ur araméernas hand; sedan bodde Israels barn i sina hyddor såsom förut.
Dock avstodo de icke från de Jerobeams hus' synder genom vilka denne hade kommit Israel att synda, utan vandrade i dem.
Aseran fick också stå kvar i Samaria.)
Ty han hade icke låtit Joahas behålla mer folk än femtio ryttare, tio vagnar och tio tusen man fotfolk; så illa förgjorde dem konungen i Aram; han slog dem, så att de blevo såsom stoft, när man tröskar.
Vad nu mer är att säga om Joahas, om allt vad han gjorde och om hans bedrifter, det finnes upptecknat i Israels konungars krönika.
Och Joahas gick till vila hos sina fäder, och man begrov honom i Samaria.
Och hans son Joas blev konung efter honom.
I Joas', Juda konungs, trettiosjunde regeringsår blev Joas, Joahas' son, konung över Israel i Samaria och regerade i sexton år.
Han gjorde vad ont var i HERRENS ögon; han avstod icke från någon av de Jerobeams, Nebats sons, synder genom vilka denne hade kommit Israel att synda, utan vandrade i dem.
Vad nu mer är att säga om Joas, om allt vad han gjorde och om hans bedrifter, om hans krig mot Amasja, Juda konung, det finnes upptecknat i Israels konungars krönika.
Och Joas gick till vila hos sina fäder, och Jerobeam besteg hans tron.
Och Joas blev begraven i Samaria, hos Israels konungar.
Men när Elisa låg sjuk i den sjukdom varav han dog, kom Joas, Israels konung, ned till honom.
Och han satt hos honom gråtande och sade: »Min fader, min fader!
Du som för Israel är både vagnar och ryttare!»
Då sade Elisa till honom: »Hämta en båge och pilar.»
Och han hämtade åt honom en båge och pilar.
Då sade han till Israels konung: »Fatta i bågen med din hand.»
Och när han hade gjort detta, lade Elisa sina händer på konungens händer.
Därefter sade han: »Öppna fönstret mot öster.»
Och när han hade öppnat det, sade Elisa: »Skjut.»
Och han sköt.
Då sade han: »En HERRENS segerpil, en segerpil mot Aram!
Du skall slå araméerna vid Afek, så att de förgöras.»
Därefter sade han: »Tag pilarna.»
Och när han hade tagit dem, sade han till Israels konung: »Slå på jorden.»
Då slog han tre gånger och sedan höll han upp.
Då blev gudsmannen vred på honom och sade: »Du skulle slagit fem eller sex gånger, ty då skulle du hava slagit araméerna så, att de hade blivit förgjorda; men nu kommer du att slå araméerna allenast tre gånger.»
Så dog då Elisa, och man begrov honom.
Men moabitiska strövskaror plägade falla in i landet, vid årets ingång.
Så hände sig, att just när några höllo på att begrava en man, fingo de se en strövskara; då kastade de mannen i Elisas grav.
När då mannen kom i beröring med Elisas ben, fick han liv igen och reste sig upp på sina fötter.
Och Hasael, konungen i Aram, hade förtryckt Israel, så länge Joahas levde.
Men HERREN blev dem nådig och förbarmade sig över dem och vände sig till dem, för det förbunds skull som han hade slutit med Abraham, Isak och Jakob; ty han ville icke fördärva dem, och han hade ännu icke kastat dem bort ifrån sitt ansikte.
Och Hasael, konungen i Aram, dog, och hans son Ben-Hadad blev konung efter honom.
Då tog Joas, Joahas' son, tillbaka från Ben-Hadad, Hasaels son, de städer som denne i krig hade tagit ifrån hans fader Joahas.
Tre gånger slog Joas honom och återtog så Israels städer.
I Joas', Joahas' sons, Israels konungs, andra regeringsår blev Amasja, Joas' son, konung i Juda.
Han var tjugufem år gammal, när han blev konung, och han regerade tjugunio år i Jerusalem.
Hans moder hette Joaddin, från Jerusalem.
Han gjorde vad rätt var i HERRENS ögon, dock icke såsom hans fader David; men han gjorde i allt såsom hans fader Joas hade gjort.
Offerhöjderna blevo likväl icke avskaffade, utan folket fortfor att frambära offer och tända offereld på höjderna.
Och sedan konungadömet hade blivit befäst i hans hand, lät han dräpa dem av sina tjänare, som hade dräpt hans fader, konungen.
Men mördarnas barn dödade han icke, i enlighet med vad föreskrivet var i Moses lagbok, där HERREN hade bjudit och sagt: »Föräldrarna skola icke dödas för sina barns skull, och barnen skola icke dödas för sina föräldrars skull, utan var och en skall dö genom sin egen synd.»
Han slog edoméerna i Saltdalen, tio tusen man, och intog Sela med strid och gav det namnet Jokteel, såsom det heter ännu i dag.
Därefter skickade Amasja sändebud till Joas, son till Joahas, son till Jehu, Israels konung, och lät säga: »Kom, låt oss drabba samman med varandra.»
Men Joas, Israels konung, sände då till Amasja, Juda konung, och lät svara: »Törnbusken på Libanon sände en gång bud till cedern på Libanon och lät säga: 'Giv din dotter åt min son till hustru.'
Men sedan gingo markens djur på Libanon fram över törnbusken och trampade ned den.
Du har slagit Edom, och däröver förhäver du dig i ditt hjärta.
Men låt dig nöja med den äran, och stanna hemma.
Varför utmanar du olyckan, dig själv och Juda med dig till fall?»
Men Amasja ville icke höra härpå, och Joas, Israels konung, drog då upp, och de drabbade samman med varandra, han och Amasja, Juda konung, vid det Bet-Semes som hör till Juda.
Och Juda män blevo slagna av Israels män och flydde, var och en till sin hydda.
Och Amasja, Juda konung, son till Joas, son till Ahasja, blev tagen till fånga i Bet-Semes av Joas, Israels konung.
Och när de kommo till Jerusalem, bröt han ned ett stycke av Jerusalems mur vid Efraimsporten, och därifrån ända till Hörnporten, fyra hundra alnar.
Och han tog allt guld och silver och alla kärl som funnos i HERRENS hus och i konungshusets skattkamrar, därtill ock gisslan, och vände så tillbaka till Samaria.
Vad nu mer är att säga om Joas, om vad han gjorde och om hans bedrifter och om hans krig mot Amasja, Juda konung, det finnes upptecknat i Israels konungars krönika.
Och Joas gick till vila hos sina fäder och blev begraven i Samaria, hos Israels konungar.
Och hans son Jerobeam blev konung efter honom.
Men Amasja, Joas' son, Juda konung, levde i femton år efter Joas', Joahas' sons, Israels konungs, död.
Vad nu mer är att säga om Amasja, det finnes upptecknat i Juda konungars krönika.
Och en sammansvärjning anstiftades mot honom i Jerusalem, så att han måste fly till Lakis.
Då sändes män efter honom till Lakis, och dessa dödade honom där.
Sedan förde man honom därifrån på hästar; och han blev begraven i Jerusalem hos sina fäder i Davids stad.
Och allt folket i Juda tog Asarja som då var sexton år gammal, och gjorde honom till konung i hans fader Amasjas ställe.
Det var han som befäste Elat; ock han lade det åter under Juda, sedan konungen hade gått till vila hos sina fäder.
I Amasjas, Joas' sons, Juda konungs, femtonde regeringsår blev Jerobeam, Joas' son, konung över Israel i Samaria och regerade i fyrtioett år.
Han gjorde vad ont var i HERRENS ögon; han avstod icke från någon av de Jerobeams, Nebats sons, synder genom vilka denne hade kommit Israel att synda.
Han återvann Israels område, från det ställe där vägen går till Hamat ända till Hedmarkshavet, i enlighet med det ord som HERREN, Israels Gud, hade talat genom sin tjänare profeten Jona, Amittais son, från Gat-Hahefer.
Ty HERREN såg att Israels betryck var mycket svårt, och att det var ute med alla och envar, och att Israel icke hade någon hjälpare.
Och HERREN hade ännu icke beslutit att utplåna Israels namn under himmelen; därför frälste han dem genom Jerobeam, Joas' son.
Vad nu mer är att säga om Jerobeam, om allt vad han gjorde och om hans bedrifter och hans krig, så ock om huru han åt Israel återvann den del av Damaskus och Hamat, som en gång hade tillhört Juda, det finnes upptecknat i Israels konungars krönika.
Och Jerobeam gick till vila hos sina fäder, Israels konungar.
Och hans son Sakarja blev konung efter honom.
I Jerobeams, Israels konungs, tjugusjunde regeringsår blev Asarja, Amasjas son, konung i Juda.
Han var sexton år gammal, när han blev konung, och han regerade femtiotvå år i Jerusalem.
Hans moder hette Jekolja, från Jerusalem.
Han gjorde vad rätt var i HERRENS ögon, alldeles såsom hans fader Amasja hade gjort.
Dock blevo offerhöjderna icke avskaffade, utan folket fortfor att frambära offer och tända offereld på höjderna.
Men HERREN hemsökte konungen, så att han blev spetälsk för hela sitt liv; och han bodde sedan i ett särskilt hus.
Jotam, konungens son, förestod då hans hus och dömde folket i landet.
Vad nu mer är att säga om Asarja och om allt vad han gjorde, det finnes upptecknat i Juda konungars krönika.
Och Asarja gick till vila hos sina fäder, och man begrov honom hos hans fäder i Davids stad.
Och hans son Jotam blev konung efter honom.
I Asarjas, Juda konungs, trettioåttonde regeringsår blev Sakarja, Jerobeams son, konung över Israel i Samaria och regerade i sex månader.
Han gjorde vad ont var i HERRENS ögon, såsom hans fäder hade gjort; han avstod icke från de Jerobeams, Nebats sons, synder genom vilka denne hade kommit Israel att synda.
Och Sallum, Jabes' son, anstiftade en sammansvärjning mot honom och slog honom till döds i folkets åsyn, och blev så konung i hans ställe
Vad nu mer är att säga om Sakarja, det finnes upptecknat i Israels konungars krönika.
Så, uppfylldes det ord som HERREN, hade talat till Jehu, när han sade: »Dina söner till fjärde led skola sitta på Israels tron.»
Det skedde så.
Sallum, Jabes' son, blev konung i Ussias, Juda konungs, trettionionde regeringsår, och han regerade en månads tid i Samaria.
Men då drog Menahem, Gadis son, upp från Tirsa och kom till Samaria och slog Sallum, Jabes' son, till döds i Samaria, och blev så konung i hans ställe
Vad nu mer är att säga om Sallum och om den sammansvärjning han anstiftade, det finnes upptecknat i Israels konungars krönika.
Vid den tiden förhärjade Menahem Tifsa med allt vad därinne var, så ock hela dess område, från Tirsa; ty staden hade icke öppnat portarna, därför härjade han den, och alla dess havande kvinnor lät han upprista.
I Asarjas, Juda konungs, trettionionde regeringsår blev Menahem, Gadis son, konung över Israel och regerade i tio år, i Samaria.
Han gjorde vad ont var i HERRENS ögon; han avstod icke, så länge han levde, från de Jerobeams Nebats sons, synder genom vilka denne hade kommit Israel att synda.
Och Pul, konungen i Assyrien, föll in i landet; då gav Menahem åt Pul tusen talenter silver, för att han skulle understödja honom och befästa konungadömet i hans hand.
Och de penningar som Menahem skulle giva åt konungen i Assyrien tog han ut genom att lägga skatt på alla rika män i Israel, en skatt av femtio siklar silver på var och en.
Så vände då konungen i Assyrien tillbaka och stannade icke där i landet.
Vad nu mer är att säga om Menahem och om allt vad han gjorde, det finnes upptecknat i Israels konungars krönika.
Och Menahem gick till vila hos sina fäder.
Och hans son Pekaja blev konung efter honom.
I Asarjas, Juda konungs, femtionde regeringsår blev Pekaja, Menahems son, konung över Israel i Samaria och regerade i två år.
Han gjorde vad ont var i HERRENS ögon; han avstod icke från de Jerobeams, Nebats sons, synder genom vilka denne hade kommit Israel att synda.
Och Peka, Remaljas son, hans livkämpe, anstiftade en sammansvärjning mot honom och dräpte honom i Samaria, i konungshusets palatsbyggnad, han tillika med Argob och Arje; därvid hade han med sig femtio gileaditer.
Så dödade han honom och blev konung i hans ställe.
Vad nu mer är att säga om Pekaja och om allt vad han gjorde, det finnes upptecknat i Israels konungars krönika.
I Asarjas, Juda konungs, femtioandra regeringsår blev Peka, Remaljas son, konung över Israel i Samaria och regerade i tjugu år.
Han gjorde vad ont var i HERRENS Ögon; han avstod icke från de Jerobeams; Nebats sons, synder genom vilka denne hade kommit Israel att synda.
I Pekas, Israels konungs, tid kom Tiglat-Pileser, konungen i Assyrien, och intog Ijon, Abel-Bet-Maaka, Janoa, Kedes, Hasor, Gilead och Galileen, hela Naftali land, och förde folket bort till Assyrien.
Och Hosea, Elas son, anstiftade en sammansvärjning mot Peka, Remaljas son, och slog honom till döds och blev så konung i hans ställe, i Jotams, Ussias sons, tjugonde regeringsår.
Vad nu mer är att säga om Peka och om allt vad han gjorde, det finnes upptecknat i Israels konungars krönika.
I Pekas, Remaljas sons, Israels konungs, andra regeringsår blev Jotam, Ussias son, konung i Juda.
Han var tjugufem år gammal, när han blev konung, och han regerade sexton år i Jerusalem.
Hans moder hette Jerusa, Sadoks dotter.
Han gjorde vad rätt var i HERRENS ögon; han gjorde alldeles såsom hans fader Ussia hade gjort.
Dock blevo offerhöjderna icke avskaffade, utan folket fortfor att frambära offer och tända offereld på höjderna.
Han byggde Övre porten till HERRENS hus.
Vad nu mer är att säga om Jotam, om vad han gjorde, det finnes upptecknat i Juda konungars krönika.
Vid den tiden begynte HERREN att låta Juda hemsökas av Resin, konungen i Aram, och av Peka, Remaljas son.
Och Jotam gick till vila hos sina fäder och blev begraven hos sina fäder i sin fader Davids stad.
Och hans son Ahas blev konung efter honom.
I Pekas, Remaljas sons, sjuttonde regeringsår blev Ahas, Jotams son, konung i Juda.
Tjugu år gammal var Ahas, när han blev konung, och han regerade sexton år i Jerusalem.
Han gjorde icke vad rätt var i HERRENS, sin Guds, ögon, såsom hans fader David,
utan vandrade på Israels konungars väg; ja, han lät ock sin son gå genom eld, efter den styggeliga seden hos de folk som HERREN hade fördrivit för Israels barn.
Och han frambar offer och tände offereld på höjderna och kullarna och under alla gröna träd.
På den tiden drogo Resin, konungen i Aram, och Peka, Remaljas son, Israels konung, upp för att erövra Jerusalem; och de inneslöto Ahas, men kunde icke erövra staden.
Vid samma tid återvann Resin, konungen i Aram, Elat åt Aram och jagade Juda män bort ifrån Elot.
Därefter kommo araméerna till Elat och bosatte sig där, och där bo de ännu i dag.
Men Ahas skickade sändebud till Tiglat-Pileser, konungen i Assyrien, och lät säga: »Jag är din tjänare och din son.
Drag hitupp och fräls mig från Arams konung och från Israels konung, ty de hava överfallit mig.»
Och Ahas tog det silver och guld som fanns i HERRENS hus och i konungshusets skattkamrar, och sände det såsom skänk till konungen i Assyrien.
Och konungen i Assyrien lyssnade till honom: konungen i Assyrien drog upp mot Damaskus och intog det och förde bort folket till Kir och dödade Resin.
Sedan for konung Ahas till Damaskus för att där möta Tiglat-Pileser, konungen i Assyrien.
Och när konung Ahas fick se altaret i Damaskus, sände han till prästen Uria en avteckning av altaret och en mönsterbild till ett sådant, alldeles såsom det var gjort.
Sedan byggde prästen Uria altaret; alldeles efter den föreskrift som konung Ahas hade sänt till honom från Damaskus gjorde prästen Uria det färdigt, till dess konung Ahas kom tillbaka från Damaskus.
När så konungen efter sin hemkomst från Damaskus fick se altaret, trädde han fram till altaret och steg upp till det.
Därefter förbrände han sitt brännoffer och sitt spisoffer och utgöt sitt drickoffer; och blodet av det tackoffer som han offrade stänkte han på altaret.
Men kopparaltaret, som stod inför HERRENS ansikte, flyttade han undan från husets framsida, från platsen mellan det nya altaret och HERRENS hus, och ställde det på norra sidan om detta altare.
Och konung Ahas bjöd prästen Uria och sade: »På det stora altaret skall du förbränna morgonens brännoffer och aftonens spisoffer, ävensom konungens brännoffer jämte hans spisoffer, så ock brännoffer, spisoffer och drickoffer för allt folket i landet; och allt blodet, såväl av brännoffer som av slaktoffer, skall du stänka därpå.
Men vad Jag skall göra med kopparaltaret, det vill jag närmare betänka.»
Och prästen Uria gjorde alldeles såsom konung Ahas bjöd honom.
Konung Ahas lösbröt ock sidolisterna på bäckenställen och tog bort bäckenet från dem; och havet lyfte han ned från kopparoxarna som stodo därunder och ställde det på ett stengolv.
Och den täckta sabbatsgången som man hade byggt vid huset, så ock konungens yttre ingångsväg, förlade han inom HERRENS hus, för den assyriske konungens skull.
Vad nu mer är att säga om Ahas, om vad han gjorde, det finnes upptecknat i Juda konungars krönika.
Och Ahab gick till vila hos sina fäder och blev begraven hos sina fäder i Davids stad.
Och hans son Hiskia blev konung efter honom.
I Ahas', Juda konungs, tolfte regeringsår blev Hosea, Elas son, konung i Samaria över Israel och regerade i nio år.
Han gjorde vad ont var i HERRENS; ögon, dock icke såsom de israelitiska konungar som hade varit före honom
Mot honom drog den assyriske konungen Salmaneser upp; och Hosea måste bliva honom underdånig och giva honom skänker.
Men sedan märkte konungen i Assyrien att Hosea förehade stämplingar, i det att han skickade sändebud till So, konungen i Egypten och icke, såsom förut, vart år sände skänker till konungen i Assyrien Då lät konungen i Assyrien spärra in honom och hålla honom bunden i fängelse.
Ty konungen i Assyrien drog upp och angrep hela landet, och drog upp mot Samaria och belägrade det i tre år.
I Hoseas nionde regeringsår intog konungen i Assyrien Samaria och förde Israel bort till Assyrien och lät dem bo i Hala och vid Habor -- en ström i Gosan -- och i Mediens städer.
Israels barn hade ju syndat mot HERREN, sin Gud, honom som hade fört dem upp ur Egyptens land, undan Faraos, den egyptiske konungens, hand, och de hade fruktat andra gudar.
De hade ock vandrat efter de folks stadgar, som HERREN hade fördrivit för Israels barn, och efter de stadgar som Israels konungar hade uppgjort.
Ja, Israels barn hade bedrivit otillbörliga ting mot HERREN, sin Gud; de hade byggt sig offerhöjder på alla sina boningsorter, vid väktartornen såväl som i de befästa städerna.
De hade rest stoder och Aseror åt sig på alla höga kullar och under alla gröna träd.
Där hade de på alla offerhöjder tänt offereld, likasom de folk som HERREN hade drivit bort för dem, och hade gjort onda ting, så att de förtörnade HERREN.
De hade tjänat de eländiga avgudarna, fastän HERREN hade sagt till dem: »I skolen icke göra så.
Och HERREN hade varnat både Israel och Juda genom alla sina profeter och siare och sagt: »Vänden om från edra onda vägar och hållen mina bud och stadgar -- efter hela den lag som jag gav edra fäder -- så ock vad jag har låtit säga eder genom mina tjänare profeterna.»
Men de ville icke höra, utan voro hårdnackade såsom deras fäder, vilka icke trodde på HERREN, sin Gud.
De förkastade hans stadgar och det förbund som han hade slutit med deras fäder, och de förordningar som han hade givit dem, och följde efter fåfängliga avgudar och bedrevo fåfänglighet, likasom de folk som voro omkring dem, fastän HERREN hade förbjudit dem att göra såsom dessa.
De övergåvo HERRENS, sin Guds, alla bud och gjorde sig gjutna beläten, två kalvar; de gjorde sig ock Aseror och tillbådo himmelens hela härskara och tjänade Baal.
Och de läto sina söner och döttrar gå genom eld och befattade sig med spådom och övade trolldom de sålde sig till att göra vad ont var i HERRENS ögon och förtörnade honom därmed.
Därför blev ock HERREN mycket vred på Israel och försköt dem från sitt ansikte, så att icke något annat blev kvar än Juda stam allena.
Dock höll icke heller Juda HERRENS, sin Guds, bud, utan vandrade efter de stadgar som Israel hade uppgjort.
Så förkastade då HERREN all Israels säd och tuktade dem och gav dem i plundrares hand, till dess att han kastade dem bort ifrån sitt ansikte.
Ty när han hade ryckt Israel från Davids hus och de hade gjort Jerobeam, Nebats son, till konung, förförde Jerobeam Israel till att avfalla från HERREN och kom dem att begå en stor synd.
Och Israels barn vandrade i alla de synder son Jerobeam hade gjort; de avstodo icke från dem.
Men till slut försköt HERREN Israel från sitt ansikte, såsom har hade hotat genom alla sina tjänare profeterna.
Så blev Israel; bortfört från sitt land till Assyrien, där de äro ännu i dag.
Och konungen i Assyrien lät folk komma från Babel, Kuta, Ava, Hamat och Sefarvaim och bosätta sig i Samariens städer, i Israels barns ställe.
Så togo då dessa Samarien i besittning och bosatte sig i dess städer.
Men då de under den första tiden av sin vistelse där icke fruktade HERREN, sände HERREN bland dem lejon, som anställde förödelse bland dem.
Och man omtalade detta för konungen i Assyrien och sade: »De folk som du har fört bort och låtit bosätta sig i Samariens städer veta icke huru landets Gud skall dyrkas därför har han sänt lejon ibland dem, och dessa döda dem nu, eftersom de icke veta huru landets Gud skall dyrkas.»
Då bjöd konungen i Assyrien och sade: »Låten en av de präster som I haven fört bort därifrån fara dit; må de fara dit och bosätta sig där.
Och må han lära dem huru landets Gud skall dyrkas.»
Så kom då en av de präster som: de hade fört bort ifrån Samarien och bosatte sig i Betel; och han lärde dem huru de skulle frukta HERREN.
Väl gjorde sig vart folk sin egen gud och ställde upp denne i de offerhöjdshus som samariterna hade uppbyggt, vart folk för sig, i de städer där det bodde.
Folket ifrån Babel gjorde sig en Suckot-Benot, folket ifrån Kut gjorde sig en Nergal, och folket ifrån Hamat gjorde sig en Asima;
aviterna gjorde sig en Nibhas och en Tartak, och sefarviterna brände upp sina barn i eld åt Adrammelek och Anammelek, Sefarvaims gudar.
Men de fruktade också HERREN.
Och de gjorde män ur sin egen krets till offerhöjdspräster åt sig, och dessa offrade åt dem i offerhöjdshusen.
Så fruktade de visserligen HERREN, men de tjänade därjämte sina egna gudar, på samma sätt som de folk ifrån vilka man hade fört bort dem.
Ännu i dag göra de likasom förut: de frukta icke HERREN och göra icke efter de stadgar och den rätt som de hava fått, icke efter den lag och de bud som HERREN har givit Jakobs barn, den mans åt vilken han gav namnet Israel.
Ty HERREN slöt ett förbund med dem och bjöd dem och sade: »I skolen icke frukta andra gudar, ej heller tillbedja dem eller tjäna dem eller offra åt dem.
Nej, HERREN allena, som förde eder upp ur Egyptens land med stor makt och uträckt arm, honom skolen I frukta, honom skolen I tillbedja och åt honom skolen I offra.
Och de stadgar och rätter, den lag och de bud som han har föreskrivit eder, dem skolen I hålla och göra i all tid; men I skolen icke frukta andra gudar.
Det förbund som jag har slutit med eder skolen I icke förgäta; I skolen icke frukta andra gudar.
Allenast HERREN, eder Gud, skolen I frukta, så skall han rädda eder ur alla edra fienders hand.»
Men de ville icke höra härpå, utan gjorde likasom förut.
Så fruktade då dessa folk HERREN, men tjänade därjämte sina beläten.
Också deras barn och deras barnbarn göra ännu i dag såsom deras fäder gjorde.
I Hoseas, Elas sons, Israels konungs, tredje regeringsår blev Hiskia, Ahas' son, konung i Juda.
Han var tjugufem år gammal, när han blev konung, och han regerade tjugunio år i Jerusalem.
Hans moder hette Abi, Sakarjas dotter.
Han gjorde vad rätt var i HERRENS ögon, alldeles såsom hans fader David hade gjort.
Han avskaffade offerhöjderna, slog sönder stoderna och högg ned Aseran.
Han krossade ock den kopparorm som Mose hade gjort; ty ända till denna tid hade Israels barn tänt offereld åt denne.
Man kallade honom Nehustan.
På HERREN, Israels Gud, förtröstade han, så att ingen var honom lik bland alla Juda konungar efter honom, ej heller bland dem som hade varit före honom.
Han höll sig till HERREN och vek icke av ifrån honom, utan höll hans bud, dem som HERREN hade givit Mose.
Och HERREN var med honom, så att han hade framgång i allt vad han företog sig.
Han avföll från konungen i Assyrien och upphörde att vara honom underdånig.
Han slog ock filistéerna och intog deras land ända till Gasa med dess område, såväl väktartorn som befästa städer.
I konung Hiskias fjärde regeringsår, som var Hoseas, Elas sons, Israels konungs, sjunde regeringsår, drog Salmaneser, konungen i Assyrien, upp mot Samaria och belägrade det.
Och de intogo det efter tre år, i Hiskias sjätte regeringsår; under detta år, som var Hoseas, Israels konungs, nionde regeringsår, blev Samaria intaget.
Och konungen i Assyrien förde Israel bort till Assyrien och förflyttade dem till Hala och till Habor, en ström i Gosan, och till Mediens städer --
detta därför att de icke hörde HERRENS, sin Guds, röst, utan överträdde hans förbund, allt vad HERRENS tjänare Mose hade bjudit; de ville varken höra eller göra det.
Och i konung Hiskias fjortonde regeringsår drog Sanherib, konungen i Assyrien, upp och angrep alla befästa städer i Juda och intog dem.
Då sände Hiskia, Juda konung, till Assyriens konung i Lakis och lät säga: »Jag har försyndat mig; vänd om och lämna mig i fred.
Vad du lägger på mig vill jag bära.»
Då ålade konungen i Assyrien Hiskia, Juda konung, att betala tre hundra talenter silver och trettio talenter guld.
Och Hiskia gav ut alla de penningar som funnos i HERRENS hus och i konungshusets skattkamrar.
Vid detta tillfälle lösbröt ock Hiskia från dörrarna till HERRENS tempel och från dörrposterna den beläggning som Hiskia, Juda konung, hade överdragit dem med, och gav detta åt konungen i Assyrien.
Men konungen i Assyrien sände från Lakis åstad Tartan, Rab-Saris och Rab-Sake med en stor här mot konung Hiskia i Jerusalem.
Dessa drogo då upp och kommo till Jerusalem; och när de hade dragit ditupp och kommit fram, stannade de vid Övre dammens vattenledning, på vägen till Valkarfältet.
Och de begärde att få tala med konungen.
Då gingo överhovmästaren Eljakim, Hilkias son, och sekreteraren Sebna och kansleren Joa, Asafs son, ut till dem.
Och Rab-Sake sade till dem: »Sägen till Hiskia: Så säger den store konungen, konungen i Assyrien: Vad är det för en förtröstan som du nu har hängivit dig åt?
Du menar väl att allenast munväder behövs för att veta råd och hava makt att föra krig.
På vem förtröstar du då, eftersom du har satt dig upp mot mig?
Du förtröstar val nu på den bräckta rörstaven Egypten, men se, när någon stöder sig på den, går den in i hans hand och genomborrar den.
Ty sådan är Farao, konungen i Egypten, för alla som förtrösta på honom.
Eller sägen I kanhända till mig: 'Vi förtrösta på HERREN, vår Gud'?
Var det då icke hans offerhöjder och altaren Hiskia avskaffade, när han sade till Juda och Jerusalem: 'Inför detta altare skolen I tillbedja, har i Jerusalem'?
Men ingå nu ett vad med min herre, konungen i Assyrien: jag vill giva dig två tusen hästar, om du kan skaffa dig ryttare till dem.
Huru skulle du då kunna slå tillbaka en enda ståthållare, en av min herres ringaste tjänare?
Och du sätter din förtröstan till Egypten, i hopp om att så få vagnar och ryttare!
Menar du då att jag utan HERRENS vilja har dragit upp till detta ställe för att fördärva det?
Nej, det är HERREN som har sagt till mig: Drag upp mot detta land och fördärva det.»
Då sade Eljakim, Hilkias son, och Sebna och Joa till Rab-Sake: »Tala till dina tjänare på arameiska, ty vi förstå det språket, och tala icke med oss på judiska inför folket som står på muren.»
Men Rab-Sake svarade dem: »Är det då till din herre och till dig som min herre har sänt mig att tala dessa ord?
Är det icke fastmer till de män som sitta på muren, och som jämte eder skola nödgas äta sin egen träck och dricka sitt eget vatten?»
Därefter trädde Rab-Sake närmare och ropade med hög röst på judiska och talade och sade: »Hören den store konungens, den assyriske konungens, ord.
Så säger konungen: Låten icke Hiskia bedraga eder, ty han förmår icke rädda eder ur min hand
Och låten icke Hiskia förleda eder att förtrösta på HERREN, därmed att han säger: 'HERREN skall förvisso rädda oss, och denna stad skall icke bliva given i den assyriske konungens hand.'
Hören icke på Hiskia.
Ty så säger konungen i Assyrien: Gören upp i godo med mig och given eder åt mig, så skolen I få äta var och en av sitt vinträd och av sitt fikonträd och dricka var och en ur sin brunn,
till dess jag kommer och hämtar eder till ett land som är likt edert eget land, ett land med säd och vin, ett land med bröd och vingårdar, ett land med ädla olivträd och honung; så skolen I få leva och icke dö.
Men hören icke på Hiskia; ty han vill förleda eder, när han säger: 'HERREN skall rädda oss.'
Har väl någon av de andra folkens gudar någonsin räddat sitt land ur den assyriske konungens hand?
Var äro Hamats och Arpads gudar?
Var äro Sefarvaims, Henas och Ivas gudar?
Eller hava de räddat Samaria ur min hand?
Vilken bland andra länders alla gudar har väl räddat sitt land ur min hand, eftersom I menen att HERREN skall rädda Jerusalem ur min hand?»
Men folket teg och svarade honom icke ett ord, ty konungen hade så bjudit och sagt: »Svaren honom icke.»
Och överhovmästaren Eljakim, Hilkias son, och sekreteraren Sebna och kansleren Joa, Asafs son, kommo till Hiskia med sönderrivna kläder och berättade för honom vad Rab-Sake hade sagt.
Då nu konung Hiskia hörde detta, rev han sönder sina kläder och höljde sig i sorgdräkt och gick in i HERRENS hus.
Och överhovmästaren Eljakim och sekreteraren Sebna och de äldste bland prästerna sände han, höljda i sorgdräkt, till profeten Jesaja, Amos' son.
Och de sade till denne: »Så säger Hiskia: En nödens, tuktans och smälekens dag är denna dag, ty fostren hava väl kommit fram till födseln, men kraft att föda finnes icke.
Kanhända skall HERREN, din Gud, höra alla Rab-Sakes ord, med vilka hans herre, konungen i Assyrien, har sänt honom till att smäda den levande Guden, så att han straffar honom för dessa ord, som han, HERREN, din Gud, har hört.
Så bed nu en bön för den kvarleva som ännu finnes.»
När nu konung Hiskias tjänare kommo till Jesaja,
sade Jesaja till dem: »Så skolen I säga till eder herre: Så säger HERREN: Frukta icke för de ord som du har hört, dem med vilka den assyriske konungens tjänare hava hädat mig.
Se, jag skall låta en sådan ande komma in i honom, att han, på grund av ett rykte som han skall få höra, vänder tillbaka till sitt land; och jag skall låta honom falla för svärd i hans eget land.
Och Rab-Sake vände tillbaka och fann den assyriske konungen upptagen med att belägra Libna; ty han hade hört att han hade brutit upp från Lakis.
Men när Sanherib fick höra säga om Tirhaka, konungen i Etiopien, att denne hade dragit ut för att strida mot honom, skickade han åter sändebud till Hiskia och sade:
»Så skolen I säga till Hiskia, Juda konung: Låt icke din Gud, som du förtröstar på, bedraga dig, i det att du tänker: 'Jerusalem skall icke bliva givet i den assyriske konungens hand.'
Du har nu hört vad konungarna i Assyrien hava gjort med alla andra länder, huru de hava givit dem till spillo.
Och du skulle nu bliva räddad!
Hava väl de folk som mina fäder fördärvade, Gosan, Haran, Resef och Edens barn i Telassar, blivit räddade av sina gudar?
Var är Hamats konung och Arpads konung och konungen över Sefarvaims stad, över Hena och Iva?»
När Hiskia hade mottagit brevet av sändebuden och läst det, gick han upp i HERRENS hus, och där bredde Hiskia ut det inför HERRENS ansikte.
Och Hiskia bad inför HERRENS ansikte och sade: »HERRE, Israels Gud, du som tronar på keruberna, du allena är Gud, den som råder över alla riken på jorden; du har gjort himmel och jord.
HERRE, böj ditt öra härtill och hör; HERRE, öppna dina ögon och se.
Ja, hör Sanheribs ord, det budskap varmed han har smädat den levande Guden.
Det är sant, HERRE, att konungarna i Assyrien hava förött folken och deras land.
Och de hava kastat deras gudar i elden; ty dessa voro inga gudar, utan verk av människohänder, trä och sten; därför kunde de förgöra dem.
Men fräls oss nu, HERRE, vår Gud, ur hans hand, så att alla riken på jorden förnimma att du, HERRE, allena är Gud.»
Då sände Jesaja, Amos' son, bud till Hiskia och låt säga: »Så säger HERREN, Israels Gud: Det varom du har bett mig angående Sanherib, konungen i Assyrien, det har jag hört.
Så är nu detta det ord som HERREN har talat om honom: Hon föraktar dig och bespottar dig, jungfrun dottern Sion; hon skakar huvudet efter dig, dottern Jerusalem.
vem har du smädat och hädat, och mot vem har du upphävt din röst?
Alltför högt har du upplyft dina ögon -- Ja, mot Israels Helige.
Genom dina sändebud smädade du Herren, när du sade: 'Med mina många vagnar drog jag upp på bergens höjder, längst upp på Libanon; jag högg ned dess höga cedrar och väldiga cypresser; jag trängde fram till dess innersta gömslen, dess frodigaste skog;
jag grävde brunnar och drack ut främmande vatten, och med min fot uttorkade jag alla Egyptens strömmar.'
Har du icke hört att jag för länge sedan beredde detta?
Av ålder bestämde jag ju så; och nu har jag fört det fram: du fick makt att ödelägga befästa städer till grusade stenhopar.
Deras invånare blevo maktlösa, de förfärades och stodo med skam.
Det gick dem såsom gräset på marken och gröna örter, såsom det som växer på taken, och säd som förbrännes, förrän strået har vuxit upp.
Om du sitter eller går ut eller går in, så vet jag det, och huru du rasar mot mig.
Men då du nu så rasar mot mig, och då ditt övermod har nått till mina öron, skall jag sätta min krok i din näsa och mitt betsel i din mun och föra dig tillbaka samma väg som du har kommit på.
Och detta skall för dig vara tecknet: man skall detta år äta vad som växer upp av spillsäd, och nästa år självvuxen säd; men det tredje året skolen I få så och skörda och plantera vingårdar och äta deras frukt.
Och den räddade skara av Juda hus, som bliver kvar, skall åter skjuta rot nedtill och bära frukt upptill.
Ty från Jerusalem skall utgå en kvarleva, en räddad skara från Sions berg.
HERRENS nitälskan skall göra detta.
Därför säger HERREN så om konungen i Assyrien: Han skall icke komma in i denna stad och icke skjuta någon pil ditin; han skall icke mot den föra fram någon sköld eller kasta upp någon vall mot den.
Samma väg han kom skall han vända tillbaka, och in i denna stad skall han icke komma, säger HERREN.
Ty jag skall beskärma och frälsa denna stad för min och min tjänare Davids skull.»
Och samma natt gick HERRENS ängel ut och slog i assyriernas läger ett hundra åttiofem tusen man; och när man bittida följande morgon kom ut, fick man se döda kroppar ligga där överallt
Då bröt Sanherib, konungen i Assyrien, upp och tågade tillbaka; och han stannade sedan i Nineve.
Men när han en gång tillbad i sin gud Nisroks tempel, blev han dräpt med svärd av Adrammelek och Sareser; därefter flydde dessa undan till Ararats land.
Och hans son Esarhaddon blev konung efter honom.
Vid den tiden blev Hiskia dödssjuk; och profeten Jesaja, Amos' son, kom till honom och sade till honom: »Så säger HERREN: Beställ om ditt hus; ty du måste dö och skall icke tillfriskna.»
Då vände han sitt ansikte mot väggen och bad till HERREN och sade:
»Ack HERRE, tänk dock på huru jag har vandrat inför dig i trohet och med hängivet hjärta och gjort vad gott är i dina ögon.»
Och Hiskia grät bitterligen.
Men innan Jesaja hade hunnit ut ur den inre staden, kom HERRENS ord till honom; han sade:
»Vänd om och säg till Hiskia, fursten över mitt folk: Så säger HERREN, din fader Davids Gud: Jag har hört din bön, jag har sett dina tårar.
Se, jag vill göra dig frisk; i övermorgon skall du få gå upp i HERRENS hus.
Och jag skall föröka din livstid med femton år; jag skall ock rädda dig och denna stad ur den assyriske konungens hand.
Ja, jag skall beskärma denna stad, för min skull och för min tjänare Davids skull.
Och Jesaja sade: »Hämten hit en fikonkaka.»
Då hämtade man en sådan och lade den på bulnaden.
Och han tillfrisknade.
Och Hiskia sade till Jesaja: »Vad för ett tecken gives mig därpå att HERREN skall göra mig frisk, så att jag i övermorgon får gå upp i HERRENS hus?»
Jesaja svarade: »Detta skall för dig vara tecknet från HERREN därpå att HERREN skall göra vad han har lovat: skuggan har gått tio steg framåt; skall den nu gå tio steg tillbaka?»
Hiskia sade: »Det är lätt för skuggan att sträcka sig tio steg framåt.
Nej, låt skuggan gå tio steg tillbaka.»
Då ropade profeten Jesaja till HERREN, och han lät skuggan på Ahas' solvisare gå tillbaka de tio steg som den redan hade lagt till rygga.
Vid samma tid sände Berodak-Baladan, Baladans son, konungen i Babel, brev och skänker till Hiskia, ty han hade sport att Hiskia hade varit sjuk.
Och när Hiskia hade hört på dem, visade han dem hela sitt förrådshus, sitt silver och guld, sina välluktande kryddor och sina dyrbara oljor, och hela sitt tyghus och allt vad som fanns i hans skattkamrar.
Intet fanns i Hiskias hus eller eljest i hans ägo, som han icke visade dem.
Men profeten Jesaja kom till konung Hiskia och sade till honom: »Vad hava dessa män sagt, och varifrån hava de kommit till dig?»
Hiskia svarade: »De hava kommit ifrån fjärran land, ifrån Babel.»
Han sade vidare: »Vad hava de sett i ditt hus?»
Hiskia svarade: »Allt som är i mitt hus hava de sett; intet finnes i mina skattkamrar, som jag icke har visat dem.»
Då sade Jesaja till Hiskia: »Hör HERRENS ord:
Se, dagar skola komma, då allt som finnes i ditt hus, och som dina fäder hava samlat ända till denna dag skall föras bort till Babel; intet skall bliva kvar, säger HERREN.
Och söner till dig, de som skola utgå av dig, och som du skall föda, dem skall man taga, och de skola bliva hovtjänare i den babyloniske konungens palats.»
Hiskia sade till Jesaja: »Gott är det HERRENS ord som du har talat.»
Och han sade ytterligare: »Ja, om nu blott frid och trygghet få råda i min tid.»
Vad nu mer är att säga om Hiskia och om alla hans bedrifter, och om huru han anlade dammen och vattenledningen och ledde vatten in i staden, det finnes upptecknat Juda konungars krönika.
Och Hiskia gick till vila hos sina fäder.
Och hans son Manasse blev konung efter honom.
Manasse var tolv år gammal, när han blev konung, och han regerade femtiofem år i Jerusalem.
Hans moder hette Hefsi-Ba.
Han gjorde vad ont var i HERRENS ögon, efter den styggeliga seden hos de folk som HERREN hade fördrivit för Israels barn.
Han byggde åter upp de offerhöjder som hans fader Hiskia hade förstört, och reste altaren åt Baal och gjorde en Asera, likasom Ahab, Israels konung, hade gjort, och tillbad och tjänade himmelens hela härskara.
Ja, han byggde altaren i HERRENS hus, det om vilket HERREN hade sagt: »Vid Jerusalem vill jag fästa mitt namn.»
Han byggde altaren åt himmelens hela härskara på de båda förgårdarna till HERRENS hus.
Han lät ock sin son gå genom eld och övade teckentyderi och svartkonst och skaffade sig andebesvärjare och spåmän och gjorde mycket som var ont i HERRENS ögon, så att han förtörnade honom.
Och Aserabelätet som han hade låtit göra satte han i det hus om vilket HERREN hade sagt till David och till hans son Salomo: »Vid detta hus och vid Jerusalem som jag har utvalt bland alla Israels stammar, vill jag fästa mitt namn för evig tid
Och jag skall icke mer låta Israel vandra flyktig bort ifrån det land som jag har givit åt deras fäder, om de allenast hålla och göra allt vad jag har bjudit dem, och det alldeles efter den lag som min tjänare Mose har givit dem.»
Men de lyssnade icke härtill, och Manasse förförde dem, så att de gjorde mer ont än de folk som HERREN hade förgjort för Israels barn.
Då talade HERREN genom sina tjänare profeterna och sade:
»Eftersom Manasse, Juda konung, har bedrivit dessa styggelser och så gjort mer ont, än allt vad amoréerna som voro före honom hava gjort, så att han med sina eländiga avgudar har kommit också Juda att synda,
därför säger HERREN, Israels Gud, så: 'Se, jag skall låta en sådan olycka komma över Jerusalem och Juda, att det skall genljuda i båda öronen på var och en som får höra det.
Och mot Jerusalem skall jag bruka det mätsnöre som jag brukade mot Samaria, och det sänklod som jag brukade mot Ahabs hus; och jag skall skölja Jerusalem tomt, såsom man sköljer ett fat och, sedan man har sköljt det, vänder det upp och ned.
Och jag skall förskjuta kvarlevan av min arvedel och giva dem i deras fienders hand, så att de skola bliva ett rov och ett byte för alla sina fiender --
detta därför att de hava gjort vad ont är i mina ögon och beständigt förtörnat mig, från den dag då deras fader drogo ut ur Egypten ända till denna dag.'»
Därtill utgöt ock Manasse oskyldigt blod i så stor myckenhet, att han därmed uppfyllde Jerusalem från den ena ändan till den andra -- detta förutom den särskilda syns genom vilken han kom Juda att synda och göra vad ont var i HERRENS ögon.
Vad nu mer är att säga om Manasse och om allt vad han gjorde så ock om den synd han begick det finnes upptecknat i Juda konungars krönika.
Och Manasse gick till vila hos sina fäder och blev begraven i trädgården till sitt hus, i Ussas trädgård.
Och hans son Amon blev konung efter honom.
Amon var tjugutvå år gammal när han blev konung, och han regerade två år i Jerusalem.
Hans moder hette Mesullemet, Harus' dotter, från Jotba.
Han gjorde vad ont var i HERRENS ögon, såsom hans fader Manasse hade gjort.
Han vandrade i allt på samma väg som hans fader hade vandrat, och tjänade och tillbad de eländiga avgudar som hans fader hade tjänat.
Han övergav HERREN, sina fäders Gud, och vandrade icke på HERRENS väg.
Och Amons tjänare sammansvuro sig mot honom och dödade konungen hemma i hans hus.
Men folket i landet dräpte alla som hade sammansvurit sig mot konung Amon.
Därefter gjorde folket i landet hans son Josia till konung efter honom.
Vad nu mer är att säga om Amon, om vad han gjorde, det finnes upptecknat i Juda konungars krönika.
Och man begrov honom i hans grav i Ussas trädgård.
Och hans son Josia blev konung efter honom.
Josia var åtta år gammal, när han blev konung, och han regerade trettioett år i Jerusalem.
Hans moder hette Jedida, Adajas dotter, från Boskat.
Han gjorde vad rätt var i HERRENS ögon och vandrade i allt på sin fader Davids väg och vek icke av vare sig till höger eller till vänster.
I sitt adertonde regeringsår sände konung Josia sekreteraren Safan, son till Asalja, Mesullams son, åstad till HERRENS hus och sade:
»Gå upp till översteprästen Hilkia, och bjud honom att göra i ordning de penningar som hava influtit till HERRENS hus, sedan de hava blivit insamlade ifrån folket av dem som hålla vakt vid tröskeln.
Och han skall överlämna dem åt de män som förrätta arbete såsom tillsyningsmän vid HERRENS hus, och dessa skola giva dem åt de män som arbeta vid HERRENS hus, för att sätta i stånd vad som är förfallet på huset,
nämligen åt timmermännen, byggningsmännen och murarna, så ock till att inköpa trävirke och huggen sten för att sätta huset i stånd.
Dock skall man icke hålla någon räkenskap med dem angående de penningar som överlämnas åt dem, utan de skola få handla på heder och tro.»
Och översteprästen Hilkia sade till sekreteraren Safan: »Jag har funnit lagboken i HERRENS hus.»
Och Hilkia gav boken åt Safan, och han läste den.
Därefter gick sekreteraren Safan in till konungen och avgav sin berättelse inför konungen; han sade: »Dina tjänare hava tömt ut de penningar som funnos i templet, och hava överlämnat dem åt de män som förrätta arbete såsom tillsyningsmän vid HERRENS hus.»
Vidare berättade sekreteraren Safan för konungen och sade: »Prästen Hilkia har givit mig en bok.»
Och Safan föreläste den för konungen.
När konungen nu hörde lagbokens ord, rev han sönder sina kläder.
Och konungen bjöd prästen Hilkia och Ahikam, Safans son, och Akbor, Mikajas son, och sekreteraren Safan och Asaja, konungens tjänare, och sade:
»Gån och frågen HERREN för mig och för folket, ja, för hela Juda, angående det som står i denna bok som nu har blivit funnen.
Ty stor är HERRENS vrede, den som är upptänd mot oss, därför att våra fäder icke hava velat lyssna till denna boks ord och icke hava gjort allt som är oss föreskrivet.
Då gingo prästen Hilkia och Ahikam, Akbor, Safan och Asaja till profetissan Hulda, hustru åt Sallum, klädkammarvaktaren, som var son till Tikva, Harhas' son; hon bodde i Jerusalem, i Nya staden.
Och de talade med henne.
Då sade hon till dem: »Så säger HERREN, Israels Gud: Sägen till den man som har sänt eder till mig:
Så säger HERREN: Se, över denna plats och över dess invånare skall jag låta olycka komma, allt vad som står i den bok som Juda konung har läst --
detta därför att de hava övergivit mig och tänt offereld åt andra gudar, och så hava förtörnat mig med alla sina händers verk.
Min vrede skall upptändas mot denna plats och skall icke bliva utsläckt.
Men till Juda konung, som har sänt eder för att fråga HERREN, till honom skolen I säga så: Så säger HERRES, Israels Gud,
angående de ord som du har hört: Eftersom ditt hjärta blev bevekt och du ödmjukade dig inför HERREN, när du hörde vad jag har talat mot denna plats och mot dess invånare, nämligen att de skola bliva ett föremål för häpnad och ett exempel som man nämner, när man förbannar, och eftersom du rev sönder dina kläder och grät inför mig, fördenskull har jag ock hört dig, säger HERREN.
Därför vill jag samla dig till dina fäder, så att du får samlas till dem i din grav med frid; och dina ögon skola slippa att se all den olycka som jag skall låta komma över denna plats.»
Och de vände till baka till konungen med detta svar.
Då sände konungen åstad män som församlade till honom alla de äldste i Juda och Jerusalem.
Och konungen gick upp i HERRENS hus, och alla Juda män och alla Jerusalems invånare följde honom, också prästerna och profeterna, ja, allt folket, ifrån den minste till den störste.
Och han läste upp för dem allt vad som stod i förbundsboken, som hade blivit funnen i HERRENS hus
Och konungen trädde fram till pelaren och slöt inför HERRENS ansikte det förbundet, att de skulle följa efter HERREN och hålla hans bud, hans vittnesbörd och hans stadgar, av allt hjärta och av all själ, och upprätthålla detta förbunds ord, dem som voro skrivna i denna bok.
Och allt folket trädde in i förbundet.
Därefter bjöd konungen översteprästen Hilkia och prästerna näst under honom, så ock dem som höllo vakt vid tröskeln, att de skulle föra bort ur HERRENS tempel alla de redskap som voro gjorda åt Baal och Aseran och åt himmelens hela härskara.
Och han lät bränna upp dem utanför Jerusalem på Kidrons fält, men askan efter dem lät han föra till Betel.
Han avsatte ock de avgudapräster som Juda konungar hade tillsatt, för att tända offereld på offerhöjderna i Juda städer och runt omkring Jerusalem, så ock dem som tände offereld åt Baal, åt solen, åt månen, åt stjärnbilderna och åt himmelens hela härskara.
Och han tog Aseran ur HERRENS hus och förde bort den utanför Jerusalem till Kidrons dal, och brände upp den där i Kidrons dal, han stötte sönder den till stoft och kastade stoftet på den allmänna begravningsplatsen.
Vidare rev han ned tempelbolarhusen som funnos i HERRENS hus, dem i vilka kvinnor vävde tyg till tält åt Aseran.
Och han lät föra alla prästerna bort ifrån Juda städer och orenade de offerhöjder där prästerna hade tänt offereld, från Geba ända till Beer-Seba; och han bröt ned offerhöjderna vid stadsportarna, både den som låg vid ingången till stadshövitsmannen Josuas port och den som låg till vänster, när man gick in genom stadsporten.
Dock fingo offerhöjdsprästerna icke stiga upp till HERRENS altare i Jerusalem; de fingo allenast äta osyrat bröd ibland sina bröder.
Han orenade ock Tofet i Hinnoms barns dal, för att ingen skulle låta sin son eller dotter gå genom eld, till offer åt Molok.
Och han skaffade bort de hästar som Juda konungar hade invigt åt solen och ställt upp så, att man icke kunde gå in i HERRENS hus, vid hovmannen Netan-Meleks kammare i Parvarim; och solens vagnar brände han upp i eld.
Och altarna på taket över Ahas' sal, vilka Juda konungar hade låtit göra, och de altaren som Manasse hade låtit göra på de båda förgårdarna till HERRENS hus, dem bröt konungen ned; sedan skyndade han bort därifrån och kastade stoftet av dem i Kidrons dal.
Och offerhöjderna öster om Jerusalem och söder om Fördärvets berg, vilka Salomo, Israels konung, hade byggt åt Astarte, sidoniernas styggelse, åt Kemos, Moabs styggelse, och åt Milkom, Ammons barns skändlighet, dem orenade konungen.
Han slog sönder stoderna och högg ned Aserorna; och platsen där de hade stått fyllde han med människoben.
Också altaret i Betel, den offerhöjd som Jerobeam, Nebats son, hade byggt upp, han som kom Israel att synda, också detta altare med offerhöjden bröt han ned; därefter brände han upp offerhöjden och stötte sönder den till stoft och brände tillika upp Aseran.
När då Josia såg sig om och fick se gravarna som voro där på berget, sände han åstad och lät hämta benen ur gravarna och brände upp dem på altaret och orenade det så -- i enlighet med det HERRENS ord som hade blivit förkunnat av gudsmannen som förkunnade att detta skulle ske.
Och han frågade: »Vad är det för en vård som jag ser där?»
Folket i staden svarade honom: »Det är den gudsmans grav, som kom från Juda och ropade mot altaret i Betel att det skulle ske, som du nu har gjort.»
Då sade han: »Låten honom vara; ingen må röra hans ben.»
Så lämnade man då hans ben i fred, och tillika benen av den profet som hade kommit dit från Samarien.
Därjämte skaffade Josia bort alla de offerhöjdshus i Samariens städer, som Israels konungar hade byggt upp, och med vilka de hade kommit förtörnelse åstad; och han gjorde med dem alldeles på samma sätt som han hade gjort i Betel.
Och alla offerhöjdspräster som funnos där slaktade han på altarna och brände människoben ovanpå dem.
Därefter vände han tillbaka till Jerusalem.
Och konungen bjöd allt folket och sade: »Hållen HERRENS, eder Guds, påskhögtid, såsom det är föreskrivet i denna förbundsbok.»
Ty en sådan påskhögtid hade icke blivit hållen sedan den tid då domarna dömde Israel, icke under Israels konungars och Juda konungars hela tid.
Först i konung Josias adertonde regeringsår hölls en sådan HERRENS påskhögtid i Jerusalem.
Därjämte skaffade Josia bort andebesvärjarna och spåmännen, husgudarna och de eländiga avgudarna, och alla styggelser som voro att se i Juda land och i Jerusalem, på det att han skulle upprätthålla lagens ord, dem som voro skrivna i den bok som prästen Hilkia hade funnit i HERRENS hus.
Ingen konung lik honom hade funnits före honom, ingen som så av allt sitt hjärta och av all sin själ och av all sin kraft hade vänt sig till HERREN, i enlighet med Moses hela lag; och efter honom uppstod ej heller någon som var honom lik.
Dock vände HERREN sig icke ifrån sin stora vredes glöd, då nu hans vrede hade blivit upptänd mot Juda, för allt det varmed Manasse hade förtörnat honom.
Och HERREN sade: »Också Juda vill jag förskjuta ifrån mitt ansikte, likasom jag har förskjutit Israel; ja, jag vill förkasta Jerusalem, denna stad som jag hade utvalt, så ock det hus varom jag hade sagt: Mitt namn skall vara där.»
Vad nu mer är att säga om Josia och om allt vad han gjorde, det finnes upptecknat i Juda konungars krönika.
I hans tid drog Farao Neko, konungen i Egypten, upp mot konungen i Assyrien, till floden Frat.
Då tågade konung Josia emot honom, men blev dödad av honom vid Megiddo, under första sammandrabbningen.
Och hans tjänare förde hans döda kropp i en vagn bort ifrån Megiddo till Jerusalem och begrovo honom i hans grav.
Men folket i landet tog Josias son Joahas och smorde honom och gjorde honom till konung efter hans fader.
Joahas var tjugutre år gammal, när han blev konung, och han regerade tre månader i Jerusalem.
Hans moder hette Hamutal, Jeremias dotter, från Libna.
Han gjorde vad ont var i HERRENS ögon, alldeles såsom hans fäder hade gjort.
Och Farao Neko lät sätta honom i fängelse i Ribla i Hamats land och gjorde så slut på hans regering i Jerusalem; och han pålade landet en skatt av ett hundra talenter silver och en talent guld.
Och Farao Neko gjorde Josias son Eljakim till konung i hans fader Josias ställe och förändrade hans namn till Jojakim.
Men Joahas tog han med sig, och denne kom så till Egypten och dog där.
Och Jojakim betalade ut silvret och guldet åt Farao; men han måste skattlägga landet för att kunna utbetala dessa penningar enligt Faraos befallning.
Efter som var och en av folket i landet blev uppskattad, indrevs från dem silvret och guldet, för att sedan utbetalas åt Farao Neko.
Jojakim var tjugufem år gammal, när han blev konung; och han regerade elva år i Jerusalem.
Hans moder hette Sebida, Pedajas dotter, från Ruma.
Han gjorde vad ont var i HERRENS ögon, alldeles såsom hans fäder hade gjort.
I hans tid drog Nebukadnessar, konungen i Babel, upp, och Jojakim blev honom underdånig och förblev så i tre år; men sedan avföll han från honom.
Då sände HERREN över honom kaldéernas; araméernas, moabiternas och Ammons barns härskaror; han sände dem över Juda för att förgöra det -- i enlighet med det ord som HERREN hade talat genom sina tjänare profeterna.
Ja, det var efter HERRENS ord som detta kom över Juda, i det att han försköt det från sitt ansikte för de synder Manasse hade begått och för allt vad denne hade förövat,
jämväl för det oskyldiga blod som han utgöt, ty han uppfyllde Jerusalem med oskyldigt blod; det ville HERREN icke förlåta.
Vad nu mer är att säga om Jojakim och om allt vad han gjorde, det finnes upptecknat i Juda konungars krönika.
Och Jojakim gick till vila hos sina fäder.
Och hans son Jojakin blev konung efter honom.
Därefter drog konungen i Egypten icke vidare ut ur sitt land, ty konungen i Babel hade intagit allt som tillhörde konungen i Egypten, från Egyptens bäck ända till floden Frat.»
Jojakin var aderton år gammal, när han blev konung, och han regerade tre månader i Jerusalem.
Hans moder hette Nehusta, Elnatans dotter, från Jerusalem.
Han gjorde vad ont var i HERRENS ögon, alldeles såsom hans fader hade gjort.
På den tiden drogo den babyloniske konungen Nebukadnessars tjänare upp till Jerusalem, och staden blev belägrad.
Och Nebukadnessar, konungen i Babel, kom till staden, medan hans tjänare belägrade den.
Då gav sig Jojakin, Juda konung, åt konungen i Babel, med sin moder och med sina tjänare, sina hövitsmän och hovmän; och konungen i Babel tog honom så till fånga i sitt åttonde regeringsår.
Och han förde bort därifrån alla skatter i HERRENS hus och skatterna i konungshuset, han lösbröt ock beläggningen från alla gyllene föremål som Salomo, Israels konung, hade låtit göra för HERRENS tempel, detta i enlighet med vad HERREN hade hotat.
Och han förde bort i fångenskap hela Jerusalem, alla hövitsmän och alla tappra stridsmän; tio tusen förde han bort, jämväl alla timmermän och smeder.
Inga andra lämnades kvar än de ringaste av folket i landet.
Han förde Jojakin bort till Babel; därjämte förde han konungens moder, konungens hustrur och hans hovmän samt de mäktige i landet såsom fångar bort ifrån Jerusalem till Babel,
så ock alla stridsmännen, sju tusen, och timmermännen och smederna, ett tusen, allasammans raska och krigsdugliga män.
Dessa fördes nu av den babyloniske konungen i fångenskap till Babel.
Men konungen i Babel gjorde hans farbroder Mattanja till konung i hans ställe och förändrade dennes namn till Sidkia.
Sidkia var tjuguett år gammal, när han blev konung, och han regerade elva år i Jerusalem.
Hans moder hette Hamital, Jeremias dotter, från Libna.
Han gjorde vad ont var i HERRENS ögon, alldeles såsom Jojakim hade gjort.
Ty på grund av HERRENS vrede skedde vad som skedde med Jerusalem och Juda, till dess att han kastade dem bort ifrån sitt ansikte.
Då, i hans nionde regeringsår, i tionde månaden; på tionde dagen i månaden, kom Nebukadnessar, konungen i Babel, med hela sin här till Jerusalem och belägrade det; och de byggde en belägringsmur runt omkring det.
Så blev staden belägrad och förblev så ända till konung Sidkias elfte regeringsår.
Men på nionde dagen i månaden var hungersnöden så stor i staden, att mängden av folket icke hade något att äta.
Och staden stormades, och allt krigsfolket flydde om natten genom porten mellan de båda murarna (den port som ledde till den kungliga trädgården), medan kaldéerna lågo runt omkring staden; och folket tog vägen åt Hedmarken till.
Men kaldéernas här förföljde konungen, och de hunno upp honom på Jerikos hedmarker, sedan hela hans här hade övergivit honom och skingrat sig.
Och de grepo konungen och förde honom till den babyloniske konungen i Ribla; där höll man rannsakning och dom med honom.
Och Sidkias barn slaktade man inför hans ögon, och på Sidkia själv stack man ut ögonen; och man fängslade honom med kopparfjättrar och förde honom till Babel.
I femte månaden, på sjunde dagen i månaden, detta i den babyloniske konungen Nebukadnessars nittonde regeringsår, kom den babyloniske konungens tjänare Nebusaradan, översten för drabanterna, till Jerusalem.
Denne brände upp HERRENS hus och konungshuset: ja, alla hus i Jerusalem, i synnerhet alla de förnämas hus, brände han upp i eld.
Och murarna runt omkring Jerusalem brötos ned av hela den här av kaldéer, som översten för drabanterna hade med sig,
och återstoden av folket, dem som voro kvar i staden, och de överlöpare som hade gått över till konungen i Babel, så ock den övriga hopen, dem förde Nebusaradan, översten för drabanterna, bort i fångenskap.
Men av de ringaste i landet lämnade översten för drabanterna några kvar till vingårdsmän och åkermän.
Kopparpelarna i HERRENS hus, bäckenställen och kopparhavet i HERRENS hus slogo kaldéerna sönder och förde kopparen till Babel.
Och askkärlen, skovlarna, knivarna, skålarna och alla kopparkärl som hade begagnats vid gudstjänsten togo de bort.
Likaledes tog översten för drabanterna bort fyrfaten och offerskålarna, allt som var av rent guld eller av rent silver.
Vad angår de två pelarna, havet, som var allenast ett, och bäckenställen, som Salomo hade låtit göra till HERRENS hus, så kunde kopparen i alla dessa föremål icke vägas.
Aderton alnar hög var den ena pelaren, och ovanpå den var ett pelarhuvud av koppar, och pelarhuvudet var tre alnar högt, och ett nätverk och granatäpplen funnos på pelarhuvudet runt omkring, alltsammans av koppar; och likadant var det på den andra pelaren, över nätverket.
Och översten för drabanterna tog översteprästen Seraja jämte Sefanja, prästen näst under honom, så ock de tre som höllo vakt vid tröskeln,
och från staden tog han en hovman, den som var anförare för krigsfolket, och fem av konungens närmaste män, som påträffades i staden, så ock sekreteraren, den härhövitsman som plägade utskriva folket i landet till krigstjänst, och sextio andra män av landets folk, som påträffades i staden --
dessa tog Nebusaradan, översten för drabanterna, och förde dem till den babyloniske konungen i Ribla.
Och konungen i Babel lät avliva dem där, i Ribla i Hamats land. blev Juda bortfört från sitt land.
Men över det folk som blev kvar i Juda land, det folk som Nebukadnessar, konungen i Babel, lät bliva kvar där, satte han Gedalja, son till Ahikam, son till Safan.
När då alla krigshövitsmännen jämte sina män fingo höra att konungen i Babel hade satt Gedalja över landet, kommo de till Gedalja i Mispa, nämligen Ismael, Netanjas son, Johanan, Kareas son, netofatiten Seraja, Tanhumets son, och Jaasanja, maakatitens son, med sina män.
Och Gedalja gav dem och deras män sin ed och sade till dem: »Frukten icke för kaldéernas tjänare.
Stannen kvar i landet, och tjänen konungen i Babel, så skall det gå eder väl.»
Men i sjunde månaden kom Ismael, son till Netanja, son till Elisama, av konungslig börd, och hade med sig tio män, och de slogo ihjäl Gedalja, så ock de judar och kaldéer som voro hos honom i Mispa.
Då bröt allt folket upp, från den minste till den störste, tillika med krigshövitsmännen, och begav sig till Egypten; ty de fruktade för kaldéerna.
Men i det trettiosjunde året sedan Jojakin, Juda konung, hade blivit bortförd i fångenskap, i tolfte månaden, på tjugusjunde dagen i månaden, tog Evil-Merodak, konungen i Babel -- samma år han blev konung -- Jojakin, Juda konung, till nåder och befriade honom ur fängelset;
Och han talade vänligt med honom och gav honom främsta platsen bland de konungar som voro hos honom i Babel.
Han fick lägga av sin fångdräkt och beständigt äta vid hans bord, så länge han levde.
Och ett ständigt underhåll gavs honom från konungen, visst för var dag, så länge han levde.
Adam, Set, Enos,
Kenan, Mahalalel, Jered,
Hanok, Metusela, Lemek,
Noa, Sem, Ham och Jafet.
Jafets söner voro Gomer, Magog, Madai, Javan, Tubal, Mesek och Tiras.
Gomers söner voro Askenas, Difat och Togarma.
Javans söner voro Elisa och Tarsisa, kittéerna och rodanéerna.
Hams söner voro Kus, Misraim, Put och Kanaan.
Kus' söner voro Seba, Havila, Sabta, Raema och Sabteka.
Raemas söner voro Saba och Dedan.
Men Kus födde Nimrod; han var den förste som upprättade ett välde på jorden.
Och Misraim födde ludéerna, anaméerna, lehabéerna, naftuhéerna,
patroséerna, kasluhéerna, från vilka filistéerna hava utgått, och kaftoréerna.
Och Kanaan födde Sidon, som var hans förstfödde, och Het,
så ock jebuséerna, amoréerna och girgaséerna,
hivéerna, arkéerna, sinéerna,
arvadéerna, semaréerna och hamatéerna.
Sems söner voro Elam, Assur, Arpaksad, Lud och Aram, så ock Us, Hul, Geter och Mesek.
Arpaksad födde Sela, och Sela födde Eber.
Men åt Eber föddes två söner; den ene hette Peleg, ty i hans tid blev jorden fördelad; och hans broder hette Joktan.
Och Joktan födde Almodad, Selef, Hasarmavet, Jera,
Hadoram, Usal, Dikla,
Ebal, Abimael, Saba,
Ofir, Havila och Jobab; alla dessa voro Joktans söner.
Sem, Arpaksad, Sela,
Eber, Peleg, Regu,
Serug, Nahor, Tera,
Abram, det är Abraham
Abrahams söner voro Isak och Ismael.
Detta är deras släkttavla: Nebajot, Ismaels förstfödde, vidare Kedar, Adbeel och Mibsam,
Misma och Duma, Massa, Hadad och Tema,
Jetur, Nafis och Kedma.
Dessa voro Ismaels söner.
Och de söner som Ketura, Abrahams bihustru, födde voro Simran, Joksan, Medan, Midjan, Jisbak och Sua.
Joksans söner voro Saba och Dedan.
Och Midjans söner voro Efa, Efer, Hanok, Abida och Eldaa.
Alla dessa voro Keturas söner.
Och Abraham födde Isak.
Isaks söner voro Esau och Israel.
Esaus söner voro Elifas, Reguel, Jeus, Jaelam och Kora.
Elifas' söner voro Teman och Omar, Sefi och Gaetam, Kenas, Timna och Amalek
Reguels söner voro Nahat, Sera, Samma och Missa.
Men Seirs söner voro Lotan, Sobal, Sibeon, Ana, Dison, Eser och Disan.
Lotans söner voro Hori och Homam; och Lotans syster var Timna.
Sobals söner voro Aljan, Manahat och Ebal, Sefi och Onam.
Och Sibeons söner voro Aja och Ana.
Anas söner voro Dison.
Och Disons söner voro Hamran, Esban, Jitran och Keran.
Esers söner voro Bilhan, Saavan, Jaakan.
Disans söner voro Us och Aran.
Och dessa voro de konungar som regerade i Edoms land, innan ännu någon israelitisk konung var konung där: Bela, Beors son, och hans stad hette Dinhaba.
När Bela dog, blev Jobab, Seras son, från Bosra, konung efter honom.
När Jobab dog, blev Husam från temanéernas land konung efter honom.
När Husam dog, blev Hadad, Bedads son, konung efter honom, han som slog midjaniterna på Moabs mark; och hans stad hette Avit.
När Hadad dog, blev Samla från Masreka konung efter honom.
När Samla dog, blev Saul, från Rehobot vid floden, konung efter honom.
När Saul dog, blev Baal-Hanan, Akbors son, konung efter honom
När Baal-Hanan dog, blev Hadad konung efter honom; och hans stad hette Pagi, och hans hustru hette Mehetabel, dotter till Matred, var dotter till Me-Sahab.
Men när Hadad hade dött, voro dessa Edoms stamfurstar: fursten Timna, fursten Alja, fursten Jetet,
fursten Oholibama, fursten Ela, fursten Pinon,
fursten Kenas, fursten Teman, fursten Mibsar,
fursten Magdiel, fursten Iram.
Dessa voro Edoms stamfurstar.
Dessa voro Israels söner: Ruben, Simeon, Levi och Juda, Isaskar och Sebulon,
Dan, Josef och Benjamin, Naftali, Gad och Aser.
Judas söner voro Er, Onan och Sela; dessa tre föddes åt honom av Suas dotter, kananeiskan.
Men Er, Judas förstfödde, misshagade HERREN; därför dödade han honom.
Och Tamar, hans sonhustru, födde åt honom Peres och Sera, så att Judas söner voro tillsammans fem.
Peres' söner voro Hesron och Hamul.
Seras söner voro Simri, Etan, Heman, Kalkol och Dara, tillsammans fem.
Men Karmis söner voro Akar, som drog olycka över Israel, när han trolöst förgrep sig på det tillspillogivna.
Och Etans söner voro Asarja.
Och de söner som föddes åt Hesron voro Jerameel, Ram och Kelubai.
Och Ram födde Amminadab, och Amminadab födde Naheson, hövding för Juda barn.
Naheson födde Salma, och Salma födde Boas.
Boas födde Obed, och Obed födde Isai.
Isai födde Eliab, som var hans förstfödde, Abinadab, den andre, och Simea, den tredje,
Netanel, den fjärde, Raddai, den femte,
Osem, den sjätte, David, den sjunde.
Och deras systrar voro Seruja och Abigail.
Och Serujas söner voro Absai, Joab och Asael, tillsammans tre.
Och Abigail födde Amasa, och Amasas fader var ismaeliten Jeter.
Och Kaleb, Hesrons son, födde ett barn av kvinnkön, Asuba, därtill ock Jeriot; och dessa voro henne söner: Jeser, Sobab och Ardon.
Och när Asuba dog, tog Kaleb Efrat till hustru åt sig, och hon födde åt honom Hur.
Och Hur födde Uri, och Uri födde Besalel.
Därefter gick Hesron in till Makirs, Gileads faders, dotter; henne tog han till hustru, när han var sextio år gammal.
Och hon födde åt honom Segub.
Och Segub födde Jair; denne hade tjugutre städer i Gileads land.
Men gesuréerna och araméerna togo ifrån dem Jairs byar jämte Kenat med underlydande orter, sextio städer.
Alla dessa voro söner till Makir, Gileads fader.
Och sedan Hesron hade dött i Kaleb-Efrata, födde Hesrons hustru Abia åt honom Ashur, Tekoas fader.
Och Jerameels, Hesrons förstföddes, söner voro Ram, den förstfödde, vidare Buna, Oren och Osem samt Ahia.
Men Jerameel hade en annan hustru som hette Atara; hon var moder till Onam.
Och Rams, Jerameels förstföddes, söner voro Maas, Jamin och Eker.
Onams söner voro Sammai och Jada; och Sammais söner voro Nadab och Abisur.
Och Abisurs hustru hette Abihail; hon födde åt honom Aban och Molid.
Nadabs söner voro Seled och Appaim.
Seled dog barnlös.
Men Appaims söner voro Jisei; Jiseis söner voro Sesan; Sesans söner voro Alai.
Jadas, Sammais broders, söner voro Jeter och Jonatan.
Jeter dog barnlös.
Men Jonatans söner voro Pelet och Sasa.
Dessa voro Jerameels söner.
Men Sesan hade inga söner, utan allenast döttrar.
Nu hade Sesan en egyptisk tjänare som hette Jarha.
Och Sesan gav sin dotter till hustru åt sin tjänare Jarha, och hon födde åt honom Attai.
Attai födde Natan, och Natan födde Sabad.
Sabad födde Eflal, och Eflal födde Obed.
Obed födde Jehu, och Jehu födde Asarja.
Asarja födde Heles, och Heles födde Eleasa.
Eleasa födde Sisamai, och Sisamai födde Sallum.
Sallum födde Jekamja, och Jekamja födde Elisama.
Och Kalebs, Jerameels broders, söner voro Mesa, hans förstfödde, som var Sifs fader, och Maresas, Hebrons faders, söner.
Men Hebrons söner voro Kora, Tappua, Rekem och Sema.
Sema födde Raham, Jorkeams fader.
Men Rekem födde Sammai.
Sammais son var Maon, och Maon var Bet-Surs fader.
Och Efa, Kalebs bihustru, födde Haran, Mosa och Gases; och Haran födde Gases.
Och Jadais söner voro Regem, Jotam, Gesan, Pelet, Efa och Saaf.
Kalebs bihustru Maaka födde Seber och Tirhana.
Hon födde ock Saaf, Madmannas fader, Seva, Makbenas fader och Gibeas fader.
Och Kalebs dotter var Aksa.
Dessa voro Kalebs söner: Hurs, Efratas förstföddes, son var Sobal Kirjat-Jearims fader,
vidare Salma, Bet-Lehems fader, och Haref, Bet-Gaders fader.
Söner till Sobal, Kirjat-Jearims fader, voro Haroe och hälften av Hammenuhot-släkten.
Men Kirjat-Jearims släkter voro jeteriterna, putiterna, sumatiterna och misraiterna.
Från dem utgingo sorgatiterna och estaoliterna.
Salmas söner voro Bet-Lehem och netofatiterna, Atrot-Bet-Joab, så ock hälften av manahatiterna, sorgiterna.
Och de skriftlärdes släkter, deras som bodde i Jaebes, voro tireatiterna, simeatiterna, sukatiterna.
Dessa voro de kainéer som härstammade från Hammat, fader till Rekabs släkt.
Dessa voro de söner som föddes åt David i Hebron: Amnon, den förstfödde, av Ahinoam från Jisreel; Daniel, den andre, av Abigail från Karmel;
Absalom, den tredje, son till Maaka, som var dotter till Talmai, konungen i Gesur; Adonia, den fjärde, Haggits son;
Sefatja, den femte, av Abital; Jitream, den sjätte, av hans hustru Egla.
Dessa sex föddes åt honom i Hebron, där han regerade i sju år och sex månader.
I Jerusalem åter regerade han i trettiotre år.
Och dessa söner föddes åt honom i Jerusalem: Simea, Sobab, Natan och Salomo, tillsammans fyra, av Bat-Sua, Ammiels dotter;
vidare Jibhar, Elisama, Elifelet,
Noga, Nefeg, Jafia,
Elisama, Eljada och Elifelet, tillsammans nio.
Detta var alla Davids söner, förutom sönerna med bihustrurna; och Tamar var deras syster.
Salomos son var Rehabeam.
Hans son var Abia; hans son var Asa; hans son var Josafat.
Hans son var Joram; hans son var Ahasja; hans son var Joas.
Hans son var Amasja; hans son var Asarja; hans son var Jotam.
Hans son var Ahas; hans son var Hiskia; hans son var Manasse.
Hans son var Amon; hans son var Josia.
Josias söner voro Johanan den förstfödde, Jojakim, den andre, Sidkia, den tredje, Sallum, den fjärde.
Jojakims söner voro hans son Jekonja och dennes son Sidkia.
Jekonjas söner voro Assir och dennes son Sealtiel,
vidare Malkiram, Pedaja, Senassar, Jekamja, Hosama och Nedabja.
Pedajas söner voro Serubbabel och Simei.
Serubbabels söner voro Mesullam och Hananja, och deras syster var Selomit,
vidare Hasuba, Ohel, Berekja, Hasadja och Jusab-Hesed, tillsammans fem.
Hananjas söner voro Pelatja och Jesaja, vidare Refajas söner, Arnans söner, Obadjas söner och Sekanjas söner.
Sekanjas söner voro Semaja, Semajas söner voro Hattus, Jigeal, Baria, Nearja och Safat, tillsammans sex.
Nearjas söner voro Eljoenai, Hiskia och Asrikam, tillsammans tre.
Eljoenais söner voro Hodauja, Eljasib, Pelaja, Ackub, Johanan, Delaja och Anani, tillsammans sju.
Judas söner voro Peres, Hesron, Karmi, Hur och Sobal.
Och Reaja, Sobals son, födde Jahat, och Jahat födde Ahumai och Lahad.
Dessa voro sorgatiternas släkter.
Och dessa voro Abi-Etams söner: Jisreel, Jisma och Jidbas, och deras syster hette Hasselelponi,
vidare Penuel, Gedors fader, och Eser, Husas fader.
Dessa voro söner till Hur, Efratas förstfödde, Bet-Lehems fader.
Och Ashur, Tekoas fader, hade två hustrur, Helea och Naara.
Naara födde åt honom Ahussam, Hefer, Timeni och ahastariterna.
Dessa voro Naaras söner.
Och Heleas söner voro Seret, Jishar och Etnan.
Och Kos födde Anub och Hassobeba, så ock Aharhels, Harums sons, släkter.
Men Jaebes var mer ansedd än sina bröder; hans moder hade givit honom namnet Jaebes, i det hon sade: »Jag har fött honom med smärta.»
Och Jaebes åkallade Israels Gud och sade: »O att du ville välsigna mig och utvidga mitt område och låta din hand vara med mig!
O att du ville avvända vad ont är, så att jag sluppe att känna någon smärta!»
Och Gud lät det ske, som han begärde.
Och Kelub, Suhas broder, födde Mehir; han var Estons fader.
Och Eston födde Bet-Rafa, Pasea och Tehinna, Ir-Nahas' fader.
Dessa voro männen från Reka.
Och Kenas söner voro Otniel och Seraja.
Otniels söner voro Hatat.
Och Meonotai födde Ofra.
Och Seraja födde Joab, fader till Timmermansdalens släkt, ty dessa voro timmermän.
Och Kalebs, Jefunnes sons, söner voro Iru, Ela och Naam, så ock Elas söner och Kenas.
Och Jehallelels söner voro Sif och Sifa, Tirja och Asarel.
Och Esras son var Jeter, vidare Mered, Efer och Jalon.
Och kvinnan blev havande och födde Mirjam, Sammai och Jisba, Estemoas fader.
Och hans judiska hustru födde Jered, Gedors fader, och Heber, Sokos fader, och Jekutiel, Sanoas fader.
Men de andra voro söner till Bitja, Faraos dotter, som Mered hade tagit till hustru.
Och söner till Hodias hustru, Nahams syster, voro Kegilas fader, garmiten, och maakatiten Estemoa.
Och Simons söner voro Amnon och Rinna, Ben-Hanan och Tilon.
Och Jiseis söner voro Sohet och Sohets son.
Söner till Sela, Judas son, voro Er, Lekas fader, och Laeda, Maresas fader, och de släkter som tillhörde linnearbetarnas hus, av Asbeas hus,
vidare Jokim och männen i Koseba samt Joas och Saraf, som blevo herrar över Moab, så ock Jasubi-Lehem.
Men detta tillhör en avlägsen tid.
Dessa voro krukmakarna och invånarna i Netaim och Gedera; de bodde där hos konungen och voro i hans arbete.
Simeons söner voro Nemuel och Jamin, Jarib, Sera och Saul.
Hans son var Sallum; hans son var Mibsam; hans son var Misma.
Mismas söner voro hans son Hammuel, dennes son Sackur och dennes son Simei.
Och Simei hade sexton söner och sex döttrar; men hans bröder hade icke många barn.
Och deras släkt i sin helhet förökade sig icke så mycket som Juda barn.
Och de bodde i Beer-Seba, Molada och Hasar-Sual,
i Bilha, i Esem och i Tolad,
i Betuel, i Horma och i Siklag,
i Bet-Markabot, i Hasar-Susim, i Bet-Birei och i Saaraim.
Dessa voro deras städer, till dess att David blev konung.
Och deras byar voro Etam och Ain, Rimmon, Token och Asan -- fem städer;
därtill alla deras byar, som lågo runt omkring dessa städer, ända till Baal.
Dessa voro deras boningsorter; och de hade sitt särskilda släktregister.
Vidare: Mesobab, Jamlek och Josa, Amasjas son,
och Joel och Jehu, son till Josibja, son till Seraja, son till Asiel,
och Eljoenai, Jaakoba, Jesohaja, Asaja, Adiel, Jesimiel och Benaja,
så ock Sisa, son till Sifei, son till Allon, son till Jedaja, son till Simri son till Semaja.
Dessa nu nämnda voro hövdingar i sina släkter, och deras familjer utbredde sig och blevo talrika.
Och de drogo fram mot Gedor, ända till östra sidan av dalen, för att söka bete för sin boskap.
Och de funno fett och gott bete, och landet hade utrymme nog, och där var stilla och lugnt, ty de som förut bodde där voro hamiter.
Men dessa som här hava blivit upptecknade vid namn kommo i Hiskias, Juda konungs, tid och förstörde deras tält och slogo de meiniter som funnos där och gåvo dem till spillo, så att de nu icke mer äro till, och bosatte sig i deras land; ty där fanns bete för deras boskap.
Och av dem, av Simeons barn, drogo fem hundra man till Seirs bergsbygd; och Pelatja, Nearja, Refaja och Ussiel, Jiseis söner, stodo i spetsen för dem.
Och de slogo den sista kvarlevan av amalekiterna; sedan bosatte de sig där och bo där ännu i dag.
Och Rubens söner, Israels förstföddes -- han var nämligen den förstfödde, men därför att han oskärade sin faders bädd, blev hans förstfödslorätt given åt Josefs, Israels sons, söner, dock icke så, att denne skulle upptagas i släktregistret såsom den förstfödde;
ty väl var Juda den mäktigaste bland sina bröder, och furste blev en av hans avkomlingar, men förstfödslorätten blev dock Josefs --
Rubens, Israels förstföddes, söner voro Hanok och Pallu, Hesron och Karmi.
Joels söner voro hans son Semaja, dennes son Gog, dennes son Simei,
dennes son Mika, dennes son Reaja, dennes son Baal,
så ock dennes son Beera, som Tillegat-Pilneeser, konungen i Assyrien, förde bort i fångenskap; han var hövding för rubeniterna.
Och hans bröder voro, efter sina släkter, när de upptecknades i släktregistret efter sin ättföljd: Jegiel, huvudmannen, Sakarja
och Bela, son till Asas, son till Sema, son till Joel; han bodde i Aroer, och hans boningsplatser nådde ända till Nebo och Baal-Meon.
Och österut nådde hans boningsplatser ända fram till öknen som sträcker sig ifrån floden Frat; ty de hade stora boskapshjordar i Gileads land.
Men i Sauls tid förde de krig mot hagariterna, och dessa föllo för deras hand; då bosatte de sig i deras hyddor utefter hela östra sidan av Gilead.
Och Gads barn hade sina boningsplatser gent emot dem i landet Basan ända till Salka:
Joel, huvudmannen, och Safam därnäst, och vidare Jaanai och Safat i Basan.
Och deras bröder voro, efter sina familjer, Mikael, Mesullam, Seba, Jorai, Jaekan, Sia och Eber, tillsammans sju.
Dessa voro söner till Abihail, son till Huri, son till Jaroa, son till Gilead, son till Mikael, son till Jesisai, son till Jado, son till Bus.
Men Ahi, son till Abdiel, son till Guni, var huvudman för deras familjer.
Och de bodde i Gilead i Basan och underlydande orter, så ock på alla Sarons utmarker, så långt de sträckte sig.
Alla dessa blevo upptecknade i släktregistret i Jotams, Juda konungs, och i Jerobeams, Israels konungs, tid.
Rubens barn och gaditerna och ena hälften av Manasse stam, de av dem, som voro krigsdugliga och buro sköld och svärd och spände båge och voro stridskunniga, utgjorde fyrtiofyra tusen sju hundra sextio stridbara män.
Och de förde krig mot hagariterna och mot Jetur, Nafis och Nodab.
Och seger beskärdes dem i striden mot dessa, så att hagariterna och alla som voro med dem blevo givna i deras hand; ty de ropade till Gud under striden, och han bönhörde dem, därför att de förtröstade på honom.
Och såsom byte förde de bort deras boskapshjordar, femtio tusen kameler, två hundra femtio tusen får och två tusen åsnor, så ock ett hundra tusen människor.
Ty många hade fallit slagna, eftersom striden var av Gud.
Sedan bosatte de sig i deras land och bodde där ända till fångenskapen.
Halva Manasse stams barn bodde ock där i landet, från Basan ända till Baal-Hermon och Senir och Hermons berg, och de voro talrika.
Och dessa voro huvudmän för sina familjer: Efer, Jisei, Eliel, Asriel, Jeremia, Hodauja och Jadiel, tappra stridsmän, namnkunniga män, huvudmän för sina familjer.
Men de blevo otrogna mot sina fäders Gud, i det att de i trolös avfällighet lupo efter de gudar som dyrkades av de folk där i landet, som Gud hade förgjort för dem.
Då uppväckte Israels Gud den assyriske konungen Puls ande och den assyriske konungen Tillegat-Pilnesers ande och lät folket föras bort i fångenskap, såväl rubeniterna och gaditerna som ena hälften av Manasse stam, och lät dem komma till Hala, Habor, Hara och Gosans ström, där de äro ännu i dag.
Levis söner voro Gerson, Kehat och Merari.
Kehats söner voro Amram, Jishar, Hebron och Ussiel.
Amrams barn voro Aron, Mose och Mirjam.
Arons söner voro Nadab och Abihu, Eleasar och Itamar.
Eleasar födde Pinehas, Pinehas födde Abisua.
Abisua födde Bucki, och Bucki födde Ussi.
Ussi födde Seraja, och Seraja födde Merajot.
Merajot födde Amarja, och Amarja födde Ahitub.
Ahitub födde Sadok, och Sadok födde Ahimaas.
Ahimaas födde Asarja, och Asarja födde Johanan.
Johanan födde Asarja; det var han som var präst i det tempel som Salomo byggde i Jerusalem.
Asarja födde Amarja, och Amarja födde Ahitub.
Ahitub födde Sadok, och Sadok födde Sallum.
Sallum födde Hilkia, och Hilkia födde Asarja.
Asarja födde Seraja, och Seraja födde Josadak.
Men Josadak måste gå med i fångenskap, när HERREN lät Juda och Jerusalem föras bort genom Nebukadnessar.
Levis söner voro Gersom, Kehat och Merari.
Och dessa voro namnen på Gersoms söner: Libni och Simei.
Och Kehats söner voro Amram, Jishar, Hebron och Ussiel.
Meraris söner voro Maheli och Musi.
Dessa voro leviternas släkter, efter deras fäder.
Från Gersom härstammade hans son Libni, dennes son Jahat, dennes son Simma,
dennes son Joa, dennes son Iddo, dennes son Sera, dennes son Jeaterai.
Kehats söner voro hans son Amminadab, dennes son Kora, dennes son Assir,
dennes son Elkana, dennes son Ebjasaf, dennes son Assir,
dennes son Tahat, dennes son Uriel, dennes son Ussia och dennes son Saul.
Elkanas söner voro Amasai och Ahimot.
Hans son var Elkana; hans son var Elkana-Sofai; hans son var Nahat.
Hans son var Eliab; hans son var Jeroham; hans son var Elkana.
Och Samuels söner voro Vasni, den förstfödde, och Abia.
Meraris söner voro Maheli, dennes son Libni, dennes son Simei, dennes son Ussa,
dennes son Simea, dennes son Haggia, dennes son Asaja.
Och dessa voro de som David anställde för att ombesörja sången i HERRENS hus, sedan arken hade fått en vilostad.
De gjorde tjänst inför uppenbarelsetältets tabernakel såsom sångare, till dess att Salomo byggde HERRENS hus i Jerusalem; de stodo där och förrättade sin tjänst, såsom det var föreskrivet för dem.
Dessa voro de som så tjänstgjorde, och dessa voro deras söner: Av kehatiternas barn: Heman, sångaren, son till Joel, son till Samuel,
son till Elkana, son till Jeroham, son till Eliel, son till Toa,
son till Sif, son till Elkana, son till Mahat, son till Amasai,
son till Elkana, son till Joel, son till Asarja, son till Sefanja,
son till Tahat, son till Assir, son till Ebjasaf, son till Kora,
son till Jishar, son till Kehat, son till Levi, son till Israel;
vidare hans broder Asaf, som hade sin plats på hans högra sida, Asaf, son till Berekja, son till Simea,
son till Mikael, son till Baaseja, son till Malkia,
son till Etni, son till Sera, son till Adaja,
son till Etan, son till Simma, son till Simei,
son till Jahat, son till Gersom, son till Levi.
Och deras bröder, Meraris barn stodo på den vänstra sidan: Etan son till Kisi, son till Abdi, son till Malluk,
son till Hasabja, son till Amasja, son till Hilkia,
son till Amsi, son till Bani, son till Semer,
son till Maheli, son till Musi, son till Merari, son till Levi.
Och deras bröder, de övriga leviterna, hade blivit givna till allt slags tjänstgöring vid tabernaklet, Guds hus.
Men Aron och hans söner ombesörjde offren på brännoffersaltaret och på rökelsealtaret, och skulle utföra all förrättning i det allraheligaste och bringa försoning för Israel, alldeles såsom Mose, Guds tjänare, hade bjudit.
Och dessa voro Arons söner: hans son Eleasar, dennes son Pinehas, dennes son Abisua,
dennes son Bucki, dennes son Ussi, dennes son Seraja,
dennes son Merajot, dennes son Amarja, dennes son Ahitub,
dennes son Sadok, dennes son Ahimaas.
Och dessa voro deras boningsorter, efter deras tältläger inom deras område: Åt Arons söner av kehatiternas släkt -- ty dem träffade nu lotten --
åt dem gav man Hebron i Juda land med dess utmarker runt omkring.
Men åkerjorden och byarna som hörde till staden gav man åt Kaleb, Jefunnes son.
Åt Arons söner gav man alltså fristäderna Hebron och Libna med dess utmarker, vidare Jattir och Estemoa med dess utmarker.
Hilen med dess utmarker, Debir med dess utmarker,
Asan med dess utmarker och Bet-Semes med dess utmarker;
och ur Benjamins stam Geba med dess utmarker, Alemet med dess utmarker och Anatot med dess utmarker, så att deras städer tillsammans utgjorde tretton städer, efter deras släkter.
Och Kehats övriga barn fingo ur en stamsläkt, nämligen den stamhalva som utgjorde ena hälften av Manasse stam, genom lottkastning tio städer.
Gersoms barn åter fingo, efter sina släkter, ur Isaskars stam, ur Asers stam, ur Naftali stam och ur Manasse stam i Basan tretton städer.
Meraris barn fingo, efter sina släkter, ur Rubens stam, ur Gads stam och ur Sebulons stam genom lottkastning tolv städer.
Så gåvo Israels barn åt leviterna dessa städer med deras utmarker.
Genom lottkastning gåvo de åt dem ur Juda barns stam, ur Simeons barns stam och ur Benjamins barns stam dessa städer, som de namngåvo.
Och bland Kehats barns släkter fingo några följande städer ur Efraims stam såsom sitt område:
Man gav dem fristäderna Sikem med dess utmarker i Efraims bergsbygd, Geser med dess utmarker,
Jokmeam med dess utmarker, Bet-Horon med dess utmarker;
vidare Ajalon med dess utmarker och Gat-Rimmon med dess utmarker;
och ur ena hälften av Manasse stam Aner med dess utmarker och Bileam med dess utmarker.
Detta tillföll Kehats övriga barns släkt.
Gersoms barn fingo ur den släkt som utgjorde ena hälften av Manasse stam Golan i Basan med dess utmarker och Astarot med dess utmarker;
och ur Isaskars stam Kedes med dess utmarker, Dobrat med dess utmarker,
Ramot med dess utmarker och Anem med dess utmarker;
och ur Asers stam Masal med dess utmarker, Abdon med dess utmarker,
Hukok med dess utmarker och Rehob med dess utmarker;
och ur Naftali stam Kedes i Galileen med dess utmarker, Hammon med dess utmarker och Kirjataim med dess utmarker.
Meraris övriga barn fingo ur Sebulons stam Rimmono med dess utmarker och Tabor med dess utmarker,
och på andra sidan Jordan mitt emot Jeriko, öster om Jordan, ur Rubens stam Beser i öknen med dess utmarker, Jahas med dess utmarker,
Kedemot med dess utmarker och Mefaat med dess utmarker;
och ur Gads stam Ramot i Gilead med dess utmarker, Mahanaim med dess utmarker,
Hesbon med dess utmarker och Jaeser med dess utmarker.
Och Isaskars söner voro Tola och Pua, Jasib och Simron, tillsammans fyra.
Tolas söner voro Ussi, Refaja, Jeriel, Jamai, Jibsam och Samuel, huvudmän för sina familjer, ättlingar av Tola, tappra stridsmän, upptecknade efter sin ättföljd.
I Davids tid var deras antal tjugutvå tusen sex hundra.
Ussis söner voro Jisraja, och Jisrajas söner voro Mikael, Obadja och Joel samt Jissia, tillhopa fem, allasammans huvudmän.
Och med dem följde stridbara härskaror, trettiosex tusen man, efter sin ättföljd och sina familjer; ty de hade många hustrur och barn.
Och deras bröder i alla Isaskars släkter voro tappra stridsmän; åttiosju tusen utgjorde tillsammans de som voro upptecknade i deras släktregister.
Benjamins söner voro Bela, Beker och Jediael, tillsammans tre.
Belas söner voro Esbon, Ussi, Ussiel, Jerimot och Iri, tillsammans fem, huvudmän för sina familjer, tappra stridsmän; de som voro upptecknade i deras släktregister utgjorde tjugutvå tusen trettiofyra.
Bekers söner voro Semira, Joas, Elieser, Eljoenai, Omri, Jeremot, Abia, Anatot och Alemet.
Alla dessa voro Bekers söner.
De som voro upptecknade i deras släktregister, efter sin ättföljd, efter huvudmannen för sina familjer, tappra stridsmän, utgjorde tjugu tusen två hundra.
Jediaels söner voro Bilhan; Bilhans söner voro Jeus, Benjamin, Ehud, Kenaana, Setan, Tarsis och Ahisahar.
Alla dessa voro Jediaels söner, upptecknade efter huvudmännen för sina familjer, tappra stridsmän, sjutton tusen två hundra stridbara krigsmän.
Och Suppim och Huppim voro Irs söner. -- Men Husim voro Ahers söner.
Naftalis söner voro Jahasiel, Guni, Jeser och Sallum, Bilhas söner.
Manasses söner voro Asriel, som kvinnan födde; hans arameiska bihustru födde Makir, Gileads fader.
Och Makir tog hustru åt Huppim och Suppim.
Hans syster hette Maaka.
Och den andre hette Selofhad.
Och Selofhad hade döttrar.
Och Maaka, Makirs hustru, födde en son och gav honom namnet Peres, men hans broder hette Seres.
Hans söner voro Ulam och Rekem.
Ulams söner voro Bedan.
Dessa voro söner till Gilead, son till Makir, son till Manasse.
Och hans syster var Hammoleket; hon födde Is-Hod, Abieser och Mahela.
Och Semidas söner voro Ajan, Sekem, Likhi och Aniam.
Och Efraims söner voro Sutela, dennes son Bered, dennes son Tahat, dennes son Eleada, dennes son Tahat,
dennes son Sabad och dennes son Sutela, så ock Eser och Elead.
Och män från Gat, som voro födda där i landet, dräpte dem, därför att de hade dragit ned för att taga deras boskapshjordar.
Då sörjde Efraim, deras fader, i lång tid, och hans bröder kommo för att trösta honom.
Och han gick in till sin hustru, och hon blev havande och födde en son; och han gav honom namnet Beria , därför att det hade skett under en olyckstid för hans hus.
Hans dotter var Seera; hon byggde Nedre och Övre Bet-Horon, så ock Ussen-Seera.
Och hans son var Refa; hans son var Resef, ävensom Tela; hans son var Tahan.
Hans son var Laedan; hans son var Ammihud; hans son var Elisama.
Hans son var Non; hans son var Josua.
Och deras besittning och deras boningsorter voro Betel med underlydande orter, österut Naaran och västerut Geser med underlydande orter, vidare Sikem med underlydande orter, ända till Aja med underlydande orter.
Men i Manasse barns ägo voro Bet-Sean med underlydande orter, Taanak med underlydande orter, Megiddo med underlydande orter, Dor med underlydande orter.
Här bodde nu Josefs, Israels sons, barn.
Asers söner voro Jimna, Jisva, Jisvi och Beria; och deras syster var Sera.
Berias söner voro Heber och Malkiel; han var Birsaits fader.
Och Heber födde Jaflet, Somer och Hotam, så ock Sua, deras syster.
Och Jaflets söner voro Pasak, Bimhal och Asvat.
Dessa voro Jaflets söner.
Semers söner voro Ahi och Rohaga, Jaba och Aram.
Hans broder Helems söner voro Sofa, Jimna, Seles och Amal.
Sofas söner voro Sua, Harnefer, Sual, Beri och Jimra,
Beser, Hod, Samma, Silsa, Jitran och Beera.
Jeters söner voro Jefunne, Pispa och Ara.
Och Ullas söner voro Ara, Hanniel och Risja.
Alla dessa voro Asers söner, huvudmän för sina familjer, utvalda tappra stridsmän, huvudmän bland hövdingarna; och de som voro upptecknade i deras släktregister såsom dugliga till krigstjänst utgjorde ett antal av tjugusex tusen man.
Och Benjamin födde Bela, sin förstfödde, Asbel, den andre, och Ahara, den tredje,
Noha, den fjärde, och Rafa, den femte.
Bela hade följande söner: Addar, Gera, Abihud,
Abisua, Naaman, Ahoa,
Gera, Sefufan och Huram.
Och dessa voro Ehuds söner, och de voro familjehuvudmän för dem som bodde i Geba, och som blevo bortförda till Manahat,
dit Gera jämte Naaman och Ahia förde bort dem: han födde Ussa och Ahihud.
Och Saharaim födde barn i Moabs land, sedan han hade skilt sig från sina hustrur, Husim och Baara;
med sin hustru Hodes födde han där Jobab, Sibja, Mesa, Malkam,
Jeus, Sakeja och Mirma.
Dessa voro hans söner, huvudmän för familjer.
Med Husim hade han fött Abitub och Elpaal.
Och Elpaals söner voro Eber, Miseam och Semed.
Han var den som byggde Ono och Lod med underlydande orter.
Beria och Sema -- vilka voro familjehuvudmän för Ajalons invånare och förjagade Gats invånare --
så ock Ajo, Sasak och Jeremot.
Och Sebadja, Arad, Eder,
Mikael, Jispa och Joha voro Berias söner.
Och Sebadja, Mesullam, Hiski, Heber,
Jismerai, Jislia och Jobab voro Elpaals söner.
Och Jakim, Sikri, Sabdi,
Elienai, Silletai, Eliel,
Adaja, Beraja och Simrat voro Simeis söner.
Och Jispan, Eber, Eliel,
Abdon, Sikri, Hanan,
Hananja, Elam, Antotja,
Jifdeja och Peniel voro Sasaks söner.
Och Samserai, Seharja, Atalja,
Jaaresja, Elia och Sikri voro Jerohams söner.
Dessa vore huvudman för familjer, huvudmän efter sin ättföljd; de bodde i Jerusalem.
I Gibeon bodde Gibeons fader, vilkens hustru hette Maaka.
Och hans förstfödde son var Abdon; vidare Sur, Kis, Baal, Nadab,
Gedor, Ajo och Seker.
Men Miklot födde Simea.
Också dessa bodde jämte sina bröder i Jerusalem, gent emot sina bröder.
Och Ner födde Kis, Kis födde Saul, och Saul födde Jonatan, Malki-Sua, Abinadab och Esbaal.
Jonatans son var Merib-Baal, och Merib-Baal födde Mika.
Mikas söner voro Piton, Melek, Taarea och Ahas.
Ahas födde Joadda, Joadda födde Alemet, Asmavet och Simri, och Simri födde Mosa.
Mosa födde Binea.
Hans son var Rafa; hans son var Eleasa; hans son var Asel.
Och Asel hade sex söner, och dessa hette Asrikam, Bokeru, Ismael, Searja, Obadja och Hanan.
Alla dessa voro Asels söner.
Och hans broder Eseks söner voro Ulam, hans förstfödde, Jeus, den andre, och Elifelet, den tredje.
Och Ulams söner voro tappra stridsmän, som voro skickliga i att spänna båge; och de hade många söner och sonsöner: ett hundra femtio.
Alla dessa voro av Benjamins barn
Och hela Israel blev upptecknat i släktregister, och de finnas uppskrivna i boken om Israels konungar.
Och Juda fördes i fångenskap bort till Babel för sin otrohets skull.
Men de förra invånarna som bodde där de hade sin arvsbesittning, i sina städer, utgjordes av vanliga israeliter, präster, leviter och tempelträlar.
I Jerusalem bodde en del av Juda barn, av Benjamins barn och av Efraims och Manasse barn, nämligen:
Utai, son till Ammihud, son till Omri, son till Imri, son till Bani, av Peres', Judas sons, barn;
av siloniterna Asaja, den förstfödde, och hans söner;
av Seras barn Jeguel och deras broder, sex hundra nittio;
av Benjamins barn Sallu, son till Mesullam, son till Hodauja, son till Hassenua,
vidare Jibneja, Jerohams son, och Ela, son till Ussi, son till Mikri, och Mesullam, son till Sefatja, son till Reguel, son till Jibneja,
så ock deras bröder, efter deras ättföljd, nio hundra femtiosex.
Alla dessa män voro huvudmän för familjer, var och en för sin familj.
Och av prästerna: Jedaja, Jojarib och Jakin,
vidare Asarja, son till Hilkia, son till Mesullam, son till Sadok, son till Merajot, son till Ahitub, fursten i Guds hus,
vidare Adaja, son till Jeroham, son till Pashur, son till Malkia, vidare Maasai, son till Adiel, son till Jasera, son till Mesullam, son till Mesillemit, son till Immer,
så ock deras bröder, huvudmän för sina familjer, ett tusen sju hundra sextio, dugande män i de sysslor som hörde till tjänstgöringen i Guds hus.
Och av leviterna: Semaja, som till Hassub, son till Asrikam, son till Hasabja, av Meraris barn,
vidare Bakbackar, Heres och Galal, så ock Mattanja, son till Mika, son till Sikri, son till Asaf,
vidare Obadja, son till Semaja, son till Galal, son till Jedutun, så ock Berekja, son till Asa, son till Elkana, som bodde i netofatiternas byar.
Och dörrvaktarna: Sallum, Ackub, Talmon och Ahiman med sina bröder; men Sallum var huvudmannen.
Och ända till nu göra de tjänst vid Konungsporten, på östra sidan.
Dessa voro dörrvaktarna i Levi barns läger.
Men Sallum, son till Kore, son till Ebjasaf, son till Kora, hade jämte sina bröder, dem som voro av hans familj, koraiterna, till tjänstgöringssyssla att hålla vakt vid tältets trösklar; deras fäder hade nämligen i HERRENS läger hållit vakt vid ingången.
Och Pinehas, Eleasars son, hade förut varit furste över dem -- med honom vare HERREN!
Sakarja, Meselemjas son, var dörrvaktare vid ingången till uppenbarelsetältet.
Alla dessa voro utvalda till dörrvaktare vid trösklarna: två hundra tolv.
De blevo i sina byar upptecknade i släktregistret.
David och siaren Samuel hade tillsatt dem att tjäna på heder och tro.
De och deras söner stodo därför vid portarna till HERRENS hus, tälthuset, och höllo vakt.
Efter de fyra väderstrecken hade dörrvaktarna sina platser: i öster, väster, norr och söder.
Och deras bröder, de som fingo bo i sina byar, skulle var sjunde dag, alltid på samma timme, infinna sig hos dem.
Ty på heder och tro voro dessa fyra anställda såsom förmän för dörrvaktarna.
Detta var nu leviterna.
De hade ock uppsikten över kamrarna och förvaringsrummen i Guds hus.
Och de vistades om natten runt omkring Guds hus, ty dem ålåg att hålla vakt, och de skulle öppna dörrarna var morgon.
Somliga av dem hade uppsikten över de kärl som användes vid tjänstgöringen.
De buro nämligen in dem, efter att hava räknat dem, och buro sedan ut dem, efter att åter hava räknat dem.
Och somliga av dem voro förordnade till att hava uppsikten över de andra kärlen, över alla andra helgedomens kärl, så ock över det fina mjölet och vinet och oljan och rökelsen och de välluktande kryddorna.
Men somliga av prästernas söner beredde salvan av de välluktande kryddorna.
Och Mattitja, en av leviterna, koraiten Sallums förstfödde, hade på heder och tro uppsikten över bakverket.
Och somliga av deras bröder, kehatiternas söner, hade uppsikten över skådebröden och skulle tillreda dem för var sabbat.
Men de andra, nämligen sångarna, huvudmän för levitiska familjer, vistades i kamrarna, fria ifrån annan tjänstgöring, ty dag och natt voro de upptagna av sina egna sysslor.
Dessa voro huvudmännen för de levitiska familjerna, huvudman efter sin ättföljd; de bodde i Jerusalem.
I Gibeon bodde Gibeons fader Jeguel, vilkens hustru hette Maaka.
Och hans förstfödde son var Abdon; vidare Sur, Kis, Baal, Ner, Nadab
Gedor, Ajo, Sakarja och Miklot.
Men Miklot födde Simeam.
Också de bodde jämte sina bröder i Jerusalem, gent emot sina bröder.
Och Ner födde Kis, Kis födde Saul, och Saul födde Jonatan, Malki-Sua, Abinadab och Esbaal.
Jonatans son var Merib-Baal, och Merib-Baal födde Mika.
Mikas söner voro Piton, Melek och Taharea.
Ahas födde Jaera, Jaera födde Alemet, Asmavet och Simri, och Simri födde Mosa.
Mosa födde Binea.
Hans son var Refaja; hans son var Eleasa; hans son var Asel.
Och Asel hade sex söner, och dessa hette Asrikam, Bokeru, Ismael, Searja, Obadja och Hanan.
Dessa voro Asels söner
Och filistéerna stridde mot Israel; och Israels män flydde för filistéerna och föllo slagna på berget Gilboa.
Och filistéerna ansatte ivrigt Saul och hans söner.
Och filistéerna dödade Jonatan, Abinadab och Malki-Sua, Sauls söner.
När då Saul själv blev häftigt anfallen och bågskyttarna kommo över honom, greps han av förskräckelse för skyttarna.
Och Saul sade till sin vapendragare: »Drag ut ditt svärd och genomborra mig därmed, så att icke dessa oomskurna komma och hantera mig skändligt.»
Men hans vapendragare ville det icke, ty han fruktade storligen.
Då tog Saul själv svärdet och störtade sig därpå.
Men när vapendragaren såg att Saul var död, störtade han sig ock på sitt svärd och dog.
Så dogo då Saul och hans tre söner; och alla som hörde till hans hus dogo på samma gång.
Och när alla israeliterna i dalen förnummo att deras här hade flytt, och att Saul och hans söner voro döda, övergåvo de sina städer och flydde; sedan kommo filistéerna och bosatte sig i dem.
Dagen därefter kommo filistéerna för att plundra de slagna och funno då Saul och hans söner, där de lågo fallna på berget Gilboa.
Och de plundrade honom och togo med sig hans huvud och hans vapen och sände dem omkring i filistéernas land och läto förkunna det glada budskapet för sina avgudar och för folket.
Och de lade hans vapen i sitt gudahus, men hans huvudskål hängde de upp i Dagons tempel.
Men när allt folket i Jabes i Gilead hörde allt vad filistéerna hade gjort med Saul,
stodo de upp, alla stridbara män, och togo Sauls och hans söners lik och förde dem till Jabes; och de begrovo deras ben under terebinten i Jabes och fastade så i sju dagar.
Detta blev Sauls död, därför att han hade begått otrohet mot HERREN, i det att han icke hade hållit HERRENS ord, så ock därför att han hade frågat en ande och sökt svar hos en sådan.
Han hade icke sökt svar hos HERREN; därför dödade HERREN honom.
Och sedan överflyttade han konungadömet på David, Isais son.
Då församlade sig hela Israel till David i Hebron och sade: »Vi äro ju ditt kött och ben.
Redan för länge sedan, redan då Saul ännu var konung, var det du som var ledare och anförare för Israel.
Och till dig har HERREN, din Gud, sagt: Du skall vara en herde för mitt folk Israel, ja, du skall vara en furste över mitt folk Israel.»
När så alla de äldste i Israel kommo till konungen i Hebron, slöt David ett förbund med dem där i Hebron, inför HERREN; och sedan smorde de David till konung över Israel, i enlighet med HERRENS ord genom Samuel.
Och David drog med hela Israel till Jerusalem, det är Jebus; där befunno sig jebuséerna, som ännu bodde kvar i landet.
Och invånarna i Jebus sade till David: »Hitin kommer du icke.»
Men David intog likväl Sions borg, det är Davids stad
Och David sade: »Vemhelst som först slår ihjäl en jebusé, han skall bliva hövding och anförare.»
Och Joab, Serujas son, kom först ditupp och blev så hövding.
Sedan tog David sin boning i bergfästet; därför kallade man det Davids stad.
Och han uppförde befästningsverk runt omkring staden, från Millo och allt omkring; och Joab återställde det övriga av staden.
Och David blev allt mäktigare och mäktigare, och HERREN Sebaot var med honom
Och dessa äro de förnämsta bland Davids hjältar, vilka gåvo honom kraftig hjälp att bliva konung, de jämte hela Israel, och så skaffade honom konungaväldet, enligt HERRENS ord angående Israel.
Detta är förteckningen på Davids hjältar: Jasobeam, son till en hakmonit, den förnämste bland kämparna, han som svängde sitt spjut över tre hundra som hade blivit slagna på en gång.
Och efter honom kom ahoaiten Eleasar, son till Dodo; han var en av de tre hjältarna.
Han var med David vid Pas-Dammim, när filistéerna där hade församlat sig till strid.
Och där var ett åkerstycke, fullt med korn.
Och folket flydde för filistéerna.
Då ställde de sig mitt på åkerstycket och försvarade det och slogo filistéerna; och HERREN lät dem så vinna en stor seger.
En gång drogo tre av de trettio förnämsta männen ned över klippan till David vid Adullams grotta, medan en avdelning filistéer var lägrad i Refaimsdalen.
Men David var då på borgen, under det att en filisteisk utpost fanns i Bet-Lehem.
Och David greps av lystnad och sade: »Ack att någon ville giva mig vatten att dricka från brunnen vid Bet-Lehems stadsport!»
Då bröto de tre sig igenom filistéernas läger och hämtade vatten ur brunnen vid Bet-Lehems stadsport och togo det och buro det till David.
Men David ville icke dricka det, utan göt ut det såsom ett drickoffer åt HERREN.
Han sade nämligen: »Gud låte det vara fjärran ifrån mig att jag skulle göra detta!
Skulle jag dricka dessa mäns blod, som hava vågat sina liv?
Ty med fara för sina liv hava de burit det hit.»
Och han ville icke dricka det.
Sådana ting hade de tre hjältarna gjort.
Absai, Joabs broder, var den förnämste av tre andra; han svängde en gång sitt spjut över tre hundra som hade blivit slagna.
Och han hade ett stort namn bland de tre.
Han var dubbelt mer ansedd än någon annan i detta tretal, och han var deras hövitsman, men upp till de tre första kom han dock icke.
Vidare Benaja, son till Jojada, som var son till en tapper, segerrik man från Kabseel; han slog ned de två Arielerna i Moab, och det var han som en snövädersdag steg ned och slog ihjäl lejonet i brunnen.
Han slog ock ned den egyptiske mannen som var så reslig: fem alnar lång.
Fastän egyptiern i handen hade ett spjut som liknade en vävbom, gick han ned mot honom, väpnad allenast med sin stav.
Och han ryckte spjutet ur egyptiern hand och dräpte honom med hans eget spjut.
Sådana ting hade Benaja, Jojadas son, gjort.
Och han hade ett stort namn bland de tre hjältarna.
Ja, han var mer ansedd än någon av de trettio, men upp till de tre första kom han icke.
Och David satte honom till anförare för sin livvakt.
De tappra hjältarna voro: Asael, Joabs broder, Elhanan, Dodos son, från Bet-Lehem;
haroriten Sammot; peloniten Heles;
tekoaiten Ira, Ickes' son; anatotiten Abieser;
husatiten Sibbekai; ahoaiten Ilai;
netofatiten Maherai; netofatiten Heled, Baanas son;
Itai, Ribais son, från Gibea i Benjamins barns stam; pirgatoniten Benaja;
Hurai från Gaas' dalar; arabatiten Abiel;
baharumiten Asmavet; saalboniten Eljaba;
gisoniten Bene-Hasem; harariten Jonatan, Sages son;
harariten Ahiam, Sakars son; Elifal, Urs son;
mekeratiten Hefer; peloniten Ahia;
Hesro från Karmel; Naarai, Esbais son;
Joel, broder till Natan; Mibhar, Hagris son;
ammoniten Selek; berotiten Naherai, vapendragare åt Joab, Serujas son;
jeteriten Ira; jeteriten Gareb;
hetiten Uria; Sabad, Alais son;
rubeniten Adina, Sisas son, en huvudman bland rubeniterna, och jämte honom trettio andra;
Hanan, Maakas son, och mitniten Josafat;
astarotiten Ussia; Sama och Jeguel, aroeriten Hotams söner;
Jediael, Simris son, och hans broder Joha, tisiten;
Eliel-Hammahavim samt Jeribai och Josauja, Elnaams söner, och moabiten Jitma;
slutligen Eliel, Obed och Jaasiel-Hammesobaja.
Och dessa voro de som kommo till David i Siklag, medan han ännu höll sig undan för Saul, Kis' son; de hörde till de hjältar som bistodo honom under kriget.
De voro väpnade med båge och skickliga i att, både med höger och med vänster hand, slunga stenar och avskjuta pilar från bågen.
Av Sauls stamfränder, benjaminiterna, kommo:
Ahieser, den förnämste, och Joas, gibeatiten Hassemaas söner; Jesuel och Pelet, Asmavets söner; Beraka; anatotiten Jehu;
gibeoniten Jismaja, en av de trettio hjältarna, anförare för de trettio; Jeremia; Jahasiel; Johanan; gederatiten Josabad;
Eleusai; Jerimot; Bealja; Semarja; harufiten Sefatja;
koraiterna Elkana, Jissia, Asarel, Joeser och Jasobeam;
Joela och Sebadja, söner till Jeroham, av strövskaran.
Och av gaditerna avföllo några och gingo till David i bergfästet i öknen, tappra män, krigsmän skickliga att strida, rustade med sköld och spjut; de hade en uppsyn såsom lejon och voro snabba såsom gaseller på bergen:
Eser, den förnämste, Obadja, den andre, Eliab, den tredje,
Masmanna, den fjärde, Jeremia, den femte,
Attai, den sjätte, Eliel, den sjunde,
Johanan, den åttonde, Elsabad, den nionde,
Jeremia, den tionde, Makbannai, den elfte.
Dessa hörde till Gads barn och till de förnämsta i hären; den ringaste av dem var ensam så god som hundra, men den ypperste så god som tusen.
Dessa voro de som i första månaden gingo över Jordan, när den var full över alla sina bräddar, och som förjagade alla dem som bodde i dalarna, åt öster och åt väster.
Av Benjamins och Juda barn kommo några män till David ända till bergfästet.
Då gick David ut emot dem och tog till orda och sade till dem: »Om I kommen till mig i fredlig avsikt och viljen bistå mig, så är mitt hjärta redo till förening med eder; men om I kommen för att förråda mig åt mina ovänner, fastän ingen orätt är i mina händer, då må våra fäders Gud se därtill och straffa det.»
Men Amasai, den förnämste bland de trettio, hade blivit beklädd med andekraft, och han sade: »Dina äro vi, David, och med dig stå vi, du Isais son.
Frid vare med dig, frid, och frid vare med dem som bistå dig ty din Gud har bistått dig!»
Och David tog emot dem och gav dem plats bland de förnämsta i sin skara.
Från Manasse gingo några över till David, när han med filistéerna drog ut i strid mot Saul, dock fingo de icke bistå dessa; ty när filistéernas hövdingar hade rådplägat, skickade de bort honom, i det de sade: »Det gäller huvudet för oss, om han går över till sin herre Saul.
När han då drog till Siklag, gingo dessa från Manasse över till honom: Adna, Josabad, Jediael, Mikael, Josabad, Elihu och Silletai, huvudmän för de ätter som tillhörde Manasse.
Dessa bistodo David mot strövskaran, ty de voro allasammans tappra stridsmän och blevo hövitsmän i hären.
Dag efter dag kommo nämligen allt flera till David för att bistå honom, så att hans läger blev övermåttan stort.
Detta är de tal som angiva summorna av det väpnade krigsfolk som kom till David i Hebron, för att efter HERRENS befallning flytta Sauls konungamakt över på honom:
Juda barn, som buro sköld och spjut, sex tusen åtta hundra, väpnade till strid;
av Simeons barn tappra krigsmän, sju tusen ett hundra;
av Levi barn fyra tusen sex hundra;
därtill Jojada, fursten inom Arons släkt, och med honom tre tusen sju hundra;
så ock Sadok, en tapper yngling, med sin familj, tjugutvå hövitsmän;
av Benjamins barn, Sauls stamfränder, tre tusen (ty ännu vid den tiden höllo de flesta av dem troget med Sauls hus);
av Efraims barn tjugu tusen åtta hundra, tappra stridsmän, namnkunniga män i sina familjer;
av ena hälften av Manasse stam aderton tusen namngivna män, som kommo för att göra David till konung;
av Isaskars barn kommo män som väl förstodo tidstecknen och insågo vad Israel borde göra, två hundra huvudmän, därtill alla deras stamfränder under deras befäl;
av Sebulon stridbara män, rustade till krig med alla slags vapen, femtio tusen, som samlades endräktigt;
av Naftali ett tusen hövitsmän, och med dem trettiosju tusen, väpnade med sköld och spjut;
av daniterna krigsrustade män, tjuguåtta tusen sex hundra;
av Aser stridbara män, rustade till krig, fyrtio tusen;
och från andra sidan Jordan, av rubeniterna, gaditerna och andra hälften av Manasse stam, ett hundra tjugu tusen, väpnade med alla slags vapen som brukas vid krigföring.
Alla dessa krigsmän, ordnade till strid, kommo i sina hjärtans hängivenhet till Hebron för att göra David till konung över hela Israel.
Också hela det övriga Israel var enigt i att göra David till konung.
Och de voro där hos David i tre dagar och åto och drucko, ty deras bröder hade försett dem med livsmedel.
De som bodde närmast dem, ända upp till Isaskar, Sebulon och Naftali, tillförde dem ock på åsnor, kameler, mulåsnor och oxar livsmedel i myckenhet till föda: mjöl, fikonkakor och russinkakor, vin och olja, fäkreatur och småboskap; ty glädje rådde i Israel.
Och David rådförde sig med över- och underhövitsmännen, med alla furstarna.
Sedan sade David till Israels hela församling: »Om I så finnen för gott, och om detta är från HERREN, vår Gud, så låt oss sända bud åt alla håll till våra övriga bröder i alla Israels landsändar, och därjämte till prästerna och leviterna i de städer kring vilka de hava sina utmarker, att de må församla sig till oss;
och låt oss flytta vår Guds ark till oss, ty i Sauls tid frågade vi icke efter den.»
Och hela församlingen svarade att man skulle göra så, ty förslaget behagade hela folket.
Så församlade då David hela Israel, från Sihor i Egypten ända dit där vägen går till Hamat, för att hämta Guds ark från Kirjat-Jearim.
Och David drog med hela Israel upp till Baala, det är Kirjat-Jearim, som hör till Juda, för att därifrån föra upp Guds, HERRENS, ark, hans som tronar på keruberna, och efter vilken den hade fått sitt namn.
Och de satte Guds ark på en ny vagn och förde den bort ifrån Abinadabs hus; och Ussa och Ajo körde vagnen.
Och David och hela Israel fröjdade sig inför Gud av all makt, med sånger och med harpor, psaltare, pukor, cymbaler och trumpeter.
Men när de kommo till Kidonslogen, räckte Ussa ut sin hand för att fatta I arken, ty oxarna snavade.
Då upptändes HERRENS vrede mot Ussa, och därför att han hade räckt ut sin hand mot arken, slog han honom, så att han föll ned död där inför Gud.
Men det gick David hårt till sinnes att HERREN så hade brutit ned Ussa ; och han kallade det stället Peres-Ussa , såsom det heter ännu i dag.
Och David betogs av sådan fruktan för Gud på den dagen, att han sade: »Huru skulle jag töras låta föra Guds ark till mig?»
Därför lät David icke flytta in arken till sig i Davids stad, utan lät sätta in den i gatiten Obed-Edoms hus.
Sedan blev Guds ark kvar vid Obed-Edoms hus, där den stod i sitt eget hus, i tre månader; men HERREN välsignade Obed-Edoms hus och allt vad som hörde honom till.
Och Hiram, konungen i Tyrus, skickade sändebud till David med cederträ, därjämte ock murare och timmermän, för att de skulle bygga honom ett hus.
Och David märkte att HERREN hade befäst honom såsom konung över Israel; ty han hade låtit hans rike bliva övermåttan upphöjt, för sitt folk Israels skull.
Och David tog sig ännu flera hustrur i Jerusalem, och David födde ännu flera söner och döttrar.
Dessa äro namnen på de söner som han fick i Jerusalem: Sammua, Sobab, Natan, Salomo,
Jibhar, Elisua, Elpelet,
Noga, Nefeg, Jafia,
Elisama, Beeljada och Elifelet.
Men när filistéerna hörde att David hade blivit smord till konung över hela Israel, drogo de allasammans upp för att fånga David.
När David hörde detta, drog han ut mot dem.
Då nu filistéerna hade fallit in i Refaimsdalen och där företogo plundringståg,
frågade David Gud: »Skall jag draga upp mot filistéerna?
Vill du då giva dem i min hand?»
HERREN svarade honom: »Drag upp; jag vill giva dem i din hand.»
Och de drogo upp till Baal-Perasim, och där slog David dem.
Då sade David: »Gud har brutit ned mina fiender genom min hand, likasom en vattenflod bryter ned.»
Därav fick det stället namnet Baal-Perasim .
De lämnade där efter sig sina gudar; och David befallde att dessa skulle brännas upp i eld.
Men filistéerna företogo ännu en gång plundringståg i dalen.
När David då åter frågade Gud, svarade Gud honom: »Du skall icke draga upp efter dem; du må kringgå dem på en omväg, så att du kommer över dem från det håll där bakaträden stå.
Så snart du sedan hör ljudet av steg i bakaträdens toppar, drag då ut till strid, ty då har Gud dragit ut framför dig till att slå filistéernas här.»
David gjorde såsom Gud hade bjudit honom; och de slogo filistéernas här och förföljde dem från Gibeon ända till Geser.
Och ryktet om David gick ut i alla länder, och HERREN lät fruktan för honom komma över alla folk.
Och han uppförde åt sig hus i Davids stad; sedan beredde han en plats åt Guds ark och slog upp ett tält åt den.
Därvid befallde David: »Inga andra än leviterna må bära Guds ark; ty dem har HERREN utvalt till att bära Guds ark och till att göra tjänst inför honom för evärdlig tid.»
Och David församlade hela Israel till Jerusalem för att hämta HERRENS ark upp till den plats som han hade berett åt den.
Och David samlade tillhopa Arons barn och leviterna;
av Kehats barn: Uriel, deras överste, och hans bröder, ett hundra tjugu;
av Meraris barn: Asaja, deras överste, och hans bröder, två hundra tjugu;
av Gersoms barn: Joel, deras överste, och hans bröder, ett hundra trettio;
av Elisafans barn: Semaja, deras överste, och hans bröder, två hundra;
av Hebrons barn: Eliel, deras överste, och hans bröder, åttio;
av Ussiels barn: Amminadab, deras överste, och hans bröder, ett hundra tolv.
Och David kallade till sig prästerna Sadok och Ebjatar jämte leviterna Uriel, Asaja, Joel, Semaja, Eliel och Amminadab.
Och han sade till dem: »I ären huvudmän för leviternas familjer.
Helgen eder tillika med edra bröder, och hämten så HERRENS, Israels Guds, ark upp till den plats som jag har berett åt den.
Ty därför att I förra gången icke voren tillstädes var det som HERREN, vår Gud, bröt ned en av oss, till straff för att vi icke sökte honom så, som tillbörligt var.»
Då helgade prästerna och leviterna sig till att hämta upp HERRENS, Israels Guds, ark.
Och såsom Mose hade bjudit i enlighet med HERRENS ord, buro nu Levi barn Guds ark med stänger, som vilade på deras axlar.
Och David sade till de översta bland leviterna att de skulle förordna sina bröder sångarna till tjänstgöring med musikinstrumenter, psaltare, harpor och cymbaler, som de skulle låta ljuda, under det att de höjde glädjesången.
Leviterna förordnade då Heman, Joels son, och av hans bröder Asaf, Berekjas son, och av dessas bröder, Meraris barn, Etan, Kusajas son,
och jämte dem deras bröder av andra ordningen Sakarja, Ben, Jaasiel, Semiramot, Jehiel, Unni, Eliab, Benaja, Maaseja, Mattitja, Elifalehu, Mikneja, Obed-Edom och Jegiel, dörrvaktarna.
Och sångarna, Heman, Asaf och Etan, skulle slå kopparcymbaler.
Sakarja, Asiel, Semiramot, Jehiel, Unni, Eliab, Maaseja och Benaja skulle spela på psaltare, till Alamót.
Mattitja, Elifalehu, Mikneja, Obed-Edom, Jegiel och Asasja skulle leda sången med harpor, till Seminit.
Kenanja, leviternas anförare, när de buro, skulle undervisa i att bära, ty han var kunnig i sådant.
Berekja och Elkana skulle vara dörrvaktare vid arken.
Sebanja, Josafat, Netanel, Amasai, Sakarja, Benaja och Elieser, prästerna, skulle blåsa i trumpeter framför Guds ark.
Slutligen skulle Obed-Edom och Jehia vara dörrvaktare vid arken.
Så gingo då David och de äldste i Israel och överhövitsmännen åstad för att hämta HERRENS förbundsark upp ur Obed-Edoms hus, under jubel.
Och då Gud skyddade leviterna som buro HERRENS förbundsark, offrade man sju tjurar och sju vädurar.
Därvid var David klädd i en kåpa av fint linne; så voro ock alla leviterna som buro arken, så ock sångarna och Kenanja, som anförde sångarna, när de buro.
Och därjämte bar David en linne-efod.
Och hela Israel hämtade upp HERRENS förbundsark under jubel och basuners ljud; och man blåste i trumpeter och slog cymbaler och lät psaltare och harpor ljuda.
När då HERRENS förbundsark kom till Davids stad, blickade Mikal, Sauls dotter, ut genom fönstret, och då hon såg konung David dansa och göra sig glad, fick hon förakt för honom i sitt hjärta.
Sedan de hade fört Guds ark ditin, ställde de den i tältet som David hade slagit upp åt den, och framburo därefter brännoffer och tackoffer inför Guds ansikte.
När David hade offrat brännoffret och tackoffret, välsignade han folket i HERRENS namn.
Och åt var och en av alla israeliterna, både man och kvinna, gav han en kaka bröd, ett stycke kött och en druvkaka.
Och han förordnade vissa leviter till att göra tjänst inför HERRENS ark, för att de skulle prisa, tacka och lova HERREN, Israels Gud:
Asaf såsom anförare, näst efter honom Sakarja, och vidare Jegiel, Semiramot, Jehiel, Mattitja, Eliab, Benaja, Obed-Edom och Jegiel med psaltare och harpor; och Asaf skulle slå cymbaler.
Men prästerna Benaja och Jahasiel skulle beständigt stå med sina trumpeter framför Guds förbundsark.
På den dagen var det som David först fastställde den ordningen att man genom Asaf och hans bröder skulle tacka HERREN på detta sätt:
»Tacken HERREN, åkallen hans namn, gören hans gärningar kunniga bland folken.
Sjungen till hans ära, lovsägen honom, talen om alla hans under.
Berömmen eder av hans heliga namn; glädje sig av hjärtat de som söka HERREN.
Frågen efter HERREN och hans makt, söken hans ansikte beständigt.
Tänken på de underbara verk som han har gjort, på hans under och hans muns domar,
I Israels, hans tjänares, säd, I Jakobs barn, hans utvalda.
Han är HERREN, vår Gud; över hela jorden gå hans domar.
Tänken evinnerligen på hans förbund, intill tusen släkten på vad han har stadgat,
på det förbund han slöt med Abraham och på hans ed till Isak.
Han fastställde det för Jakob till en stadga, för Israel till ett evigt förbund;
han sade: 'Åt dig vill jag giva Kanaans land, det skall bliva eder arvedels lott.'
Då voren I ännu en liten hop, I voren ringa och främlingar därinne.
Och de vandrade åstad ifrån folk till folk ifrån ett rike bort till ett annat.
Han tillstadde ingen att göra dem skada, han straffade konungar för deras skull:
'Kommen icke vid mina smorda, och gören ej mina profeter något ont.'
Sjungen till HERRENS ära, alla länder, båden glädje var dag, förkunnen hans frälsning.
Förtäljen bland hedningarna hans ära, bland alla folk hans under.
Ty stor är HERREN och högt lovad, och fruktansvärd är han mer än alla gudar.
Ty folkens alla gudar äro avgudar, men HERREN är den som har gjort himmelen.
Majestät och härlighet äro inför hans ansikte, makt och fröjd i hans boning.
Given åt HERREN, I folkens släkter, given åt HERREN ära och makt;
given åt HERREN hans namns ära, bären fram skänker och kommen inför hans ansikte, tillbedjen HERREN i helig skrud.
Bäven för hans ansikte, alla länder; se, jordkretsen står fast och vacklar icke.
Himmelen vare glad, och jorden fröjde sig, och bland hedningarna säge man: 'HERREN är nu konung!'
Havet bruse och allt vad däri är, marken glädje sig och allt som är därpå;
ja, då juble skogens träd inför HERREN, ty han kommer för att döma jorden.
Tacken HERREN, ty han är god, ty hans nåd varar evinnerligen,
och sägen: 'Fräls oss, du vår frälsnings Gud, församla oss och rädda oss från hedningarna, så att vi få prisa ditt heliga namn och berömma oss av ditt lov.'
Lovad vare HERREN, Israels Gud, från evighet till evighet!»
Och allt folket sade: »Amen», och lovade HERREN.
Och han gav där, inför HERRENS förbundsark, åt Asaf och hans bröder uppdraget att beständigt göra tjänst inför arken, var dag med de för den dagen bestämda sysslorna.
Men Obed-Edom och deras bröder voro sextioåtta; och Obed-Edom, Jedituns son, och Hosa gjorde han till dörrvaktare.
Och prästen Sadok och hans bröder, prästerna, anställde han inför HERRENS tabernakel, på offerhöjden i Gibeon,
för att de beständigt skulle offra åt HERREN brännoffer på brännoffersaltaret, morgon och afton, och göra allt vad som var föreskrivet i HERRENS lag, den som han hade givit åt Israel;
och jämte dem Heman och Jedutun och de övriga namngivna utvalda, på det att de skulle tacka HERREN, därför att hans nåd varar evinnerligen.
Och hos dessa, nämligen Heman och Jedutun, förvarades trumpeter och cymbaler åt dem som skulle spela, så ock andra instrumenter som hörde till gudstjänsten.
Och Jedutuns söner gjorde han till dörrvaktare.
Sedan gick allt folket hem, var och en till sitt; men David vände om för att hälsa sitt husfolk.
Då nu David satt i sitt hus, sade han till profeten Natan: »Se, jag bor i ett hus av cederträ, under det att HERRENS förbundsark står under ett tält.»
Natan sade till David: »Gör allt vad du har i sinnet; ty Gud är med dig.»
Men om natten kom Guds ord till Natan; han sade:
»Gå och säg till min tjänare David: Så säger HERREN: Icke du skall bygga mig det hus som jag skall bo i.
Jag har ju icke bott i något hus, från den dag då jag förde Israel hitupp ända till denna dag, utan jag har flyttat ifrån tält till tält, ifrån tabernakel till tabernakel.
Har jag då någonsin, varhelst jag flyttade omkring med hela Israel, talat och sagt så till någon enda av Israels domare, som jag har förordnat till herde för mitt folk: 'Varför haven I icke byggt mig ett hus av cederträ?'
Och nu skall du säga så till min tjänare David: Så säger HERREN Sebaot: Från betesmarken, där du följde fåren, har jag hämtat dig, för att du skulle bliva en furste över mitt folk Israel.
Och jag har varit med dig på alla dina vägar och utrotat alla dina fiender för dig.
Och jag vill göra dig ett namn, sådant som de störstes namn på jorden.
Jag skall bereda en plats åt mitt folk Israel och plantera det, så att det får bo kvar där, utan att vidare bliva oroat.
Orättfärdiga människor skola icke mer föröda det, såsom fordom skedde,
och såsom det har varit allt ifrån den tid då jag förordnade domare över mitt folk Israel; och jag skall kuva alla dina fiender.
Så förkunnar jag nu för dig att HERREN skall bygga ett hus åt dig.
Ty det skall ske, att när din tid är ute och du går till dina fäder skall jag efter dig upphöja din son, en av dina avkomlingar; och jag skall befästa hans konungamakt.
Han skall bygga ett hus åt mig, och jag skall befästa hans tron för evig tid.
Jag skall vara hans fader, och han skall vara min son; och min nåd skall jag icke låta vika ifrån honom, såsom jag lät den vika ifrån din företrädare.
Jag skall hålla honom vid makt i mitt hus och i mitt rike för evig tid, och hans tron skall vara befäst för evig tid.»
Alldeles i överensstämmelse med dessa ord och med denna syn talade nu Natan till David.
Då gick konung David in och satte sig ned inför HERRENS ansikte och sade: »Vem är jag, HERRE Gud, och vad är mitt hus, eftersom du har låtit mig komma härtill?
Och detta har likväl synts dig vara för litet, o Gud; du har talat angående din tjänares hus om det som ligger långt fram i tiden.
Ja, du har sett till mig på människosätt, for att upphöja mig, HERRE Gud.
Vad skall nu David vidare säga till dig om den ära du har bevisat din tjänare?
Du känner ju din tjänare.
HERRE, för din tjänares skull och efter ditt hjärta har du gjort allt detta stora och förkunnat alla dessa stora ting.
HERRE, ingen är dig lik, och ingen Gud finnes utom dig, efter allt vad vi hava hört med våra öron.
Och var finnes på jorden något enda folk som är likt ditt folk Israel, vilket Gud själv har gått åstad att förlossa åt sig till ett folk -- för att så göra dig ett stort och fruktansvärt namn, i det att du förjagade hedningarna för ditt folk, det som du hade förlossat ifrån Egypten?
Och du har gjort ditt folk Israel till ett folk åt dig för evig tid, och du, HERRE, har blivit deras Gud
Så må nu, HERRE, vad du har talat om din tjänare och om hans hus bliva fast för evig tid; gör såsom du har talat.
Då skall ditt namn anses fast och bliva stort till evig tid, så att man skall säga: 'HERREN Sebaot, Israels Gud, är Gud över Israel.'
Och så skall din tjänare Davids hus bestå inför dig.
Ty du, min Gud, har uppenbarat för din tjänare att du skall bygga honom ett hus; därför har din tjänare dristat att bedja inför dig.
Och nu, HERRE, du är Gud; och då du har lovat din tjänare detta goda,
så må du nu ock värdigas välsigna din tjänares hus, så att det förbliver evinnerligen inför dig.
Ty vad du, HERRE, välsignar, det är välsignat evinnerligen.»
En tid härefter slog David filistéerna och kuvade dem.
Därvid tog han Gat med underlydande orter ur filistéernas hand.
Han slog ock moabiterna; så blevo moabiterna David underdåniga och förde till honom skänker.
Likaledes slog David Hadareser, konungen i Soba, vid Hamat, när denne hade dragit åstad för att befästa sitt välde vid floden Frat.
Och David tog ifrån honom ett tusen vagnar och tog till fånga sju tusen ryttare och tjugu tusen man fotfolk; och David lät avskära fotsenorna på alla vagnshästarna, utom på ett hundra hästar, som han skonade.
När sedan araméerna från Damaskus kommo för att hjälpa Hadareser, konungen i Soba, nedgjorde David tjugutvå tusen man av dem.
Och David insatte fogdar bland araméerna i Damaskus; och araméerna blevo David underdåniga och förde till honom skänker.
Så gav HERREN seger åt David, varhelst han drog fram.
Och David tog de gyllene sköldar som Hadaresers tjänare hade burit och förde dem till Jerusalem.
Och från Hadaresers städer Tibhat och Kun tog David koppar i stor myckenhet; därav gjorde sedan Salomo kopparhavet, pelarna och kopparkärlen.
Då nu Tou, konungen i Hamat, hörde att David hade slagit Hadaresers, konungens i Soba, hela här,
sände han sin son Hadoram till konung David för att hälsa honom och lyckönska honom, därför att han hade givit sig i strid med Hadareser och slagit honom; ty Hadareser hade varit Tous fiende.
Han sände ock alla slags kärl av guld, silver och koppar.
Också dessa helgade konung David åt HERREN, likasom han hade gjort med det silver och guld han hade hemfört från alla andra folk: från edoméerna, moabiterna, Ammons barn, filistéerna och amalekiterna.
Och sedan Absai, Serujas son, hade slagit edoméerna i Saltdalen, aderton tusen man,
insatte han fogdar i Edom; och alla edoméer blevo David underdåniga.
Så gav HERREN seger åt David, varhelst han drog fram.
David regerade nu över hela Israel; och han skipade lag och rätt åt allt sitt folk.
Joab, Serujas son, hade befälet över krigshären, och Josafat, Ahiluds son, var kansler.
Sadok, Ahitubs son, och Abimelek, Ebjatars son, voro präster, och Sausa var sekreterare.
Benaja, Jojadas son, hade befälet över keretéerna och peletéerna; men Davids söner voro de förnämste vid konungens sida.
En tid härefter dog Nahas, Ammons barns konung, och hans son blev konung efter honom.
Då sade David: »Jag vill bevisa Hanun, Nahas' son, vänskap, eftersom hans fader bevisade mig vänskap.»
Och David skickade sändebud för att trösta honom i hans sorg efter fadern.
När så Davids tjänare kommo till Ammons barns land, till Hanun, för att trösta honom,
sade Ammons barns furstar till Hanun: »Menar du att David därmed att han sänder tröstare till dig vill visa dig att han ärar din fader?
Nej, för att undersöka och fördärva och bespeja landet hava hans tjänare kommit till dig.»
Då tog Hanun Davids tjänare och lät raka dem och skära av deras kläder mitt på, ända uppe vid sätet, och lät dem så gå.
Och man kom och berättade för David vad som hade hänt männen; då sände han bud emot dem, ty männen voro ju mycket vanärade.
Och konungen lät säga: »Stannen i Jeriko, till dess edert skägg hinner växa ut, och kommen så tillbaka.»
Då nu Ammons barn insågo att de hade gjort sig förhatliga för David, sände Hanun och Ammons barn ett tusen talenter silver för att leja sig vagnar och ryttare från Aram-Naharaim, från Aram-Maaka och från Soba.
De lejde sig trettiotvå tusen vagnar, ävensom hjälp av konungen i Maaka med hans folk; dessa kommo och lägrade sig framför Medeba.
Ammons barn församlade sig ock från sina städer och kommo för att strida.
När David hörde detta, sände han åstad Joab med hela hären, de tappraste krigarna.
Och Ammons barn drogo ut och ställde upp sig till strid vid ingången till staden; men de konungar som hade kommit dit ställde upp sig för sig själva på fältet.
Då Joab nu såg att han hade fiender både framför sig och bakom sig, gjorde han ett urval bland allt Israels utvalda manskap och ställde sedan upp sig mot araméerna.
Men det övriga folket överlämnade han åt sin broder Absai, och dessa fingo ställa upp sig mot Ammons barn.
Och han sade: »Om araméerna bliva mig övermäktiga, så skall du komma mig till hjälp; och om Ammons barn bliva dig övermäktiga, så vill jag hjälpa dig.
Var nu vid gott mod; ja, låt oss visa mod i striden för vårt folk och för vår Guds städer.
Sedan må HERREN göra vad honom täckes.
Därefter ryckte Joab fram med sitt folk till strid mot araméerna, och de flydde för honom.
Men när Ammons barn sågo att araméerna flydde, flydde också de för hans broder Absai och begåvo sig in i staden.
Då begav sig Joab till Jerusalem.
Då alltså araméerna sågo att de hade blivit slagna av Israel, sände de bud att de araméer som bodde på andra sidan floden skulle rycka ut, anförda av Sofak, Hadaresers härhövitsman.
När detta blev berättat för David, församlade han hela Israel och gick över Jordan, och då han kom fram till dem, ställde han upp sig i slagordning mot dem; och när David hade ställt upp sig till strid mot araméerna, gåvo dessa sig i strid med honom.
Men araméerna flydde undan för Israel, och David dräpte av araméerna manskapet på sju tusen vagnar, så ock fyrtio tusen man fotfolk; härhövitsmannen Sofak dödade han ock.
Då, alltså Hadaresers tjänare sågo att de hade blivit slagna av israeliterna, ingingo de fred med David och blevo honom underdåniga.
Efter detta ville araméerna icke vidare hjälpa Ammons barn.
Följande år, vid den tid då konungarna plägade draga i fält, tågade Joab ut med krigshären och härjade Ammons barns land, och kom så och belägrade Rabba, medan David stannade kvar i Jerusalem.
Och Joab intog Rabba och förstörde det.
Och David tog deras konungs krona från hans huvud, den befanns väga en talent guld och var prydd med en dyrbar sten.
Den sattes nu på Davids huvud.
Och han förde ut byte från staden i stor myckenhet.
Och folket därinne förde han ut och söndersargade dem med sågar och tröskvagnar av järn och med bilor.
Så gjorde David mot Ammons barns alla städer.
Sedan vände David med allt folket tillbaka till Jerusalem.
Därefter uppstod en strid med filistéerna vid Geser; husatiten Sibbekai slog då ned Sippai, en av rafaéernas avkomlingar; så blevo de kuvade.
Åter stod en strid med filistéerna; Elhanan, Jaurs son, slog då ned Lami, gatiten Goljats broder, som hade ett spjut vars skaft liknade en vävbom.
Åter stod en strid vid Gat.
Där var en reslig man som hade sex fingrar och sex tår, tillsammans tjugufyra; han var ock en avkomling av rafaéerna.
Denne smädade Israel; då blev han nedgjord av Jonatan, son till Simea, Davids broder.
Dessa voro avkomlingar av rafaéerna i Gat; och de föllo för Davids och hans tjänares hand.
Men Satan trädde upp mot Israel och uppeggade David till att räkna Israel.
Då sade David till Joab och till folkets andra hövitsman: »Gån åstad och räknen Israel, från Beer-Seba ända till Dan, och given mig besked därom, så att jag får veta huru många de äro.»
Joab svarade: »Må HERREN än vidare föröka sitt folk hundrafalt.
Äro de då icke, min herre konung, allasammans min herres tjänare?
Varför begär då min herre sådant?
Varför skulle man därmed draga skuld över Israel?
Likväl blev konungens befallning gällande, trots Joab.
Alltså drog Joab ut och for omkring i hela Israel, och kom så hem igen till Jerusalem.
Och Joab uppgav för David vilken slutsumma folkräkningen utvisade: i Israel funnos tillsammans elva hundra tusen svärdbeväpnade män, och i Juda funnos fyra hundra sjuttio tusen svärdbeväpnade man.
Men Levi och Benjamin hade han icke räknat jämte de andra, ty konungens befallning var en styggelse för Joab.
Vad som hade skett misshagade Gud, och han hemsökte Israel.
Då sade David till Gud: »Jag har syndat storligen däri att jag har gjort detta; men tillgiv nu din tjänares missgärning, ty jag har handlat mycket dåraktigt.»
Men HERREN talade till Gad, Davids siare, och sade:
»Gå och tala till David och säg: Så säger HERREN: Tre ting lägger jag fram för dig; välj bland dem ut åt dig ett som du vill att jag skall göra dig.»
Då gick Gad in till David och sade till honom: »Så säger HERREN:
Tag vilketdera du vill: antingen hungersnöd i tre år, eller förödelse i tre månader genom dina ovänners anfall, utan att du kan undkomma dina fienders svärd, eller HERRENS svärd och pest i landet under tre dagar, i det att HERRENS ängel sprider fördärv inom hela Israels område.
Eftersinna nu vilket svar jag skall giva honom som har sänt mig.»
David svarade Gad: »Jag är i stor vånda.
Men låt mig då falla i HERRENS hand, ty hans barmhärtighet är mycket stor; i människohand vill jag icke falla.»
Så lät då HERREN pest komma i Israel, så att sjuttio tusen män av Israel föllo.
Och Gud sände en ängel mot Jerusalem till att fördärva det.
Men när denne höll på att fördärva, såg HERREN därtill och ångrade det onda, så att han sade till ängeln, Fördärvaren: »Det är nog; drag nu din hand tillbaka.»
Och HERRENS ängel stod då vid jebuséen Ornans tröskplats.
När nu David lyfte upp sina ögon och fick se HERRENS ängel stående mellan jorden och himmelen med ett blottat svärd i sin hand, uträckt över Jerusalem, då föllo han och de äldste, höljda i sorgdräkt, ned på sina ansikten.
Och David sade till Gud: »Det var ju jag som befallde att folket skulle räknas.
Det är då jag som har syndat och gjort vad ont är; men dessa, min hjord, vad hava de gjort?
HERRE, min Gud, må din hand vända sig mot mig och min faders hus, men icke mot ditt folk, så att det bliver hemsökt.»
Men HERRENS ängel befallde Gad att säga till David att David skulle gå åstad och resa ett altare åt HERREN på jebuséen Ornans tröskplats.
Och David gick åstad på grund av det ord som Gad hade talat i HERRENS namn.
Då Ornan nu vände sig om, fick han se ängeln; och hans fyra söner som voro med honom, gömde sig.
Men Ornan höll på att tröska vete.
Och David kom till Ornan; när då Ornan såg upp och fick se David, gick han fram ifrån tröskplatsen och föll ned till jorden på sitt ansikte för David.
Och David sade till Ornan: »Giv mig den plats där du tröskar din säd, så att jag där kan bygga ett altare åt HERREN; giv mig den för full betalning; och må så hemsökelsen upphöra bland folket.»
Då sade Ornan till David: »Tag den, och må sedan min herre konungen göra vad honom täckes.
Se, här giver jag dig fäkreaturen till brännoffer och tröskvagnarna till ved och vetet till spisoffer; alltsammans giver jag.»
Men konung David svarade Ornan: »Nej, jag vill köpa det för full betalning; ty jag vill icke taga åt HERREN det som är ditt, och offra brännoffer som jag har fått för intet.»
Och David gav åt Ornan för platsen sex hundra siklar guld, i full vikt.
Och David byggde där ett altare åt HERREN och offrade brännoffer och tackoffer.
Han ropade till HERREN, och han svarade honom med eld från himmelen på brännoffersaltaret.
Och på HERRENS befallning stack ängeln sitt svärd tillbaka i skidan.
Då, när David förnam att HERREN hade bönhört honom på jebuséen Ornans tröskplats, offrade han där.
Men HERRENS tabernakel, som Mose hade låtit göra i öknen, stod jämte brännoffersaltaret, vid den tiden på offerhöjden i Gibeon.
Dock vågade David icke komma inför Guds ansikte för att söka honom; så förskräckt var han för HERRENS ängels svärd.
Och David sade: »Här skall HERREN Guds hus stå, och här altaret för Israels brännoffer.»
Och David befallde att man skulle samla tillhopa de främlingar som funnos i Israels land; och han anställde hantverkare, som skulle hugga ut stenar för att därmed bygga Guds hus.
Och David anskaffade järn i myckenhet till spikar på dörrarna i portarna och till krampor, så ock koppar i sådan myckenhet att den icke kunde vägas,
och cederbjälkar i otalig mängd; ty sidonierna och tyrierna förde cederträ i myckenhet till David.
David tänkte nämligen: »Min son Salomo är ung och späd, men huset som skall byggas åt HERREN måste göras övermåttan stort, så att det bliver namnkunnigt och prisat i alla länder; jag vill därför skaffa förråd åt honom.»
Så skaffade David förråd i myckenhet före sin död.
Och han kallade till sig sin son Salomo och bjöd honom att bygga ett hus åt HERREN, Israels Gud.
Och David sade till sin son Salomo: »Jag hade själv i sinnet att bygga ett hus åt HERRENS, min Guds, namn.
Men HERRENS ord kom till mig; han sade: Du har utgjutit blod i myckenhet och fört stora krig; du skall icke bygga ett hus åt mitt namn, eftersom du har utgjutit så mycket blod på jorden, i min åsyn.
Men se, åt dig skall födas en son; han skall bliva en fridsäll man, och jag skall låta honom få fred med alla sina fiender runt omkring; ty Salomo skall han heta, och frid och ro skall jag låta vila över Israel i hans dagar.
Han skall bygga ett hus åt mitt namn; han skall vara min son, och jag skall vara hans fader.
Och jag skall befästa hans konungatron över Israel för evig tid.
Så vare nu HERREN med dig, min son; må du bliva lyckosam och få bygga HERRENS, din Guds, hus, såsom han har lovat om dig.
Må HERREN allenast giva dig klokhet och förstånd, när han sätter dig till härskare över Israel, och förhjälpa dig till att hålla HERRENS, din Guds, lag.
Då skall du bliva lyckosam, om du håller och gör efter de stadgar och rätter som HERREN har bjudit Mose att ålägga Israel.
Var frimodig och oförfärad; frukta icke och var icke försagd.
Och se, trots mitt betryck har jag nu anskaffat till HERRENS hus ett hundra tusen talenter guld och tusen gånger tusen talenter silver, därtill av koppar och järn mer än som kan vägas, ty så mycket är det; trävirke och sten har jag ock anskaffat, och mer må du själv anskaffa.
Arbetare har du ock i myckenhet hantverkare, stenhuggare och timmermän, och därtill allahanda folk som är kunnigt i allt slags annat arbete.
På guldet, silvret, kopparen och järnet kan ingen räkning hållas.
Upp då och gå till verket; och vare HERREN med dig!»
Därefter bjöd David alla Israels furstar att de skulle understödja hans son Salomo; han sade:
»HERREN, eder Gud, är ju med eder och har låtit eder få ro på alla sidor; ty han har givit landets förra inbyggare i min hand, och landet har blivit HERREN och hans folk underdånigt.
Så vänden nu edert hjärta och eder själ till att söka HERREN, eder Gud; och stån upp och byggen HERREN Guds helgedom, så att man kan föra HERRENS förbundsark och vad annat som hör till Guds helgedom in i det hus som skall byggas åt HERRENS namn.»
Och när David blev gammal och levnadsmätt, gjorde han sin son Salomo till konung över Israel.
Och han församlade alla Israels furstar, så ock prästerna och leviterna.
Och leviterna blevo räknade, de nämligen som voro trettio år gamla eller därutöver; och deras antal, antalet av alla personer av mankön, utgjorde trettioåtta tusen.
»Av dessa», sade han, »skola tjugufyra tusen förestå sysslorna vid HERRENS hus, och sex tusen vara tillsyningsmän och domare;
fyra tusen skola vara dörrvaktare och fyra tusen skola lovsjunga HERREN till de instrumenter som jag har låtit göra för lovsången.»
Och David delade dem i avdelningar efter Levis söner, Gerson Kehat och Merari.
Till gersoniterna hörde Laedan och Simei.
Laedans söner voro Jehiel, huvudmannen, Setam och Joel, tillsammans tre.
Simeis söner voro Selomot, Hasiel och Haran, tillsammans tre.
Dessa voro huvudmän för Laedans familjer.
Och Simeis söner voro Jahat, Sina, Jeus och Beria.
Dessa voro Simeis söner, tillsammans fyra.
Jahat var huvudmannen, och Sisa var den andre.
Men Jeus och Beria hade icke många barn; därför fingo de utgöra allenast en familj, en ordning.
Kehats söner voro Amram, Jishar, Hebron och Ussiel, tillsammans fyra.
Amrams söner voro Aron och Mose.
Och Aron blev jämte sina söner för evärdlig tid avskild till att helgas såsom höghelig, till att för evärdlig tid antända rökelse inför HERREN och göra tjänst inför honom och välsigna i hans namn.
Men gudsmannen Moses söner räknades till Levi stam.
Moses söner voro Gersom och Elieser.
Gersoms söner voro Sebuel, huvudmannen.
Och Eliesers söner voro Rehabja, huvudmannen.
Elieser hade inga andra söner; men Rehabjas söner voro övermåttan talrika.
Jishars söner voro Selomit, huvudmannen.
Hebrons söner voro Jeria, huvudmannen, Amarja, den andre, Jahasiel, den tredje, och Jekameam, den fjärde.
Ussiels söner voro Mika, huvudmannen, och Jissia, den andre.
Meraris söner voro Maheli och Musi.
Mahelis söner voro Eleasar och Kis.
När Eleasar dog, lämnade han inga söner efter sig, utan allenast döttrar; men Kis' söner, deras fränder, togo dessa till hustrur.
Musis söner voro Maheli, Eder och Jeremot, tillsammans tre.
Dessa voro Levi barn, efter deras familjer, huvudmännen för familjerna, så många av dem som inmönstrades, vart namn räknat särskilt, var person för sig, de som kunde förrätta sysslor vid tjänstgöringen i HERRENS hus, nämligen de som voro tjugu år gamla eller därutöver.
Ty David sade: »HERREN, Israels Gud, har låtit sitt folk komma till ro, och han har nu sin boning i Jerusalem till evig tid;
därför behöva icke heller leviterna mer bära tabernaklet och alla redskap till tjänstgöringen därvid.»
(Enligt berättelsen om Davids sista tid räknades nämligen av Levi barn de som voro tjugu år gamla eller därutöver.)
De fingo i stället sin plats vid Arons söners sida för tjänstgöringen i HERRENS hus, i vad som rörde förgårdarna och kamrarna och reningen av allt heligt och sysslorna vid tjänstgöringen i Guds hus,
vare sig det gällde skådebröden eller det fina mjölet till spisoffret eller de osyrade tunnkakorna eller plåtarna eller det hopknådade mjölet, eller något mått och mål,
eller att var morgon göra tjänst genom att tacka och lova HERREN, och likaledes var afton,
eller att offra alla brännoffer åt HERREN på sabbaterna, vid nymånaderna och vid högtiderna, till bestämt antal och såsom det var föreskrivet för dem, beständigt, inför HERRENS ansikte.
De skulle iakttaga vad som var att iakttaga vid uppenbarelsetältet och vid det heliga, vad Arons söner, deras bröder, hade att iakttaga vid tjänstgöringen i HERRENS hus.
Och Arons söner hade följande avdelningar: Arons söner voro Nadab och Abihu, Eleasar och Itamar.
Men Nadab och Abihu dogo före sin fader; och de hade inga söner.
Så blevo allenast Eleasar och Itamar präster.
Och David jämte Sadok, av Eleasars söner, och Ahimelek, av Itamars söner, indelade dem och bestämde den ordning i vilken de skulle göra tjänst.
Då nu Eleasars söner befunnos hava flera huvudmän än Itamars söner, indelade man dem så, att Eleasars söner fingo sexton huvudmän för sina familjer och Itamars söner åtta huvudmän för sina familjer.
Man indelade dem genom lottkastning, de förra såväl som de senare, ty helgedomens furstar och Guds furstar togos både av Eleasars söner och av Itamars söner.
Och Semaja, Netanels son, sekreteraren, av Levi stam, tecknade upp dem i närvaro av konungen, furstarna och prästen Sadok och Ahimelek, Ebjatars son, och i närvaro av huvudmännen för prästernas och leviternas familjer.
Lotterna drogos skiftevis för Eleasars och för Itamars familjer.
Den första lotten föll ut för Jojarib, den andra för Jedaja,
den tredje för Harim, den fjärde för Seorim,
den femte för Malkia, den sjätte för Mijamin,
den sjunde för Hackos, den åttonde för Abia,
den nionde för Jesua, den tionde för Sekanja,
den elfte för Eljasib, den tolfte för Jakim,
den trettonde för Huppa, den fjortonde för Jesebab,
den femtonde för Bilga, den sextonde för Immer,
den sjuttonde för Hesir, den adertonde för Happisses,
den nittonde för Petaja, den tjugonde för Hesekiel,
den tjuguförsta för Jakin, den tjuguandra för Gamul,
den tjugutredje for Delaja, den tjugufjärde för Maasja.
Detta blev den ordning i vilken de skulle göra tjänst, när de gingo in i HERRENS hus, såsom det var föreskrivet för dem genom deras fader Aron, i enlighet med vad HERREN, Israels Gud, hade bjudit honom.
Vad angår de övriga Levi barn, så hörde till Amrams barn Subael, till Subaels barn Jedeja,
till Rehabja, det är till Rehabjas barn, huvudmannen Jissia,
till jishariterna Selomot, till Selomots barn Jahat.
Och benajiter voro Jeria, Amarja, den andre, Jahasiel, den tredje, och Jekameam, den fjärde.
Ussiels barn voro Mika; till Mikas barn hörde Samur.
Mikas broder var Jissia; till Jissias barn hörde Sakarja.
Meraris barn voro Maheli och Musi, Jaasia-Benos söner.
Meraris barn voro dessa av Jaasia-Beno, och vidare Soham, Sackur och Ibri.
Mahelis son var Eleasar, men denne hade inga söner.
Till Kis, det är Kis' barn, hörde Jerameel.
Men Musis barn voro Maheli, Eder och Jerimot.
Dessa voro leviternas barn, efter deras familjer.
Också dessa kastade lott likasåväl som deras bröder, Arons söner, i närvaro av konung David, Sadok, Ahimelek och huvudmännen för prästernas och leviternas familjer, huvudmännen för familjerna likasåväl som deras yngsta bröder.
Och David jämte härhövitsmännen avskilde till tjänstgöring Asafs, Hemans och Jedutuns söner, som hade profetisk anda till att spela på harpor, psaltare och cymbaler.
Och detta är förteckningen på dem, på de män som fingo denna tjänstgöring till åliggande.
Av Asafs söner: Sackur, Josef, Netanja och Asarela, Asafs söner, under ledning av Asaf, som hade profetisk anda till att spela, under konungens ledning.
Av Jedutun: Jedutuns söner Gedalja, Seri, Jesaja, Hasabja och Mattitja, tillsammans sex, med harpor, under ledning av sin fader Jedutun, som hade profetisk anda till att spela tack- och lovsånger till HERREN.
Av Heman: Hemans söner Buckia, Mattanja, Ussiel, Sebuel och Jerimot, Hananja, Hanani, Eliata, Giddalti och Romamti-Eser, Josbekasa, Malloti, Hotir, Mahasiot.
Alla dessa voro söner till Heman, som var konungens siare, enligt det löfte Gud hade givit, att han ville upphöja hans horn; därför gav Gud Heman fjorton söner och tre döttrar.
Alla dessa stodo var och en under sin faders ledning, när de utförde sången i HERRENS hus till cymbaler, psaltare och harpor och så gjorde tjänst i Guds hus; de stodo under konungens, Asafs, Jedutuns och Hemans ledning.
Och antalet av dem jämte deras bröder, av dem som hade blivit undervisade i sången till HERREN ära, alla de däri kunniga, utgjorde två hundra åttioåtta.
Och de kastade lott om tjänstgöringen, alla, den minste likasåväl som den störste, den kunnige jämte lärjungen.
Den första lotten kom ut för Asaf och föll på Josef; den andre blev Gedalja, han själv med sina bröder och söner, tillsammans tolv;
den tredje blev Sackur, med sin söner och bröder, tillsammans tolv
den fjärde lotten kom ut för Jisri, med hans söner och bröder, tillsammans tolv;
den femte blev Netanja, med sina söner och bröder, tillsammans tolv;
den sjätte blev Buckia, med sina söner och bröder, tillsammans tolv;
den sjunde blev Jesarela, med sina söner och bröder, tillsammans tolv;
den åttonde blev Jesaja, med sin söner och bröder, tillsammans tolv
den nionde blev Mattanja, med sina söner och bröder, tillsammans tolv;
den tionde blev Simei, med sina söner och bröder, tillsammans tolv
den elfte blev Asarel, med sin söner och bröder, tillsammans tolv
den tolfte lotten kom ut för Hasabja, med hans söner och bröder tillsammans tolv;
den trettonde blev Subael, med sina söner och bröder, tillsammans tolv;
den fjortonde blev Mattitja, med sina söner och bröder, tillsammans tolv;
den femtonde lotten kom ut för Jeremot, med hans söner och bröder, tillsammans tolv;
den sextonde för Hananja, med hans söner och bröder, tillsammans tolv;
den sjuttonde för Josbekasa, med hans söner och bröder, tillsammans tolv;
den adertonde för Hanani, med hans söner och bröder, tillsammans tolv;
den nittonde för Malloti, med hans söner och bröder, tillsammans tolv;
den tjugonde för Elijata, med hans söner och bröder, tillsammans tolv;
den tjuguförsta för Hotir, med hans söner och bröder, tillsammans tolv;
den tjuguandra för Giddalti, med hans söner och bröder, tillsammans tolv;
den tjugutredje för Mahasiot, med hans söner och bröder, tillsammans tolv;
den tjugufjärde för Romamti-Eser, med hans söner och bröder, tillsammans tolv.
Vad angår dörrvaktarnas avdelningar, så hörde till koraiterna Meselemja, Kores son, av Asafs barn.
Och Meselemja hade söner: Sakarja var den förstfödde, Jediael den andre, Sebadja den tredje, Jatniel den fjärde,
Elam den femte, Johanan den sjätte, Eljoenai den sjunde.
Och Obed-Edom hade söner: Semaja var den förstfödde, Josabad den andre, Joa den tredje, Sakar den fjärde, Netanel den femte,
Ammiel den sjätte, Isaskar den sjunde, Peulletai den åttonde; ty Gud hade välsignat honom.
Åt hans son Semaja föddes ock söner, som blevo furstar inom sin familj, ty de voro dugande män.
Semajas söner voro Otni, Refael och Obed, Elsabad och hans bröder, dugliga män, Elihu och Semakja.
Alla dessa hörde till Obed-Edoms avkomlingar, de själva och deras söner och bröder, dugliga och kraftfulla män i tjänsten, tillsammans sextiotvå avkomlingar av Obed-Edom.
Meselemja hade ock söner och bröder, dugliga män, tillsammans aderton.
Och Hosa, av Meraris barn, hade söner: Simri var huvudmannen, ty visserligen var han icke förstfödd, men hans fader insatte honom till huvudman;
Hilkia var den andre, Tebalja den tredje, Sakarja den fjärde.
Hosas söner och bröder voro tillsammans tretton.
Dessa avdelningar av dörrvaktarna, nämligen dessa deras huvudmän, fingo nu, likasåväl som deras bröder, sina åligganden för att göra tjänst i HERRENS hus.
Och om var port kastade de lott, den minste såväl som den störste, efter sina familjer.
Den lott som angav öster föll då på Selemja; och för hans son Sakarja, en rådklok man, kastade man lott, och för honom kom ut den lott som angav norr;
för Obed-Edom den lott som angav söder, under det att hans söner fingo på sin del förrådshuset;
för Suppim och för Hosa den lott som angav platsen västerut, vid Salleketporten, där vägen höjer sig uppåt, det ena vaktstället invid det andra.
Österut voro sex leviter, norrut fyra för var dag, söderut fyra för var dag, och vid förrådshuset två i sänder;
vid Parbar västerut voro fyra vid vägen och två vid själva Parbar.
Dessa voro dörrvaktarnas avdelningar, av koraiternas barn och av Meraris barn.
Och av leviterna hade Ahia uppsikten över Guds hus skatter och vården om de förråd som utgjordes av vad som hade blivit helgat åt HERREN.
Laedans barn, nämligen gersoniternas barn av Laedans släkt, huvudmannen för gersoniten Laedans familj, jehieliterna,
det är jehieliternas barn, Setam och hans broder Joel, hade uppsikten över skatterna i HERRENS hus.
Vad angår amramiterna, jishariterna, hebroniterna och ossieliterna,
så var Sebuel, son till Gersom, son till Mose, överuppsyningsman över skatterna.
Och hans bröder av Eliesers släkt voro dennes son Rehabja, dennes son Jesaja, dennes son Joram, dennes son Sikri och dennes son Selomot.
Denne Selomot och hans bröder hade uppsikten över alla förråd som utgjordes av vad som hade blivit helgat åt HERREN av konung David, så ock av huvudmännen för familjerna, ävensom av över- och underhövitsmännen och av härhövitsmännen.
Från krigen och av bytet hade de helgat detta för att hålla HERRENS hus vid makt;
likaledes allt vad siaren Samuel och Saul, Kis' son, och Abner, Ners son, och Joab, Serujas son, hade helgat -- korteligen, var och en som helgade något lämnade det under Selomits och hans bröders vård.
Av jishariterna togos Kenanja och hans söner till de världsliga sysslorna i Israel, till att vara tillsyningsmän och domare.
Av hebroniterna togos Hasabja och hans bröder, dugliga män, ett tusen sju hundra, till ämbetsförvaltningen i Israel på andra sidan Jordan, på västra sidan, till alla slags sysslor åt HERREN och till konungens tjänst.
För hebroniterna var Jeria huvudman, för hebroniterna efter deras ättföljd och familjer.
(I Davids fyrtionde regeringsår anställdes undersökning rörande dem; och bland dem funnos då dugande män i Jaeser i Gilead.)
Hans bröder, dugliga män, vore två tusen sju hundra, huvudmän för familjer.
Dem satte konung David över rubeniterna, gaditerna och ena hälften av Manasse stam, för att ombesörja alla Guds och konungens angelägenheter.
Och detta är förteckningen på Israels barn, efter deras antal med huvudmännen för deras familjer och med över- och underhövitsmännen och med deras tillsyningsmän vilka tjänade konungen i allt som rörde krigsfolkets avdelningar, vilka avdelningar kommo och avgingo skiftevis för var och en av årets alla månader, var avdelning tjugufyra tusen man stark.
Över den första avdelningen, den som tjänstgjorde under första månaden, hade Jasobeam, Sabdiels son, befälet.
Och i hans avdelning voro tjugufyra tusen.
Han hörde till Peres' barn och var huvudanförare för alla härhövitsmän som tjänstgjorde under första månaden.
Över den andra månadens avdelning hade ahoaiten Dodai befälet, det var hans avdelning; där var ock fursten Miklot.
Och i hans avdelning voro tjugufyra tusen.
Den tredje härhövitsmannen, den som tjänstgjorde under tredje månaden, var Benaja, prästen Jojadas son, såsom huvudanförare.
Och i hans avdelning voro tjugufyra tusen.
Denne Benaja var en hjälte bland de trettio och hade befälet över de trettio.
Och vid hans avdelning var hans son Ammisabad.
Den fjärde, den som tjänstgjorde under fjärde månaden, var Asael, Joabs broder, och efter honom hans son Sebadja.
Och i hans avdelning voro tjugufyra tusen
Den femte, den som tjänstgjorde under femte månaden, var hövitsmannen Samhut, jisraiten.
Och i hans avdelning voro tjugufyra tusen.
Den sjätte, den som tjänstgjorde under sjätte månaden, var tekoaiten Ira, Ickes' son.
Och i hans avdelning voro tjugufyra tusen.
Den sjunde, den som tjänstgjorde under sjunde månaden, var peloniten Heles, av Efraims barn.
Och i hans avdelning voro tjugufyra tusen.
Den åttonde, den som tjänstgjorde under åttonde månaden, var husatiten Sibbekai, som hörde till seraiterna.
Och i hans avdelning voro tjugufyra tusen.
Den nionde, den som tjänstgjorde under nionde månaden, var anatotiten Abieser, som hörde till benjaminiterna.
Och i hans avdelning voro tjugufyra tusen.
Den tionde, den som tjänstgjorde under tionde månaden, var netofatiten Maherai, som hörde till seraiterna.
Och i hans avdelning voro tjugufyra tusen.
Den elfte, den som tjänstgjorde under elfte månaden, var pirgatoniten Benaja, av Efraims barn.
Och i hans avdelning voro tjugufyra tusen.
Den tolfte, den som tjänstgjorde under tolfte månaden, var netofatiten Heldai, som hörde till Otniels släkt.
Och i hans avdelning voro tjugufyra tusen.
Och Israels stamhövdingar voro dessa: furste för rubeniterna var Elieser, Sikris son; för simeoniterna Sefatja, Maakas son;
för Levi Hasabja, Kemuels son; för Arons släkt Sadok;
för Juda Elihu, en av Davids bröder; för Isaskar Omri, Mikaels son;
för Sebulon Jismaja, Obadjas son; för Naftali Jerimot, Asriels son;
för Efraims barn Hosea, Asasjas son; för ena hälften av Manasse stam Joel, Pedajas son;
för andra hälften av Manasse, den i Gilead, Jiddo, Sakarjas son; för Benjamin Jaasiel, Abners son;
för Dan Asarel, Jerohams son.
Dessa voro Israels stamhövdingar.
Men David tog i förteckningen icke upp dem som voro under tjugu år, ty HERREN hade lovat att han ville föröka Israel såsom stjärnorna på himmelen.
Joab, Serujas son, begynte räkningen, men fullbordade den icke, ty genom den kom förtörnelse över Israel; och antalet togs icke upp i någon förteckning i konung Davids krönika.
Uppsikten över konungens skatter hade Asmavet, Adiels son; över förråden på fälten, i städerna och byarna och fästningstornen Jonatan, Ussias son;
över dem som arbetade på fältet med jordbruket Esri, Kelubs son;
över vingårdarna ramatiten Simei; över de vinförråd som man hade samlat i vingårdarna sifmiten Sabdi;
över olivplanteringarna och mullbärsfikonträden i Låglandet gaderiten Baal-Hanan; över oljeförråden Joas.
Över de fäkreatur som betade i Saron saroniten Sitrai, och över fäkreaturen i dalarna Safat, Adlais son;
över kamelerna ismaeliten Obil; över åsninnorna meronotiten Jedeja;
över småboskapen hagariten Jasis.
Alla dessa voro uppsyningsmän över konung Davids ägodelar.
Men Jonatan, Davids farbroder, var rådgivare; han var en förståndig och skriftlärd man.
Jehiel, Hakmonis son, var anställd hos konungens söner.
Ahitofel var konungens rådgivare, och arkiten Husai var konungens vän.
Efter Ahitofel kom Jojada, Benajas son, och Ebjatar.
Och Joab var konungens härhövitsman.
Och David församlade till Jerusalem alla Israels hövdingar, stamhövdingarna och häravdelningarnas hövitsmän, dem som voro i konungens tjänst, och över- och underhövitsmännen och uppsyningsmännen över alla konungens och hans söners ägodelar och boskap, så ock hovmännen och hjältarna och alla tappra stridsmän.
Och konung David stod upp från sin plats och sade: »Hören mig, mina bröder och mitt folk.
Jag hade själv i sinnet att bygga ett hus till vilostad för HERRENS förbundsark och för vår Guds fotapall, och jag hade skaffat förråd till byggnadsverket.
Men Gud sade till mig: 'Du skall icke bygga ett hus åt mitt namn, ty du är en krigsman och har utgjutit blod.'
Dock utvalde HERREN, Israels Gud mig ur hela min faders hus till att vara konung över Israel evärdligen.
Ty Juda utvalde han till furste, och i Juda hus min faders hus, och bland min faders söner hade han behag till mig, så att han gjorde mig till konung över hela Israel.
Och bland alla mina söner -- ty HERREN har givit mig många söner -- utvalde han min son Salomo till att sitta på HERRENS konungatron och härska över Israel.
Och han sade till mig: 'Din son Salomo är den som skall bygga mitt hus och mina förgårdar; ty honom har jag utvalt till min son, och jag skall vara hans fader.
Och jag skall befästa hans konungamakt för evigt, om han är ståndaktig i att göra efter mina bud och rätter, såsom han nu gör.'
Och nu säger jag inför hela Israel, HERRENS församling, och inför vår Gud, som hör det: Hållen och akten på alla HERRENS, eder Guds, bud, så att I fån besitta det goda landet och lämna det såsom arv åt edra barn efter eder till evärdlig tid.
Och du, min son Salomo, må lära känna din faders Gud och tjäna honom med hängivet hjärta och med villig själ; ty HERREN rannsakar alla hjärtan och förstår alla uppsåt och tankar.
Om du söker honom, så låter han sig finnas av dig, men om du övergiver honom, då förkastar han dig evinnerligen.
Så se nu till; ty HERREN har utvalt dig att bygga ett hus till helgedomen.
Var frimodig och gå till verket.»
Och David gav åt sin son Salomo en mönsterbild av förhuset och tempelbyggnaderna, och av förrådskamrarna, de övre salarna och de inre rummen, och av nådastolens boning;
vidare en mönsterbild av allt som han hade tänkt ut i sitt sinne rörande förgårdarna till HERRENS hus, och rörande alla kamrarna runt omkring för Guds hus' skatter och för de förråd som utgjordes av vad som hade blivit helgat åt HERREN;
vidare föreskrifter rörande prästernas och leviternas avdelningar och alla sysslor som skulle förekomma vid tjänstgöringen i HERRENS hus, och rörande alla kärl som skulle användas vid tjänstgöringen i HERRENS hus,
och rörande guldet, med uppgift på den vikt i guld, som kom på vart särskilt kärl till tjänstgöringen, och rörande alla kärl av silver, med uppgift på den vikt som kom på vart särskilt kärl till tjänstgöringen.
Och han angav vikten på de gyllene ljusstakarna med tillhörande lampor av guld, med uppgift på vikten i var särskild ljusstake med dess lampor, så ock rörande silverljusstakarna, med uppgift på vikten i var ljusstake med dess lampor, alltefter beskaffenheten av den tjänstförrättning vid vilken ljusstaken skulle användas;
likaledes rörande vikten på guldet till skådebrödsborden, vart bord för sig, och rörande silvret till silverborden.
Och han gav honom föreskrifter rörande gafflarna och skålarna och kannorna av rent guld, och rörande de gyllene bägarna, med uppgift på vikten i var särskild bägare, och rörande silverbägarna, med uppgift på vikten i var särskild bägare;
likaså rörande rökelsealtaret av rent guld, med uppgift på vikten; så ock en mönsterbild av vagnen, de gyllene keruberna, som skulle breda ut sina vingar och övertäcka HERRENS förbundsark.
»Om alltsammans», sade han, »har HERREN undervisat mig genom en skrift av sin hand, om allt som skall utföras enligt mönsterbilden.»
Och David sade till sin son Salomo: »Var frimodig och oförfärad och gå till verket; frukta icke och var icke försagd.
Ty HERREN Gud, min Gud, skall vara med dig.
Han skall icke lämna dig och icke övergiva dig, till dess att allt som skall utföras för tjänstgöringen i HERRENS hus har blivit fullbordat.
Och se, här äro prästernas och leviternas avdelningar, som skola förrätta allt slags tjänst i Guds hus.
Och till allt som skall utföras har du hos dig allahanda villigt folk, utrustat med vishet till allt slags arbete; därjämte äro hövdingarna och allt folket redo till allt vad du befaller.»
Och konung David sade till hela församlingen: »Min son Salomo den ende som Gud har utvalt, är ung och späd, och arbetet är stort, ty denna borg är icke avsedd för en människa, utan för HERREN Gud.
Därför har jag, så vitt jag har förmått, för min Guds hus anskaffat guld till det som skall vara av guld, silver till det som skall vara av silver, koppar till det som skall vara av koppar, järn till det som skall vara av järn, och trä till det som skall vara av trä, dessutom onyxstenar och andra infattningsstenar, svartglänsande och brokiga stenar, korteligen, alla slags dyrbara stenar, så ock marmor i myckenhet.
Och därjämte, eftersom jag har min Guds hus kärt, giver jag nu vad jag själv äger i guld och silver till min Guds hus, utöver allt vad jag förut har anskaffat för det heliga huset:
tre tusen talenter guld, guld från Ofir, och sju tusen talenter renat silver till att därmed överdraga byggnadernas väggar,
till att göra av guld vad som skall vara av guld, och till att göra av silver vad som skall vara av silver, ja, till allt slags arbete som utföres av konstnärer.
Vill då någon annan nu i dag frivilligt fylla sin hand med gåvor åt HERREN?»
Då kommo frivilligt familjehövdingarna och Israels stamhövdingar, så ock över- och underhövitsmännen och tillika uppsyningsmännen över konungens arbeten,
och de gåvo till arbetet på Guds hus fem tusen talenter guld, tio tusen dariker, tio tusen talenter silver, aderton tusen talenter koppar och ett hundra tusen talenter järn.
Och var och en som hade ädla stenar i sin ägo gav dem till skatten i HERRENS hus, under gersoniten Jehiels vård.
Då gladde sig folket över deras frivilliga gåvor, ty av hängivet hjärta buro de fram sina frivilliga gåvor åt HERREN; konung David gladde sig ock högeligen.
Och David lovade HERREN inför hela församlingen; David sade: »Lovad vare du, HERRE, vår fader Israels Gud, från evighet till evighet!
Dig, HERRE, tillhör storhet och makt och härlighet och glans och majestät, ja, allt vad i himmelen och på jorden är.
Ditt, o HERRE, är riket, och du har upphöjt dig till ett huvud över allt.
Rikedom och ära komma från dig, du råder över allt, och i din hand är kraft och makt; det står i din hand att göra vad som helst stort och starkt.
Så tacka vi dig nu, vår Gud, och lova ditt härliga namn.
Ty vad är väl jag, och vad är mitt folk, att vi själva skulle förmå att giva sådana frivilliga gåvor?
Nej, från dig kommer allt, och ur din hand hava vi givit det åt dig.
Ty vi äro främlingar hos dig och gäster såsom alla våra fäder; såsom en skugga äro våra dagar på jorden, och intet är här att lita på.
HERRE, vår Gud, alla dessa håvor som vi hava anskaffat för att bygga dig ett hus åt ditt heliga namn -- från din hand hava de kommit, och ditt är alltsammans.
Och jag vet, min Gud, att du prövar hjärtat och har behag till vad rätt är.
Med rättsinnigt hjärta har jag burit fram alla dessa frivilliga gåvor; och nu har jag ock sett med glädje huru ditt folk, som står har, har burit fram åt dig sina frivilliga gåvor.
HERRE, Abrahams, Isaks och Israels, våra fäders, Gud, låt evinnerligen ditt folks hjärtas håg och tankar vara redo till sådant, och vänd deras hjärtan till dig.
Och giv min son Salomo ett hängivet hjärta, så att han håller dina bud, dina vittnesbörd och dina stadgar, och utför allt detta och bygger denna borg, vartill jag har skaffat förråd.»
Därefter sade David till hela församlingen: »Loven HERREN, eder Gud.»
Då lovade hela församlingen HERREN, sina fäders Gud, och de bugade sig och föllo ned för HERREN och för konungen.
Och dagen efter denna dag slaktade de slaktoffer åt HERREN och offrade brännoffer åt HERREN: tusen tjurar, tusen vädurar och tusen lamm med tillhörande drickoffer, därtill slaktoffer i myckenhet för hela Israel.
Och de åto och drucko inför HERRENS ansikte på den dagen med stor glädje.
Och de gjorde för andra gången Salomo, Davids son, till konung; de smorde honom till en HERRENS furste, och Sadok till präst.
Och så satt Salomo på HERRENS tron såsom konung efter sin fader David, och han blev lyckosam; och hela Israel lydde honom.
Och alla hövdingarna och hjältarna och därjämte alla konung Davids söner underkastade sig konung Salomo.
Och HERREN gjorde Salomo övermåttan stor inför hela Israel, och lät hans konungsliga härlighet bliva större än någons som före honom hade varit konung över Israel.
Men David, Isais son, hade regerat över hela Israel.
Den tid han regerade över Israel var fyrtio år; i Hebron regerade han i sju år, och i Jerusalem regerade han i trettiotre år.
Och han dog i en god ålder, mätt på att leva och mätt på rikedom och ära.
Och hans son Salomo blev konung efter honom.
Och vad som är att säga om konung David, om hans första tid såväl som om hans sista, det finnes upptecknat i siaren Samuels krönika, i profeten Natans krönika och i siaren Gads krönika,
tillika med hela hans regering och hans bedrifter och de skickelser som övergingo honom och Israel och alla andra länder och riken.
Salomo, Davids son, befäste sig nu i sin konungamakt, i det att HERREN, hans Gud, var med honom och gjorde honom övermåttan stor.
Och sedan Salomo hade låtit kallelse utgå till hela Israel, till över- och underhövitsmännen, till domarna och till alla hövdingar i hela Israel, huvudmännen för familjerna,
begav han sig med hela denna församling till offerhöjden i Gibeon, ty där stod Guds uppenbarelsetält, som HERRENS tjänare Mose hade gjort i öknen.
Guds ark däremot hade David hämtat från Kirjat-Jearim upp till den plats som David hade berett åt den, ty han hade åt den slagit upp ett tält i Jerusalem.
Men kopparaltaret, som Besalel, son till Uri, son till Hur, hade gjort, det hade man ställt upp framför HERRENS tabernakel; och Salomo och församlingen gingo dit för att fråga honom.
Där offrade nu Salomo inför HERRENS ansikte på kopparaltaret, som stod vid uppenbarelsetältet; han offrade på det tusen brännoffer.
Och om natten uppenbarade sig Gud för Salomo; han sade till honom: »Bed mig om vad du vill att jag skall giva dig.»
Salomo svarade Gud: »Du har gjort stor nåd med min fader David och har låtit mig bliva konung efter honom.
Så låt nu, HERRE Gud, ditt ord till min fader David visa sig vara sant; ty du har själv gjort mig till konung över ett folk som är så talrikt som stoftet på jorden.
Giv mig nu vishet och förstånd till att vara detta folks ledare och anförare; ty vem skulle eljest kunna vara domare för detta ditt stora folk?»
Då sade Gud till Salomo: »Eftersom du är så till sinnes, och icke har bett om rikedom, skatter och ära eller om dina ovänners liv, och ej heller bett om långt liv, utan har bett om vishet och förstånd, så att du kan vara domare för mitt folk, över vilket jag har gjort dig till konung,
därför vare vishet och förstånd dig givna; därtill vill jag ock giva dig rikedom och skatter och ära, så att ingen konung före dig har haft och ej heller någon efter dig skall hava så mycket därav.»
Sedan nu Salomo hade varit vid offerhöjden i Gibeon, begav han sig från uppenbarelsetältet till Jerusalem och regerade där över Israel.
Och Salomo samlade vagnar och ridhästar, så att han hade ett tusen fyra hundra vagnar och tolv tusen ridhästar; dem förlade han dels i vagnsstäderna, dels i Jerusalem, hos konungen själv.
Och konungen styrde så, att silver och guld blev lika vanligt i Jerusalem som stenar, och cederträ lika vanligt som mullbärsfikonträ i Låglandet.
Och hästarna som Salomo lät anskaffa infördes från Egypten; ett antal kungliga uppköpare hämtade ett visst antal av dem till bestämt pris.
Var vagn som de hämtade upp från Egypten och införde kostade sex hundra siklar silver, och var häst ett hundra femtio.
Sammalunda infördes ock genom deras försorg sådana till hetiternas alla konungar och till konungarna i Aram.
Och Salomo tänkte nu på att bygga ett hus åt HERRENS namn och ett hus åt sig själv till konungaboning.
Därför avräknade Salomo sjuttio tusen män till att vara bärare, åttio tusen man till att hugga sten i bergen, och tre tusen sex hundra till att hava uppsikt över de andra.
Och Salomo sände till Huram, konungen i Tyrus, och lät säga: »Visa samma vänskap mot mig som mot min fader David, till vilken du sände cederträ, för att han skulle bygga sig ett hus att bo i.
Nu vill jag bygga ett hus åt HERRENS, min Guds, namn och helga det åt honom, för att man där må antända välluktande rökelse inför hans ansikte, och hava skådebröden beständigt upplagda, och offra brännoffer morgon och afton, på sabbaterna, vid nymånaderna och vid HERRENS, vår Guds, högtider; ty så är det för evärdlig tid stadgat för Israel.
Och det hus som jag vill bygga skall vara stort, ty vår Gud är större än alla andra gudar.
Vem förmår väl att bygga honom ett hus?
Himlarna och himlarnas himmel rymma honom ju icke.
Vem är då jag, att jag skulle kunna bygga honom ett hus, om icke för att antända rökelse inför hans ansikte?
Så sänd mig nu en konstförfaren man som kan arbeta i guld, silver, koppar och järn, så ock i purpurrött, karmosinrött och mörkblått garn, och som är skicklig i att utföra snidverk, tillsammans med de konstförfarna män som jag har hos mig här i Juda och Jerusalem, och som min fader David har anställt.
Och sänd mig cederträ, cypressträ och algumträ från Libanon, ty jag vet att dina tjänare äro skickliga i att hugga virke på Libanon; och mina tjänare äro redo att vara dina tjänare behjälpliga.
Må du skaffa mig virke i myckenhet, ty huset som jag vill bygga skall vara stort och härligt.
Och jag är villig att åt timmermännen som hugga virket giva, för dina tjänares räkning, tjugu tusen korer tröskat vete, tjugu tusen korer korn, tjugu tusen bat vin och tjugu tusen bat olja.»
Härpå svarade Huram, konungen i Tyrus, i ett brev som han sände till Salomo: »Därför att HERREN älskar sitt folk, har han satt dig till konung över dem.»
Och Huram skrev ytterligare: »Lovad vare HERREN, Israels Gud, himmelens och jordens skapare, han som har givit konung David en vis son, så utrustad med klokhet och förstånd, att han kan bygga ett hus åt HERREN och ett hus åt sig själv till konungaboning!
Så sänder jag nu en konstförfaren och förståndig man, nämligen Huram-Abi.
Han är son till en av Dans döttrar, och hans fader är en tyrisk man; han är skicklig att arbeta i guld och silver, i koppar, järn, sten och trä, så ock i purpurrött, mörkblått, vitt och karmosinrött garn, och tillika att utföra alla slags snidverk och att väva alla slags konstvävnader; honom må du låta utföra arbetet tillsammans med dina och min herres, din fader Davids, konstförfarna män.
Må alltså nu min herre sända till sina tjänare vetet och kornet, oljan och vinet som han har talat om.
Då vilja vi hugga virke på Libanon, så mycket du behöver, och flotta det till dig på havet till Jafo; men därifrån må du själv låta föra det upp till Jerusalem.»
Och Salomo lät räkna alla främmande män i Israels land, likasom hans fader David förut hade anställt en räkning av dem.
Och de befunnos vara ett hundra femtiotre tusen sex hundra.
Av dem utsåg han sjuttio tusen till att vara bärare, åttio tusen till att hugga sten i bergen, och tre tusen sex hundra till att hava uppsikt över folket och hålla det till arbete.
Och Salomo begynte att bygga HERRENS hus i Jerusalem, på berget Moria, där hans fader David hade fått sin uppenbarelse, och där han nu själv hade berett rum, på det ställe som David hade utsett, nämligen på jebuséen Ornans tröskplats.
Han begynte att bygga på andra dagen i andra månaden, i sitt fjärde regeringsår.
När Salomo då skulle bygga Guds hus, lade han grunden så, att det blev sextio alnar långt och tjugu alnar brett, efter det gamla alnmåttet.
Förhuset, som låg framför långhuset, framför husets kortsida, mätte tjugu alnar, och dess höjd var ett hundra tjugu, och han överdrog det innantill med rent guld.
Huvudbyggnaden beklädde han med cypressträ, detta åter beklädde han med bästa guld, och prydde det med palmer och kedjeverk.
Därjämte smyckade han huset med dyrbara stenar.
Men guldet var från Parvaim.
Och han beklädde huset, bjälkarna, trösklarna, ävensom väggarna och dörrarna däri med guld, och lät inrista keruber på väggarna.
Vidare tillredde han det rum som skulle vara det allraheligaste; det låg utefter husets kortsida och var tjugu alnar långt och tjugu alnar brett.
Och han beklädde det med bästa guld, sex hundra talenter i vikt.
Och spikarna däri vägde femtio siklar i guld.
De övre salarna beklädde han ock med guld.
Och till det rum som var det allraheligaste gjorde han två keruber, i bildhuggeriarbete, och man överdrog dem med guld.
Längden på kerubernas vingar tillsammans var tjugu alnar.
Den enas ena vinge, fem alnar lång, rörde vid husets ena vägg, och hans andra vinge, fem alnar lång, rörde vid den andra kerubens vinge.
Och den andra kerubens ena vinge, fem alnar lång, rörde vid husets andra vägg, och hans andra vinge, fem alnar lång, nådde intill den första kerubens vinge.
Alltså bredde dessa keruber ut sina vingar tjugu alnar vitt, under det att de stodo på sina fötter, med ansiktena vända inåt.
Och han gjorde förlåten av mörkblått, purpurrött, karmosinrött och vitt garn och prydde den med keruber.
Och han gjorde två pelare till att stå framför huset, trettiofem alnar höga; och huvudet som satt ovanpå var och en av dem var fem alnar.
Och han gjorde kedjor till koret och satte ock sådana upptill på pelarna.
Och vidare gjorde han hundra granatäpplen och satte dem på kedjorna.
Och pelarna ställde han upp framför tempelsalen, den ena på högra sidan och den andra på vänstra; åt den högra gav han namnet Jakin och åt den vänstra namnet Boas.
Och han gjorde ett altare av koppar, tjugu alnar långt, tjugu alnar brett och tio alnar högt.
Han gjorde ock havet, i gjutet arbete.
Det var tio alnar från den ena kanten till den andra, runt allt omkring, och fem alnar högt; och ett trettio alnar långt snöre mätte dess omfång.
Och runt omkring nedantill voro bilder som föreställde oxar, och omgåvo det runt omkring -- tio alnar brett som det var -- så att de omslöto havet runt omkring; oxarna bildade två rader och voro gjutna i ett stycke med det övriga.
Det stod ock på tolv oxar, tre vända mot norr, tre vända mot väster, tre vända mot söder och tre vända mot öster; havet stod ovanpå dessa, och deras bakdelar voro alla vända inåt.
Dess tjocklek var en handsbredd; och dess kant var gjord såsom kanten på en bägare, i form av en utslagen lilja.
Det rymde och höll tre tusen bat.
Vidare gjorde han tio bäcken och ställde fem på högra sidan och fem på vänstra, för att brukas vid tvagning; i dem skulle man nämligen skölja vad som hörde till brännoffret.
Men havet var för prästerna till att två sig i.
Vidare gjorde han de gyllene ljusstakarna, tio till antalet, sådana de skulle vara, och ställde dem i tempelsalen, fem på högra sidan och fem på vänstra.
Vidare gjorde han tio bord och satte dem i tempelsalen, fem på högra sidan och fem på vänstra.
Han gjorde ock ett hundra skålar av guld.
Och han gjorde prästernas förgård och den stora yttre förgården, så ock dörrar till denna förgård; och dörrarna överdrog han med koppar.
Och havet ställde han på högra sidan, åt sydost.
Dessutom gjorde Huram askkärlen, skovlarna och skålarna.
Så förde Hiram det arbete till slut, som han fick utföra åt konung Salomo för Guds hus:
nämligen två pelare, och de två kloten och pelarhuvudena ovanpå pelarna, och de två nätverk som skulle betäcka de båda klotformiga pelarhuvuden som sutto ovanpå pelarna,
och därjämte de fyra hundra granatäpplena till de båda nätverken, två rader granatäpplen till vart nätverk, för att de båda klotformiga pelarhuvuden som sutto uppe på pelarna så skulle bliva betäckta.
Vidare gjorde han bäckenställen och gjorde tillika bäckenen på bäckenställen,
så ock havet, som var allenast ett, och de tolv oxarna därunder.
Och askkärlen, skovlarna och gafflarna och alla dithörande föremål gjorde Huram-Abiv åt konung Salomo till HERRENS hus.
Allt var av blank koppar.
På Jordanslätten lät konungen gjuta det i lerformar, mellan Suckot och Sereda.
Och Salomo lät göra en så stor myckenhet av alla dessa föremål, att kopparens vikt icke kunde utrönas.
Alltså gjorde Salomo alla föremål som skulle finnas i Guds hus: det gyllene altaret, borden som skådebröden skulle ligga på,
så ock ljusstakarna med sina lampor, som skulle tändas på föreskrivet sätt, framför koret, av fint guld,
med blomverket, lamporna och lamptängerna av guld -- allt av yppersta guld;
vidare knivarna, de båda slagen av skålar och fyrfaten, av fint guld.
Och vad angår ingångarna i huset, så voro både de dörrar i dess innersta, som ledde till det allraheligaste, och de dörrar i huset, som ledde till tempelsalen, gjorda av guld.
Sedan allt det arbete som Salomo lät utföra för HERRENS hus var färdigt, förde Salomo ditin vad hans fader David hade helgat åt HERREN: silvret, guldet och alla kärlen; detta lade han in i skattkamrarna i Guds hus.
Därefter församlade Salomo de äldste i Israel, alla huvudmännen för stammarna, Israels barns familjehövdingar, till Jerusalem, för att hämta HERRENS förbundsark upp från Davids stad, det är Sion.
Så församlade sig då till konungen alla Israels män under högtiden, den som firades i sjunde månaden.
När då alla de äldste i Israel hade kommit tillstädes, lyfte leviterna upp arken.
Och de hämtade arken och uppenbarelsetältet ditupp, jämte alla heliga föremål som funnos i tältet; de levitiska prästerna hämtade det ditupp.
Och konung Salomo stod framför arken jämte Israels hela menighet, som hade församlats till honom; och de offrade därvid småboskap och fäkreatur i sådan myckenhet, att de icke kunde täljas eller räknas.
Och prästerna buro in HERRENS förbundsark till dess plats i husets kor, i det allraheligaste, till platsen under kerubernas vingar.
Keruberna höllo nämligen sina vingar utbredda över den plats där arken stod, så att arken och dess stänger ovantill övertäcktes av keruberna.
Och stängerna voro så långa, att deras ändar, som sköto ut från arken, väl kunde ses framför koret, men däremot icke voro synliga längre ute.
Och den har blivit kvar där ända till denna dag.
I arken fanns intet annat än de två tavlor som Mose hade lagt dit vid Horeb, när HERREN slöt förbund med Israels barn, sedan de hade dragit ut ur Egypten.
Men när prästerna gingo ut ur helgedomen (ty alla präster som funnos där hade helgat sig, utan avseende på vilken avdelning de tillhörde;
och leviterna, samtliga sångarna, Asaf, Heman och Jedutun med sina söner och bröder, stodo, klädda i vitt linne, med cymbaler, psaltare och harpor öster om altaret, och jämte dem ett hundra tjugu präster som blåste i trumpeter;
och trumpetblåsarna och sångarna stämde på en gång och enhälligt upp HERRENS lov och pris), och när man nu lät trumpeter och cymbaler och andra instrumenter ljuda och begynte lova HERREN, därför att han är god, och därför att hans nåd varar evinnerligen, då blev huset, HERRENS hus, uppfyllt av en molnsky,
så att prästerna för molnskyns skull icke kunde stå där och göra tjänst; ty HERRENS härlighet uppfyllde Guds hus.
Då sade Salomo: »HERREN har sagt att han vill bo i töcknet.
Men jag har byggt ett hus till boning åt dig och berett en plats där du må förbliva till evig tid.»
Sedan vände konungen sig om och välsignade Israels hela församling, under det att Israels hela församling förblev stående.
Han sade: »Lovad vare HERREN, Israels Gud, som med sina händer har fullbordat vad han med sin mun lovade min fader David, i det han sade:
'Från den dag då jag förde mitt folk ut ur Egyptens land har jag icke i någon av Israels stammar utvalt en stad, till att i den bygga ett hus där mitt namn skulle vara, ej heller har jag utvalt någon man till att vara en furste över mitt folk Israel;
men Jerusalem har jag nu utvalt, för att mitt namn skall vara där, och David har jag utvalt till att råda över mitt folk Israel.'
Och min fader David hade väl i sinnet att bygga ett hus åt HERRENS, Israels Guds, namn;
men HERREN sade till min fader David: 'Då du nu har i sinnet att bygga ett hus åt mitt namn, så gör du visserligen väl däri att du har detta i sinnet;
dock skall icke du få bygga detta hus, utan din son, den som har utgått från din länd, han skall bygga huset åt mitt namn.'
Och HERREN har uppfyllt det löfte han gav; ty jag har kommit upp i min fader Davids ställe och sitter nu på Israels tron, såsom HERREN lovade, och jag har byggt huset åt HERRENS, Israels Guds, namn.
Och där har jag satt arken, i vilken förvaras det förbund som HERREN slöt med Israels barn.»
Därefter trädde han fram för HERRENS altare inför Israels hela församling och uträckte sina händer.
Ty Salomo hade gjort en talarstol av koppar, fem alnar lång, fem alnar bred och tre alnar hög, och ställt den mitt på den yttre förgården, på den stod han nu.
Och han föll ned på sina knän inför Israels hela församling, och uträckte sina händer mot himmelen
och sade: »HERRE, Israels Gud, ingen gud är dig lik, i himmelen eller på jorden, du som håller förbund och bevarar nåd mot dina tjänare, när de vandra inför dig av allt sitt hjärta,
du som har hållit vad du lovade din tjänare David, min fader; ty vad du med din mun lovade, det fullbordade du med din hand, så som nu har skett.
Så håll nu ock, HERRE, Israels Gud, vad du lovade din tjänare David, min fader, i det att du sade: 'Aldrig skall den tid komma, då på Israels tron icke inför mig sitter en avkomling av dig, om allenast dina barn hava akt på sin väg, så att de vandra efter min lag, såsom du har vandrat inför mig.'
Så låt nu, HERRE, Israels Gud, det ord som du har talat till din tjänare David bliva sant.
Men kan då Gud verkligen bo på jorden bland människorna?
Himlarna och himlarnas himmel rymma dig ju icke; huru mycket mindre då detta hus som jag har byggt!
Men vänd dig ändå till din tjänares bön och åkallan, HERRE, min Gud, så att du hör på det rop och den bön som din tjänare uppsänder till dig
och låter dina ögon dag och natt vara öppna och vända mot detta hus -- den plats varom du har sagt att du där vill fästa ditt namn -- så att du ock hör den bön som din tjänare beder, vänd mot denna plats.
Ja, hör på de böner som din tjänare och ditt folk Israel uppsända, vända mot denna plats.
Må du höra dem från himmelen, där du bor; och när du hör, så må du förlåta.
Om någon försyndar sig mot sin nästa och man ålägger honom en ed och låter honom svärja, och han så kommer och svär inför ditt altare i detta hus,
må du då höra det från himmelen och utföra ditt verk och skaffa dina tjänare rätt, i det att du vedergäller den skyldige och låter hans gärningar komma över hans huvud, men skaffar rätt åt den som har rätt och låter honom få efter hans rättfärdighet.
Och om ditt folk Israel bliver slaget av en fiende, därför att de hava syndat mot dig, men de omvända sig och prisa ditt namn och bedja och åkalla inför ditt ansikte i detta hus
må du då höra det från himmelen och förlåta ditt folk Israels synd och låta dem komma tillbaka till det land som du har givit åt dem och deras fäder.
Om himmelen bliver tillsluten, så att regn icke faller, därför att de hava syndat mot dig, men de då bedja, vända mot denna plats, och prisa ditt namn och omvända sig från sin synd, när du bönhör dem,
må du då höra det i himmelen och förlåta dina tjänares och ditt folk Israels synd, i det att du lär dem den goda väg som de skola vandra; och må du låta det regna över ditt land, det som du har givit åt ditt folk till arvedel.
Om hungersnöd uppstår i landet, om pest uppstår, om sot och rost, om gräshoppor och gräsmaskar komma, om fienderna tränga folket i det land där deras städer stå, eller om någon annan plåga och sjukdom kommer, vilken det vara må,
och om då någon bön och åkallan höjes från någon människa, vilken det vara må, eller ock från hela ditt folk Israel, när de var för sig känna den plåga och smärta som har drabbat dem, och de så uträcka sina händer mot detta hus,
må du då höra det från himmelen, där du bor, och förlåta och giva var och en efter alla hans gärningar, eftersom du känner hans hjärta -- ty du allena känner människornas hjärtan --
på det att de alltid må frukta dig och vandra på dina vägar, så länge de leva i det land som du har givit åt våra fäder.
Också om en främling, en som icke är av ditt folk Israel, kommer ifrån fjärran land, för ditt stora namns och din starka hands och din uträckta arms skull, om någon sådan kommer och beder, vänd mot detta hus,
må du då från himmelen, där du bor, höra det och göra allt varom främlingen ropar till dig, på det att alla jordens folk må känna ditt namn och frukta dig, likasom ditt folk Israel gör, och förnimma att detta hus som jag har byggt är uppkallat efter ditt namn.
Om ditt folk drager ut till strid mot sina fiender, på den väg du sänder dem, och de då bedja till dig, vända i riktning mot denna stad som du har utvalt och mot det hus som jag har byggt åt ditt namn,
må du då från himmelen höra deras bön och åkallan och skaffa dem rätt.
Om de synda mot dig -- eftersom ingen människa finnes, som icke syndar -- och du bliver vred på dem och giver dem i fiendens våld, så att man tager dem till fånga och för dem bort till något annat land, fjärran eller nära,
men de då besinna sig i det land där de äro i fångenskap, och omvända sig och åkalla dig i fångenskapens land och säga: 'Vi hava syndat, vi hava gjort illa och varit ogudaktiga',
om de så omvända sig till dig av allt sitt hjärta och av all sin själ, i fångenskapens land, dit man har fört dem i fångenskap, och bedja, vända i riktning mot sitt land, det som du har givit åt deras fäder, och mot den stad som du har utvalt, och mot det hus som jag har byggt åt ditt namn,
må du då från himmelen, där du bor, höra deras bön och åkallan och skaffa dem rätt och förlåta ditt folk vad de hava syndat mot dig.
Ja, min Gud, låt nu dina ögon vara öppna och dina öron akta på vad som bedes på denna plats.
Ja: Stå upp, HERRE Gud, och kom till din vilostad, du och din makts ark.
Dina präster, HERRE Gud, vare klädda i frälsning, och dina fromma glädje sig över ditt goda.
HERRE Gud, visa icke tillbaka din smorde; tänk på den nåd du har lovat din tjänare David.
När Salomo hade slutat sin bön, kom eld ned från himmelen och förtärde brännoffret och slaktoffren, och HERRENS härlighet uppfyllde huset.
Och prästerna kunde icke gå in i HERRENS hus, eftersom HERRENS härlighet uppfyllde HERRENS hus.
Då nu alla Israels barn sågo huru elden kom ned, och sågo HERRENS härlighet över huset, föllo de ned på den stenlagda gården, med ansiktena mot jorden, och tillbådo HERREN och tackade honom, därför att han är god, och därför att hans nåd varar evinnerligen.
Och konungen och allt folket offrade slaktoffer inför HERRENS ansikte.
Konung Salomo offrade såsom slaktoffer tjugutvå tusen tjurar och ett hundra tjugu tusen av småboskapen.
Så invigdes Guds hus av konungen och allt folket.
Och prästerna stodo där i sina tjänstförrättningar, och leviterna stodo med HERRENS musikinstrumenter, som konung David hade låtit göra, för att de med dem skulle tacka HERREN, därför att hans nåd varar evinnerligen; David lät nämligen dem utföra lovsången.
Men prästerna stodo mitt emot dem och blåste i trumpeter, medan hela Israel förblev stående.
Och Salomo helgade den mellersta delen av förgården framför HERRENS hus; ty där offrade han brännoffren och fettstyckena av tackoffret eftersom kopparaltaret som Salomo hade låtit göra icke kunde rymma brännoffret, spisoffret och fettstyckena.
Tid detta tillfälle firade Salomo högtiden i sju dagar, och med honom hela Israel, en mycket stor församling ifrån hela landet, allt ifrån det ställe där vägen går till Hamat ända till Egyptens bäck.
Och på åttonde dagen höllo de högtidsförsamling.
Ty altarets invigning firade de i sju dagar och högtiden i sju dagar.
Men på tjugutredje dagen i sjunde månaden lät han folket gå hem till sina hyddor; och de voro fulla av glädje och fröjd över det goda som HERREN hade gjort mot David och Salomo och mot sitt folk Israel.
Så fullbordade Salomo HERRENS hus och konungshuset; och allt vad Salomo hade haft i sinnet att utföra i HERRENS hus och i sitt eget hus hade lyckats honom väl.
Och HERREN uppenbarade sig för Salomo om natten och sade till honom: »Jag har hört din bön och utvalt denna plats åt mig till offerplats.
Om jag tillsluter himmelen, så att regn icke faller, om jag bjuder gräshoppor att fördärva landet, eller om jag sänder pest bland mitt folk,
men mitt folk, det som är uppkallat efter mitt namn, då ödmjukar sig och beder och söker mitt ansikte och omvänder sig från sina onda vägar, så vill jag höra det från himmelen och förlåta deras synd och skaffa bot åt deras land.
Så skola nu mina ögon vara öppna och mina öron akta på vad som bedes på denna plats.
Och nu har jag utvalt och helgat detta hus, för att mitt namn skall vara där till evig tid.
Och mina ögon och mitt hjärta skola vara där alltid.
Om du nu vandrar inför mig, såsom din fader David vandrade, så att du gör allt vad jag har bjudit dig och håller mina stadgar och rätter,
då skall jag upprätthålla din konungatron, såsom jag lovade din fader David, när jag sade: 'Aldrig skall den tid komma, då en avkomling av dig icke råder över Israel.'
Men om I vänden om och övergiven de stadgar och bud som jag har förelagt eder, och gån bort och tjänen andra gudar och tillbedjen dem,
då skall jag rycka upp dem som så göra ur mitt land, det som jag har givit dem; och detta hus som jag har helgat åt mitt namn skall jag förkasta ifrån mitt ansikte; och jag skall göra det till ett ordspråk och en visa bland alla folk.
Och över detta hus, som har varit så upphöjt, skall då var och en som går därförbi bliva häpen.
Och när någon frågar: 'Varför har HERREN gjort så mot detta land och detta hus?',
då skall man svara: 'Därför att de övergåvo HERREN, sina fäders Gud, som hade fört dem ut ur Egyptens land, och höllo sig till andra gudar och tillbådo dem och tjänade dem, därför har han låtit allt detta onda komma över dem.'»
När de tjugu år voro förlidna, under vilka Salomo byggde på HERRENS hus och på sitt eget hus,
byggde Salomo upp de städer som Huram hade givit honom och lät Israels barn bosätta sig i dem.
Och Salomo drog till Hamat-Soba och bemäktigade sig det.
Och han byggde upp Tadmor i öknen och alla de förrådsstäder som i Hamat äro byggda av honom.
Vidare byggde han upp Övre Bet-Horon och Nedre Bet-Horon och gjorde dem till fasta städer med murar, portar och bommar,
så ock Baalat och alla Salomos förrådsstäder, ävensom alla vagnsstäderna och häststäderna, och allt annat som Salomo kände åstundan att bygga i Jerusalem, på Libanon och eljest i hela det land som lydde under hans välde.
Allt det folk som fanns kvar av hetiterna, amoréerna, perisséerna, hivéerna och jebuséerna, korteligen, alla de som icke voro av Israel --
deras avkomlingar, så många som funnos kvar i landet efter dem, i det att Israels barn icke hade utrotat dem, dessa pålade Salomo att vara arbetspliktiga, såsom de äro ännu i dag.
Men somliga av Israels barn gjorde Salomo icke till trälar vid de arbeten han utförde, utan de blevo krigare och hövitsmän för hans kämpar, eller uppsyningsmän över hans vagnar och ridhästar.
Och konung Salomos överfogdar voro två hundra femtio; dessa hade befälet över folket.
Och Salomo lät Faraos dotter flytta upp från Davids stad till det hus som han hade byggt åt henne; ty han sade: »Jag vill icke att någon kvinna skall bo i Davids, Israels konungs, hus, ty det är en helig plats, eftersom HERRENS ark har kommit dit.»
Nu offrade Salomo brännoffer åt HERREN på HERRENS, altare, det som han hade byggt framför förhuset;
han offrade var dag de för den dagen bestämda offren, efter Moses bud, på sabbaterna, vid nymånaderna och vid högtiderna tre gånger om året, nämligen vid det osyrade brödets högtid, vid veckohögtiden och vid lövhyddohögtiden.
Och efter sin fader Davids anordning fastställde han de avdelningar i vilka prästerna skulle tjänstgöra, ävensom leviternas åligganden, att de skulle utföra lovsången och betjäna prästerna -- var dag de för den dagen bestämda åliggandena -- så ock huru dörrvaktarna, efter sina avdelningar, skulle hålla vakt vid de särskilda portarna; ty så hade gudsmannen David bjudit.
Och man vek icke av ifrån vad konungen hade bjudit angående prästerna och leviterna, varken i fråga om någon annan angelägenhet eller i fråga om förråden.
Så utfördes allt Salomos arbete, först intill den dag då grunden lades till HERRENS hus, och sedan intill dess det blev fullbordat.
Och så var då HERRENS hus färdigt.
Vid denna tid drog Salomo till Esjon-Geber och till Elot, på havsstranden, i Edoms land.
Och Huram sände till honom skepp genom sitt folk, och därjämte av sitt folk sjökunnigt manskap.
De foro med Salomos folk till Ofir och hämtade därifrån fyra hundra femtio talenter guld, som de förde till konung Salomo.
När drottningen av Saba fick höra ryktet om Salomo, kom hon för att i Jerusalem sätta Salomo på prov med svåra frågor.
Hon kom med ett mycket stort följe och förde med sig kameler, som buro välluktande kryddor och guld i myckenhet, så ock ädla stenar.
Och när hon kom inför konung Salomo, förelade hon honom allt vad hon hade i tankarna.
Men Salomo gav henne svar på alla hennes frågor; intet var förborgat för Salomo, utan han kunde giva henne svar på allt.
När nu drottningen av Saba såg Salomos vishet, och såg huset som han hade byggt,
och såg rätterna på hans bord och såg huru hans tjänare sutto där, och huru de som betjänade honom utförde sina åligganden, och huru de voro klädda, och vidare såg hans munskänkar, och huru de voro klädda, och när hon såg den trappgång på vilken han gick upp till HERRENS hus, då blev hon utom sig av förundran.
Och hon sade till konungen: »Sant var det tal som jag hörde i mitt land om dig och om din vishet.
Jag ville icke tro vad man sade förrän jag själv kom och med egna ögon fick se det; men nu finner jag att vidden av din vishet icke ens till hälften har blivit omtalad för mig.
Du är vida förmer, än jag genom ryktet hade hört.
Sälla äro dina män, och sälla äro dessa dina tjänare, som beständigt få stå inför dig och höra din visdom.
Lovad vare HERREN, din Gud, som har funnit sådant behag i dig, att han har satt dig på sin tron till att vara konung inför HERREN, din Gud!
Ja, därför att din Gud älskar Israel och vill hålla det vid makt evinnerligen, därför har han satt dig till konung över dem, för att du skall skipa lag och rätt.»
Och hon gav åt konungen ett hundra tjugu talenter guld, så och välluktande kryddor i stor myckenhet, därtill ädla stenar; sådana välluktande kryddor som de vilka drottningen av Saba gav åt konung Salomo hava eljest icke funnits.
När Hirams folk och Salomos folk hämtade guld från Ofir, hemförde också de algumträ och ädla stenar.
Av algumträet lät konungen göra tillbehör till HERRENS hus och till konungshuset, så ock harpor och psaltare för sångarna.
Sådant hade aldrig förut blivit sett i Juda land.
Konung Salomo åter gav åt drottningen av Saba allt vad hon åstundade och begärde, förutom vad som svarade emot det hon hade medfört åt konungen.
Sedan vände hon om och for till sitt land igen med sina tjänare.
Det guld som årligen inkom till Salomo vägde sex hundra sextiosex talenter,
förutom det som infördes genom kringresande handelsmän och andra köpmän; också Arabiens alla konungar och ståthållarna i landet förde guld och silver till Salomo.
Och konung Salomo lät göra två hundra stora sköldar av uthamrat guld och använde till var sådan sköld sex hundra siklar uthamrat guld;
likaledes tre hundra mindre sköldar av uthamrat guld och använde till var sådan sköld tre hundra siklar guld; och konungen satte upp dem i Libanonskogshuset.
Vidare lät konungen göra en stor tron av elfenben och överdrog den med rent guld.
Tronen hade sex trappsteg och en pall av guld, fastsatta vid tronen; på båda sidor om sitsen voro armstöd, och två lejon stodo utmed armstöden;
och tolv lejon stodo där på de sex trappstegen, på båda sidor.
Något sådant har aldrig blivit förfärdigat i något annat rike.
Och alla konung Salomos dryckeskärl voro av guld, och alla kärl i Libanonskogshuset voro av fint guld; silver aktades icke för något i Salomos tid.
Ty konungen hade skepp som gingo till Tarsis med Hurams folk; en gång vart tredje år kommo Tarsis-skeppen hem och förde med sig guld och silver, elfenben, apor och påfåglar.
Och konung Salomo blev större än någon annan konung på jorden, både i rikedom och i vishet.
Alla konungar på jorden kommo för att besöka Salomo och höra den vishet som Gud hade nedlagt i hans hjärta.
Och var och en av dem förde med sig skänker: föremål av silver och av guld, kläder, vapen, välluktande kryddor, hästar och mulåsnor.
Så skedde år efter år.
Och Salomo hade fyra tusen spann hästar med vagnar och tolv tusen ridhästar; dem förlade han dels i vagnsstäderna, dels i Jerusalem, hos konungen själv.
Och han var herre över alla konungar ifrån floden ända till filistéernas land och sedan ända ned till Egyptens gräns.
Och konungen styrde så, att silver blev lika vanligt i Jerusalem som stenar, och cederträ lika vanligt som mullbärsfikonträ i Låglandet.
Och hästar infördes till Salomo från Egypten och från alla andra länder.
Vad nu vidare är att säga om Salomo, om hans första tid såväl som om hans sista, det finnes upptecknat i profeten Natans krönika, i siloniten Ahias profetia och i siaren Jedais syner om Jerobeam, Nebats son.
Salomo regerade i Jerusalem över hela Israel i fyrtio år.
Och Salomo gick till vila hos sina fäder, och man begrov honom i hans fader Davids stad.
Och hans son Rehabeam blev konung efter honom.
Och Rehabeam drog till Sikem, ty hela Israel hade kommit till Sikem för att göra honom till konung.
När Jerobeam, Nebats son, hörde detta, där han var i Egypten -- dit hade han nämligen flytt för konung Salomo -- vände han tillbaka från Egypten.
Och de sände bort och läto kalla honom åter.
Då kom Jerobeam tillstädes jämte hela Israel och talade till Rehabeam och sade:
»Din fader gjorde vårt ok för svårt; men lätta nu du det svåra arbete och det tunga ok som din fader lade på oss, så vilja vi tjäna dig.»
Han svarade dem: »Vänten ännu tre dagar, och kommen så tillbaka till mig.»
Och folket gick.
Då rådförde sig konung Rehabeam med de gamle som hade varit i tjänst hos hans fader Salomo, medan denne ännu levde; han sade: »Vilket svar råden I mig att giva detta folk?»
De svarade honom och sade: »Om du visar dig god mot detta folk och är nådig mot dem och talar goda ord till dem, så skola de för alltid bliva dina tjänare.»
Men han aktade icke på det råd som de gamle hade givit honom, utan rådförde sig med de unga män som hade vuxit upp med honom, och som nu voro i hans tjänst.
Han sade till dem: »Vilket svar råden I oss att giva detta folk som har talat till mig och sagt: 'Lätta det ok som din fader har lagt på oss'?»
De unga männen som hade vuxit upp med honom svarade honom då och sade: »Så bör du säga till folket som har talat till dig och sagt: 'Din fader gjorde vårt ok tungt, men lätta du det för oss' -- så bör du säga till dem: 'Mitt minsta finger är tjockare än min faders länd.
Så veten nu, att om min fader har belastat eder med ett tungt ok, så skall jag göra edert ok ännu tyngre; har min fader tuktat eder med ris, så skall jag göra det med skorpiongissel.'»
Så kom nu Jerobeam med allt folket till Rehabeam på tredje dagen, såsom konungen hade befallt, i det han sade: »Kommen tillbaka till mig på tredje dagen.»
Då gav konungen dem ett hårt svar; ty konung Rehabeam aktade icke på de gamles råd.
Han talade till dem efter de unga männens råd och sade: »Jag skall göra edert ok tungt, ja, jag skall göra det ännu tyngre än förut; har min fader tuktat eder med ris, så skall jag göra det med skorpiongissel.»
Alltså hörde konungen icke på folket; ty det var så skickat av Gud, för att HERRENS ord skulle uppfyllas, det som han hade talat till Jerobeam, Nebats son, genom Ahia från Silo.
Då nu hela Israel förnam att konungen icke ville höra på dem, gav folket konungen detta svar: »Vad del hava vi i David?
Ingen arvslott hava vi i Isais son.
Israel drage hem, var och en till sin hydda.
Se nu själv om ditt hus, du David.»
Därefter drog hela Israel hem till sina hyddor.
Allenast över de israeliter som bodde i Juda städer förblev Rehabeam konung.
Och när konung Rehabeam sände åstad Hadoram, som hade uppsikten över de allmänna arbetena, stenade Israels barn denne till döds; och konung Rehabeam själv måste med hast stiga upp i sin vagn och fly till Jerusalem.
Så avföll Israel från Davids hus och har varit skilt därifrån ända till denna dag.
Och när Rehabeam kom till Jerusalem, församlade han Juda hus och Benjamin, ett hundra åttio tusen utvalda krigare, för att de skulle strida mot Israel och återvinna konungadömet åt Rehabeam.
Men HERRENS ord kom till gudsmannen Semaja; han sade:
»Säg till Rehabeam, Salomos son, Juda konung, och till alla israeliter i Juda och Benjamin:
Så säger HERREN: I skolen icke draga upp och strida mot edra bröder.
Vänden tillbaka hem, var och en till sitt, ty vad som har skett har kommit från mig.»
Och de lyssnade till HERRENS ord och vände om och drogo icke mot Jerobeam.
Men Rehabeam bodde i Jerusalem, och han befäste städer i Juda och gjorde dem till fasta platser.
Han befäste Bet-Lehem, Etam, Tekoa,
Bet-Sur, Soko, Adullam
Gat, Maresa, Sif,
Adoraim, Lakis, Aseka,
Sorga, Ajalon och Hebron, alla i Juda och Benjamin, och gjorde dem till fasta städer.
Och han gjorde deras befästningar starka och tillsatte hövdingar i dem och lade in i dem förråd av mat, olja och vin;
var och en särskild av dessa städer försåg han med sköldar och spjut; han befäste dem mycket starkt.
Och Juda och Benjamin förblevo under hans välde.
Och prästerna och leviterna i hela Israel gingo över till honom från alla sina områden;
ty leviterna övergåvo sina utmarker och sina andra besittningar och begåvo sig till Juda och Jerusalem, eftersom Jerobeam med sina söner drev dem bort ifrån deras tjänst såsom HERRENS präster,
och anställde åt sig andra präster för offerhöjderna och för de onda andarna och för kalvarna som han hade låtit göra.
Och dem följde ifrån alla Israels stammar de som vände sina hjärtan till att söka HERREN, Israels Gud; dessa kommo till Jerusalem för att offra åt HERREN, sina fäders Gud.
I tre år befäste de så konungamakten i Juda och gjorde Rehabeams, Salomos sons, välde starkt; ty i tre år vandrade de på Davids och Salomos väg.
Och Rehabeam tog till hustru åt sig Mahalat, dotter till Jerimot, Davids son, och till Abihail, Eliabs, Isais sons, dotter.
Hon födde åt honom sönerna Jeus, Semarja och Saham.
Och efter henne tog han till hustru Maaka, Absaloms dotter.
Hon födde åt honom Abia, Attai, Sisa och Selomit.
Och Rehabeam hade Maaka, Absaloms dotter, kärare än alla sina andra hustrur och bihustrur -- ty han hade tagit aderton hustrur och sextio bihustrur -- och han födde tjuguåtta söner och sextio döttrar.
Och Rehabeam satte Abia, Maakas son, till huvud och furste bland sina bröder, ty han hade i sinnet att göra honom till konung.
Och på lämpligt sätt fördelade han alla Judas och Benjamins landskap och alla fasta städer mellan några av sina söner och gav dem rikligt underhåll; han skaffade dem ock hustrur i mängd.
När Rehabeams konungamakt nu hade blivit befäst och han hade blivit mäktig, övergav han HERRENS lag, han jämte hela Israel.
Men i konung Rehabeams femte regeringsår drog Sisak, konungen i Egypten, upp mot Jerusalem, därför att de hade varit otrogna mot HERREN;
han kom med ett tusen två hundra vagnar och sextio tusen ryttare, och ingen kunde räkna det folk som följde honom från Egypten: libyer, suckéer och etiopier.
Och han intog de fasta städerna i Juda och kom ända till Jerusalem.
Och profeten Semaja hade kommit till Rehabeam och till Juda furstar, som hade församlat sig i Jerusalem av fruktan för Sisak; och han sade till dem: »Så säger HERREN: I haven övergivit mig, därför har ock jag övergivit eder och givit eder i Sisaks hand.»
Då ödmjukade sig Israels furstar och konungen själv och sade: »HERREN är rättfärdig.»
När nu HERREN såg att de ödmjukade sig, kom HERRENS ord till Semaja; han sade: »Eftersom de hava ödmjukat sig, vill jag icke fördärva dem; jag skall låta dem med knapp nöd komma undan, och min vrede skall icke bliva utgjuten över Jerusalem genom Sisaks hand.
Dock skola de nödgas bliva honom underdåniga, för att de må lära sig förstå vilken skillnad det är mellan att tjäna mig och att tjäna främmande konungadömen.»
Så drog nu Sisak, konungen i Egypten, upp mot Jerusalem.
Och han tog skatterna i HERRENS hus och skatterna i konungshuset; alltsammans tog han.
Han tog ock de gyllene sköldar som Salomo hade låtit göra.
I deras ställe lät konung Rehabeam göra sköldar av koppar, och dessa lämnade han i förvar åt hövitsmännen för drabanterna som höllo vakt vid ingången till konungshuset.
Och så ofta konungen gick till HERRENS hus, gingo ock drabanterna och buro dem; sedan förde de dem tillbaka till drabantsalen.
Därför att nu Rehabeam ödmjukade sig, vände sig HERRENS vrede ifrån honom, så att han icke alldeles fördärvade honom.
Också fanns ännu något gott i Juda.
Alltså befäste konung Rehabeam sitt välde i Jerusalem och fortsatte att regera.
Rehabeam var nämligen fyrtioett år gammal, när han blev konung, och han regerade sjutton år i Jerusalem, den stad som HERREN hade utvalt ur alla Israel stammar, till att där fästa sitt namn.
Hans moder hette Naama, ammonitiskan.
Och han gjorde vad ont var, ty han vände icke sitt hjärta till att söka HERREN.
Men vad som är att säga om Rehabeam, om hans första tid såväl som om hans sista, det finnes upptecknat i profeten Semajas och siaren Iddos krönikor, enligt släktregistrens sätt.
Och Rehabeam och Jerobeam lågo i krig med varandra, så länge de levde.
Men Rehabeam gick till vila hos sina fäder och blev begraven i Davids stad.
Och hans son Abia blev konung efter honom.
I konung Jerobeams adertonde regeringsår blev Abia konung över Juda.
Han regerade tre år i Jerusalem.
Hans moder hette Mikaja, Uriels dotter, från Gibea.
Men Abia och Jerobeam lågo i krig med varandra.
Och Abia begynte kriget med en här av tappra krigsmän, fyra hundra tusen utvalda män; men Jerobeam ställde upp sig till strid mot honom med åtta hundra tusen utvalda tappra stridsmän.
Och Abia steg upp på berget Semaraim i Efraims bergsbygd och sade: »Hören mig, du, Jerobeam, och I, hela Israel.
Skullen I icke veta att det är HERREN, Israels Gud, som har givit åt David konungadömet över Israel för evig tid, åt honom själv och hans söner, genom ett saltförbund?
Men Jerobeam, Nebats son, Salomos, Davids sons, tjänare, uppreste sig och avföll från sin herre.
Och till honom församlade sig löst folk, onda män, och de blevo Rehabeam, Salomos son, för starka, eftersom Rehabeam ännu var ung och försagd och därför icke kunde stå dem emot.
Och nu menen I eder kunna stå emot HERRENS konungadöme, som tillhör Davids söner, eftersom I ären en stor hop och haven hos eder de guldkalvar som Jerobeam har låtit göra åt eder till gudar.
Haven I icke fördrivit HERRENS präster, Arons söner, och leviterna, och själva gjort eder präster, såsom de främmande folken göra?
Vemhelst som kommer med en ungtjur och sju vädurar for att taga handfyllning, han får bliva präst åt dessa gudar, som icke äro gudar.
Men vi hava HERREN till vår Gud, och vi hava icke övergivit honom.
Vi hava präster av Arons söner, som göra tjänst inför HERREN, och leviter, som sköta tempelsysslorna;
och de förbränna åt HERREN brännoffer var morgon och var afton och antända välluktande rökelse och lägga upp bröd på det gyllene bordet och tända var afton den gyllene ljusstaken med dess lampor.
Ty vi hålla vad HERREN, vår Gud, har bjudit oss hålla, men I haven övergivit honom.
Och se, vi hava Gud i spetsen för oss, och vi hava hans präster med larmtrumpeterna för att blåsa till strid mot eder.
I Israels barn, striden icke mot HERREN, edra fäders Gud; ty då skall det icke gå eder väl.»
Men Jerobeam hade låtit kringgå dem och lagt ett bakhåll för att falla dem i ryggen; så stodo de nu mitt emot Juda män och hade sitt bakhåll bakom dem.
När då Juda män vände sig om, fingo de se att de hade fiender både framför sig och bakom sig.
Då ropade de till HERREN, och prästerna blåste i trumpeterna.
Därefter hovo Juda män upp ett härskri; och när Juda män hovo upp sitt härskri, lät Gud Jerobeam och hela Israel bliva slagna av Abia och Juda.
Och Israels barn flydde för Juda, och Gud gav dem i deras hand.
Och Abia med sitt folk anställde ett stort nederlag bland dem, så att fem hundra tusen unga män av Israel föllo slagna.
Alltså blevo Israels barn på den tiden kuvade; men Juda barn voro starka, ty de stödde sig på HERREN sina fäders Gud.
Och Abia förföljde Jerobeam och tog ifrån honom några städer: Betel med underlydande orter, Jesana med underlydande orter och Efron med underlydande orter.
Och Jerobeam förmådde ingenting mer, så länge Abia levde; och han blev hemsökt av HERREN, så att han dog.
Men Abia befäste sitt välde; och han tog sig fjorton hustrur och födde tjugutvå söner och sexton döttrar.
Vad nu mer är att säga om Abia, om hans företag och om annat som rör honom, det finnes upptecknat i profeten Iddos »Utläggning».
Och Abia gick till vila hos sina fäder, och man begrov honom i Davids stad.
Och hans son Asa blev konung efter honom.
Under hans tid hade landet ro i tio år.
Och Asa gjorde vad gott och rätt var i HERRENS, sin Guds, ögon.
Han skaffade bort de främmande altarna och offerhöjderna och slog sönder stoderna och högg ned Aserorna.
Och han uppmanade Juda att söka HERREN, sina fäders Gud, och hålla lagen och budorden.
Ur alla Juda städer skaffade han bort offerhöjderna och solstoderna; och riket hade ro under honom.
Och han byggde fasta städer i Juda, eftersom landet hade ro och han under dessa år icke hade något krig; ty HERREN hade givit honom lugn.
Han sade nämligen till Juda: »Låt oss bygga dessa städer och förse dem runt omkring med murar och torn, med portar och bommar, medan vi ännu hava landet i vår makt, därför att vi hava sökt HERREN, vår Gud; ty vi hava sökt honom, och han har låtit oss få lugn på alla sidor.»
Så byggde de då, och allt gick väl.
Och Asa hade en här som var väpnad med stora sköldar och med spjut, och som utgjordes av tre hundra tusen man från Juda, vartill kommo två hundra åttio tusen man från Benjamin, som voro väpnade med små sköldar och spände båge.
Alla dessa voro tappra stridsmän.
Men Sera från Etiopien drog ut mot dem med en här av tusen gånger tusen man och tre hundra vagnar; och han kom till Maresa.
Och Asa drog ut mot honom, och de ställde upp sig till strid i Sefatas dal vid Maresa.
Och Asa ropade till HERREN, sin Gud, och sade: »HERRE, förutom dig finnes ingen som kan hjälpa i striden mellan den starke och den svage.
Så hjälp oss, HERRE, vår Gud, ty på dig stödja vi oss, och i ditt namn hava vi kommit hit mot denna hop.
HERRE, du är vår Gud; mot dig förmår ju ingen människa något.»
Och HERREN lät etiopierna bliva slagna av Asa och Juda, så att etiopierna flydde.
Och Asa och hans folk förföljde dem ända till Gerar; och av etiopierna föllo så många, att ingen av dem kom undan med livet, ty de blevo nedgjorda av HERREN och hans här.
Och folket tog byte i stor myckenhet.
Och de intogo alla städer runt omkring Gerar, ty en förskräckelse ifrån HERREN hade kommit över dessa; och de plundrade alla städerna, ty i dem fanns mycket att plundra.
Till och med boskapsskjulen bröto de ned och förde bort småboskap i myckenhet och kameler, och vände så tillbaka till Jerusalem.
Och över Asarja, Odeds son, kom Guds Ande.
Han gick ut mot Asa och sade till honom: »Hören mig, du, Asa, och I, hela Juda och Benjamin.
HERREN är med eder, när I ären med honom, och om I söken honom, så låter han sig finnas av eder; men om I övergiven honom, så övergiver han ock eder.
En lång tid var ju Israel utan den sanne Guden, utan präster som undervisade dem, och utan någon lag.
Men i sin nöd omvände de sig till HERREN, Israels Gud, och när de sökte honom, lät han sig finnas av dem.
Under de tiderna fanns ingen trygghet, när man gick ut eller in; utan stor förvirring rådde bland alla dem som bodde här i länderna,
och folk drabbade samman med folk och stad med stad; ty Gud förvirrade dem med allt slags nöd.
Men varen I frimodiga, låten icke modet falla, ty edert verk skall få sin lön.»
När Asa hörde dessa ord och denna profetia av profeten Oded, tog han mod till sig och skaffade bort styggelserna ur Judas och Benjamins hela land och ur de städer som han hade tagit i Efraims bergsbygd, och upprättade åter HERRENS altare, det som stod framför HERRENS förhus.
Och han församlade hela Juda och Benjamin, så ock de främlingar ifrån Efraim, Manasse och Simeon, som bodde ibland dem; ty många från Israel hade gått över till honom, när de sågo att HERREN, hans Gud, var med honom.
Och de församlade sig till Jerusalem i tredje månaden av Asas femtonde regeringsår,
och offrade på den dagen åt HERREN sju hundra tjurar och sju tusen djur av småboskapen, uttagna av det byte som de hade fört med sig.
Och de ingingo det förbundet att de skulle söka HERREN, sina fäders Gud, av allt sitt hjärta och av all sin själ,
och att var och en som icke sökte HERREN, Israels Gud, han skulle bliva dödad, liten eller stor, man eller kvinna.
Och de gåvo HERREN sin ed med hög röst och under jubel, och under det att trumpeter och basuner ljödo.
Och hela Juda gladde sig över eden; ty de hade svurit den av allt sitt hjärta, och de sökte HERREN med hela sin vilja, och han lät sig finnas av dem, och han lät dem få ro på alla sidor.
Konung Asa avsatte ock sin moder Maaka från hennes drottningsvärdighet, därför att hon hade satt upp en styggelse åt Aseran; Asa högg nu ned styggelsen och krossade de och brände upp den i Kidrons dal.
Men offerhöjderna blevo icke avskaffade ur Israel; dock var Asas hjärta gudhängivet, så länge han levde.
Och han förde in i Guds hus både vad hans fader och vad han själv hade helgat åt HERREN: silver, guld och kärl.
Och intet krig uppstod förrän i Asas trettiofemte regeringsår.
I Asas trettiosjätte regeringsår drog Baesa, Israels konung, upp mot Juda och begynte befästa Rama, för att hindra att någon komme vare sig från eller till Asa, Juda konung.
Då tog Asa silver och guld ur skattkamrarna i HERRENS hus och i konungshuset, och sände det till Ben-Hadad, konungen i Aram, som bodde i Damaskus, och lät säga:
»Ett förbund består ju mellan mig och dig, såsom det var mellan min fader och din fader.
Se, här sänder jag dig silver och guld; så bryt då ditt förbund med Baesa, Israels konung, för att han må lämna mig i fred.»
Och Ben-Hadad lyssnade till konung Asa och sände sina krigshövitsmän mot Israels städer, och de förhärjade Ijon, Dan och Abel-Maim samt alla förrådshus i Naftali städer.
När Baesa hörde detta, avstod han från att befästa Rama och lät sina arbeten där upphöra.
Men konung Asa tog med sig hela Juda, och de förde bort ifrån Rama stenar och trävirke som Baesa använde till att befästa det.
Därmed befäste han så Geba och Mispa.
Vid samma tid kom siaren Hanani till Asa, Juda konung, och sade till honom: »Eftersom du stödde dig på konungen i Aram och icke stödde dig på HERREN, din Gud, därför har den arameiske konungens här sluppit undan din hand.
Voro icke etiopierna och libyerna en väldig här, med vagnar och ryttare i stor myckenhet?
Men därför att du då stödde dig på HERREN, gav han dem i din hand.
TY HERRENS ögon överfara hela jorden, för att han med sin kraft skall bistå dem som med sina hjärtan hängiva sig åt honom.
Härutinnan har du handlat dåraktigt.
Därför skall du hädanefter hava ständiga strider.»
Men Asa blev förtörnad på siaren och satte honom i stockhuset; så förbittrad var han på honom för vad han hade sagt.
Vid samma tid förfor Asa ock våldsamt mot andra av folket.
Men vad som är att säga om Asa, om hans första tid såväl som om hans sista, det finnes upptecknat i boken om Judas och Israels konungar.
Och i sitt trettionionde regeringsår fick Asa en sjukdom i sina fötter, och sjukdomen blev övermåttan svår; men oaktat sin sjukdom sökte han icke HERREN, utan allenast läkares hjälp.
Och Asa gick till vila hos sina fäder och dog i sitt fyrtioförsta regeringsår.
Och man begrov honom i den grav som han hade låtit hugga ut åt sig i Davids stad; och man lade honom på en bädd som man hade fyllt med vällukter och kryddor av olika slag, konstmässigt beredda, och anställde till hans ära en mycket stor förbränning.
Och hans son Josafat blev konung; efter honom.
Han befäste sitt välde mot Israel.
Han lade in krigsfolk i alla Juda fasta städer och lade in besättningar i Juda land och i de Efraims städer som hans fader Asa hade intagit.
Och HERREN var med Josafat, ty han vandrade på sin fader Davids första vägar och sökte icke Baalerna,
utan sökte sin faders Gud och vandrade efter hans bud och gjorde icke såsom Israel.
Därför befäste HERREN konungadömet i hans hand, och hela Juda gav skänker åt Josafat, så att hans rikedom och ära blev stor.
Och då hans frimodighet växte på HERRENS vägar, skaffade han också bort offerhöjderna och Aserorna ur Juda.
Och i sitt tredje regeringsår sände han ut sina hövdingar Ben-Hail, Obadja, Sakarja, Netanel och Mikaja, till att undervisa i Juda städer,
och med dem några leviter, nämligen leviterna Semaja, Netanja, Sebadja, Asael, Semiramot, Jonatan, Adonia, Tobia och Tob-Adonia; och de hade med sig prästerna Elisama och Joram.
Dessa undervisade nu i Juda och hade HERRENS lagbok med sig; de foro omkring i alla Juda städer och undervisade bland folket.
Och en förskräckelse ifrån HERREN kom över alla riken i de länder som lågo omkring Juda, så att de icke vågade kriga mot Josafat.
Och en del av filistéerna förde skänker till Josafat och gåvo silver i skatt.
Därtill förde ock araberna till honom småboskap, sju tusen sju hundra vädurar och sju tusen sju undra bockar.
Så blev Josafat allt mäktigare och till slut övermåttan mäktig.
Och han byggde borgar och förrådsstäder i Juda.
Han hade stora upplag i Juda städer; och krigsfolk, tappra stridsmän, hade han i Jerusalem.
Och detta var ordningen bland dem, efter deras familjer.
Till Juda hörde följande överhövitsmän: hövitsmannen Adna och med honom tre hundra tusen tappra stridsmän;
därnäst hövitsmannen Johanan och med honom två hundra åttio tusen;
därnäst Amasja, Sikris son, som frivilligt hade givit sig i HERRENS tjänst, och med honom två hundra tusen tappra stridsmän.
Men från Benjamin voro: Eljada, en tapper stridsman, och med honom två hundra tusen, väpnade med båge och sköld;
därnäst Josabad och med honom ett hundra åttio tusen, rustade till strid.
Dessa voro de som gjorde tjänst hos konungen; därtill kommo de som konungen hade förlagt i de befästa städerna i hela Juda.
När Josafat nu hade kommit till stor rikedom och ära, befryndade han sig med Ahab.
Och efter några års förlopp for han ned till Ahab i Samaria.
Och Ahab lät för honom och folket som han hade med sig slakta får och fäkreatur i myckenhet; och han sökte intala honom att draga upp mot Ramot i Gilead.
Ahab, Israels konung, frågade alltså Josafat, Juda konung: »Vill du draga med mig mot Ramot i Gilead?»
Han svarade honom: »Jag såsom du, och mitt folk såsom ditt folk!
Jag vill följa med dig i striden.»
Men Josafat sade ytterligare till Israels konung: »Fråga dock först HERREN härom.»
Då församlade Israels konung profeterna, fyra hundra män, och frågade dem: »Skola vi draga åstad till Ramot i Gilead för att belägra det, eller skall jag avstå därifrån?»
De svarade: »Drag ditupp; Gud skall giva det i konungens hand.»
Men Josafat sade: »Finnes här ingen annan HERRENS profet, så att vi kunna fråga genom honom?»
Israels konung svarade Josafat: »Här finnes ännu en man, Mika, Jimlas son, genom vilken vi kunna fråga HERREN; men han är mig förhatlig, ty han profeterar aldrig lycka åt mig, utan beständigt allenast olycka.»
Josafat sade: »Konungen säge icke så.»
Då kallade Israels konung till sig en hovman och sade: »Skaffa skyndsamt hit Mika, Jimlas son.»
Israels konung och Josafat, Juda konung, sutto nu var och en på sin tron, iklädda sina skrudar; de sutto på en tröskplats vid Samarias port, under det att alla profeterna profeterade inför dem.
Då gjorde sig Sidkia, Kenaanas son, horn av järn och sade: »Så säger HERREN: Med dessa skall du stånga araméerna, så att de förgöras.»
Och alla profeterna profeterade på samma sätt och sade: »Drag upp mot Ramot i Gilead, så skall du bliva lyckosam; HERREN skall giva det i konungens hand.»
Och budet som hade gått för att kalla på Mika talade till honom och sade: »Det är så, att profeterna med en mun lova konungen lycka; så låt nu ock ditt tal stämma överens med deras, och lova också du lycka.»
Men Mika svarade: »Så sant HERREN lever, jag skall allenast tala det som min Gud säger.»
När han sedan kom till konungen, frågade konungen honom: »Mika, skola vi draga åstad till Ramot i Gilead för att belägra det, eller skall jag avstå därifrån?»
Han svarade: »Dragen ditupp, så skolen I bliva lyckosamma; de skola bliva givna i eder hand.»
Men konungen sade till honom: »Huru många gånger skall jag besvärja dig att icke tala till mig annat än sanning i HERRENS namn?»
Då sade han: »Jag såg hela Israel förskingrat på bergen, likt får som icke hava någon herde.
Och HERREN sade: 'Dessa hava icke någon herre; må de vända tillbaka hem i frid, var och en till sitt.'»
Då sade Israels konung till Josafat: »Sade jag dig icke att denne aldrig profeterar lycka åt mig, utan allenast olycka?»
Men han sade: »Hören alltså HERRENS ord.
Jag såg HERREN sitta på sin tron och himmelens hela härskara stå på hans högra sida och på hans vänstra.
Och HERREN sade: 'Vem vill locka Ahab, Israels konung, att draga upp mot Ramot i Gilead, för att han må falla där?'
Då sade den ene så och den andre så.
Slutligen kom anden fram och ställde sig inför HERREN och sade: 'Jag vill locka honom därtill.'
HERREN frågade honom: 'På vad sätt?'
Han svarade: 'Jag vill gå ut och bliva en lögnens ande i alla hans profeters mun.»
Då sade han: 'Du må försöka att locka honom därtill och du skall också lyckas; gå ut och gör så.'
Och se, nu har HERREN lagt en lögnens ande i dessa dina profeters mun, medan HERREN ändå har beslutit att olycka skall komma över dig.»
Då trädde Sidkia, Kenaanas son, fram och gav Mika ett slag på kinden och sade: »På vilken väg har då HERRENS Ande gått bort ifrån mig för att tala med dig?»
Mika svarade: »Du skall få se det på den dag då du nödgas springa från kammare till kammare för att gömma dig.»
Men Israels konung sade: »Tagen Mika och fören honom tillbaka till Amon, hövitsmannen i staden, och till Joas, konungasonen.
Och sägen: Så säger konungen: Sätten denne i fängelse och bespisen honom med fångkost, till dess jag kommer välbehållen tillbaka.»
Mika svarade: »Om du kommer välbehållen tillbaka, så har HERREN icke talat genom mig.»
Och han sade ytterligare: »Hören detta, I folk, allasammans.»
Så drog nu Israels konung jämte Josafat, Juda konung, upp till Ramot i Gilead.
Och Israels konung sade till Josafat: »Jag vill förkläda mig, när jag drager ut i striden, men du må vara klädd i dina egna kläder.»
Så förklädde sig Israels konung, när de drogo ut i striden.
Men konungen i Aram hade bjudit och sagt till sina vagnshövitsmän: »I skolen icke giva eder i strid med någon, vare sig liten eller stor, utom med Israels konung allena.»
När då hövitsmannen över vagnarna fingo se Josafat, tänkte de: »Detta är Israels konung», och omringade honom därför, i avsikt att anfalla honom.
Då gav Josafat upp ett rop, och HERREN hjälpte honom, Gud vände dem bort ifrån honom.
Så snart nämligen hövitsmännen över vagnarna märkte att det icke var Israels konung, vände de om och läto honom vara.
Men en man som spände sin båge och sköt på måfå träffade Israels konung i en fog på rustningen.
Då sade denne till sin körsven: »Sväng om vagnen och för mig ut ur hären, ty jag är sårad.»
Och striden blev på den dagen allt häftigare, och Israels konung höll sig ända till aftonen upprätt i sin vagn, vänd mot araméerna; men vid den tid då solen gick ned gav han upp andan.
Men Josafat, Juda konung, vände välbehållen hem igen till Jerusalem.
Då gick siaren Jehu, Hananis son, ut mot konung Josafat och sade till honom: »Skall man då hjälpa den ogudaktige?
Skall du då älska dem som hata HERREN?
För vad du har gjort vilar nu HERRENS förtörnelse över dig.
Dock har något gott blivit funnet hos dig, ty du har utrotat Aserorna ur landet och har vänt ditt hjärta till att söka Gud.»
Och Josafat stannade nu i Jerusalem, men sedan drog han åter ut bland folket, ifrån Beer-Seba ända till Efraims bergsbygd, och förde dem tillbaka till HERREN, deras fäders Gud.
Och han anställde domare i landet, i alla Juda befästa städer, särskilda för var stad.
Och han sade till dessa domare: »Sen till, vad I gören; ty I dömen icke människodom, utan HERRENS dom, och han är närvarande, så ofta I dömen.
Låten alltså nu fruktan för HERREN vara över eder.
Given akt på vad I gören; ty hos HERREN, vår Gud, finnes ingen orätt, och han har icke anseende till personen, ej heller tager han mutor.»
Också i Jerusalem hade Josafat anställt några av leviterna och prästerna och några av huvudmännen för Israels familjer till att döma HERRENS dom och avgöra rättstvister.
När de sedan vände tillbaka till Jerusalem,
bjöd han dem och sade: »Så skolen I göra i HERRENS fruktan, redligt och med hängivet hjärta.
Och så ofta någon rättssak drages inför eder av edra bröder, som bo i sina städer, det må gälla dom i en blodssak eller eljest tillämpning av lag och bud, stadgar och rätter, då skolen I varna dem, så att de icke ådraga sig skuld inför HERREN, varigenom förtörnelse kommer över eder och edra bröder.
Så skolen I göra, för att I icke mån ådraga eder skuld.
Och se, översteprästen Amarja skall vara eder förman i alla HERRENS saker, och Sebadja, Ismaels son, fursten för Juda hus, i alla konungens saker; och leviterna skola vara tillsyningsmän under eder.
Varen nu ståndaktiga i vad I gören, och HERREN skall vara med den som är god.»
Därefter kommo Moabs barn och Ammons barn och med dem en del av ammoniterna för att strida mot Josafat.
Och man kom och berättade detta för Josafat och sade: »En stor hop kommer mot dig från landet på andra sidan havet, från Aram, och de äro redan i Hasason-Tamar (det är En-Gedi).»
Då blev Josafat förskräckt och vände sin håg till att söka HERREN; och han lät lysa ut en fasta över hela Juda.
Och Juda församlade sig för att söka hjälp hos HERREN; ja, från alla Juda städer kom man för att söka HERREN.
Och Josafat trädde upp i Juda mäns och Jerusalems församling i HERRENS hus, framför den nya förgården,
och sade: »HERRE, våra fäders Gud, är icke du Gud i himmelen och den som råder över alla hednafolkens riken?
I din hand är kraft och makt; och ingen finnes, som kan stå dig emot.
Var det icke du, vår Gud, som fördrev detta lands inbyggare för ditt folk Israel och gav det åt Abrahams, din väns, säd för evig tid?
De fingo bo där, och de byggde dig där en helgedom åt ditt namn, i det de sade:
'Om något ont kommer över oss, svärd, straffdom eller pest eller hungersnöd, så vilja vi träda upp inför detta hus och inför dig, ty ditt namn är i detta hus; och vi vilja ropa till dig i vår nöd, och du skall då höra och hjälpa.'
Se därför nu huru Ammons barn och Moab och folket i Seirs bergsbygd -- genom vilkas område du icke tillstadde Israel att gå, när de kommo från Egyptens land, varför de ock togo en omväg bort ifrån dem och icke förgjorde dem --
se huru dessa nu vedergälla oss, i det att de komma för att förjaga oss ur det land som är din besittning, och som du har givit oss till besittning.
Du, vår Gud, skall du icke hålla dom över dem?
Ty vi förmå intet mot denna stora hop som kommer emot oss, och själva veta vi icke vad vi skola göra, utan till dig se våra ögon.»
Och hela Juda stod där inför HERREN med sina späda barn, sina hustrur och söner.
Då kom HERRENS Ande mitt i församlingen över Jahasiel, son till Sakarja, son till Benaja, son till Jegiel, son till Mattanja, en levit, av Asafs söner,
och han sade: »Akten härpå, alla I av Juda, och I Jerusalems invånare, och du konung Josafat.
Så säger HERREN till eder: Frukten icke och varen icke förfärade för denna stora hop, ty striden är icke eder, utan Guds.
Dragen i morgon ned mot dem.
De draga då upp på Hassishöjden, och I skolen träffa dem vid andan av dalen, framför Jeruels öken.
Men därvid bliver det icke eder sak att strida.
I skolen allenast träda fram och stå stilla och se på, huru HERREN frälsar eder, I av Juda och Jerusalem.
Frukten icke och varen icke förfärade.
Dragen i morgon ut mot dem, och HERREN skall vara med eder.»
Då böjde Josafat sig ned med ansiktet mot jorden, och alla Juda män och Jerusalems invånare föllo ned för HERREN och tillbådo HERREN.
Och de av leviterna, som tillhörde kehatiternas och koraiternas barn, stodo upp och lovade HERREN, Israels Gud, med hög och stark röst.
Men bittida följande morgon drogo de ut till Tekoas öken.
Och när de drogo ut, trädde Josafat fram och sade: »Hören mig, I av Juda och I Jerusalems invånare.
Haven tro på HERREN, eder Gud, så skolen I hava ro.
Och tron på hans profeter, så skolen I bliva lyckosamma.»
Och sedan han hade rådfört sig med folket, ställde han upp män som skulle sjunga till HERRENS ära och lova honom i helig skrud, under det att de drogo ut framför den väpnade hären; de skulle sjunga: »Tacken HERREN, ty hans nåd varar evinnerligen.»
Och just som de begynte med sången och lovet, lät HERREN ett angrepp ske bakifrån på Ammons barn och Moab och folket ifrån Seirs bergsbygd, dem som hade kommit mot Juda; och de blevo slagna.
Och Ammons barn och Moab reste sig mot folket ifrån Seirs bergsbygd och gåvo dem till spillo och förgjorde dem; och när de hade gjort ände på folket ifrån Seir, hjälptes de åt att nedgöra varandra.
När sedan Juda män kommo upp på höjden, varifrån man kunde se ut över öknen, och vände sig mot fiendernas hop, fingo de se dessa ligga döda på jorden, och ingen hade undkommit.
Och när Josafat begav sig dit med sitt folk för att plundra och taga byte från dem, funno de där en myckenhet av gods och av döda kroppar och av dyrbara ting; och de togo for sig så mycket att de icke kunde bära det.
Och de fortsatte plundringen i tre dagar; så stort var bytet.
Men på fjärde dagen församlade de sig i Berakadalen; där lovade de HERREN, och därav fick det stället namnet Berakadalen , såsom det heter ännu i dag.
Därefter vände alla Judas och Jerusalems män, med Josafat i spetsen, glada tillbaka igen till Jerusalem; ty HERREN hade berett dem glädje genom vad som hade skett med deras fiender.
Och de drogo in i Jerusalem med psaltare, harpor och trumpeter och tågade till HERRENS hus.
Och en förskräckelse ifrån Gud kom över alla de främmande rikena, när de hörde att HERREN hade stritt mot Israels fiender.
Och Josafats rike hade nu ro, ty hans Gud lät honom få lugn på alla sidor.
Så regerade Josafat över Juda. han var trettiofem år gammal, när han blev konung, och han regerade tjugufem år i Jerusalem.
Hans moder hette Asuba, Silhis dotter.
Och han vandrade på sin fader Asas väg, utan att vika av ifrån den; han gjorde nämligen vad rätt var i HERRENS ögon.
Dock blevo offerhöjderna icke avskaffade, och ännu hade folket icke vänt sina hjärtan till sina fäders Gud.
Vad nu mer är att säga om Josafat, om hans första tid såväl som om hans sista, det finnes upptecknat i Jehus, Hananis sons, krönika, som är upptagen i boken om Israels konungar.
Men sedan förband sig Josafat, Juda konung, med Ahasja, Israels konung, fastän denne var ogudaktig i sina gärningar;
han förband sig med honom för att bygga skepp som skulle gå till Tarsis.
Och de byggde skepp i Esjon-Geber.
Då profeterade Elieser, Dodavahus son, från Maresa, mot Josafat; han sade: »Därför att du har förbundit dig med Ahasja, skall HERREN låta ditt företag bliva om intet.»
Och somliga av skeppen ledo skeppsbrott, så att de icke kunde gå till Tarsis.
Och Josafat gick till vila hos sina fäder och blev begraven hos sina fäder i Davids stad.
Och hans son Joram blev konung efter honom.
Denne hade bröder, söner till Josafat: Asarja, Jehiel, Sakarja, Asarjahu, Mikael och Sefatja; alla dessa voro söner till Josafat, Israels konung.
Och deras fader gav dem stora skänker i silver och guld och dyrbarheter, därtill ock fasta städer i Juda; men konungadömet hade han givit åt Joram, ty denne var den förstfödde.
När Joram nu hade övertagit sin faders konungadöme och befäst sig däri, dräpte han alla sina bröder med svärd, så ock några av Israels furstar,
Joram var trettiotvå år gammal, är han blev konung, och han regerade åtta år i Jerusalem.
Men han vandrade på Israels konungars väg, såsom Ahabs hus hade gjort, ty en dotter till Ahab var hans hustru; han gjorde vad ont var i HERRENS ögon.
Dock ville HERREN icke fördärva Davids hus, för det förbunds skull som han hade slutit med David, och enligt sitt löfte, att han skulle låta honom och hans söner hava en lampa för alltid.
I hans tid avföll Edom från Juda välde och satte en egen konung över sig.
Då drog Joram dit med sina hövitsmän och med alla sina stridsvagnar.
Och om natten gjorde han ett anfall på edoméerna, som hade omringat honom, och slog dem och hövitsmännen över deras vagnar.
Så avföll Edom från Juda välde, och det har varit skilt därifrån ända till denna dag.
Vid samma tid avföll ock Libna från hans välde, därför att han hade övergivit HERREN, sina fäders Gud.
Också han uppförde offerhöjder på bergen i Juda och förledde så Jerusalems invånare till trolös avfällighet och förförde Juda.
Men en skrivelse kom honom till handa från profeten Elia, så lydande: »Så säger HERREN, din fader Davids Gud: Se, du har icke vandrat på din fader Josafats vägar eller på Asas, Juda konungs, vägar,
utan du har vandrat på Israels konungars väg och förlett Juda och Jerusalems invånare till trolös avfällighet, på samma sätt som Ahabs hus förledde till avfällighet; du har också dräpt dina bröder, dem som hörde till din faders hus, och som voro bättre än du.
Därför skall HERREN låta en stor hemsökelse drabba ditt folk, så ock dina barn och dina hustrur och allt vad du äger;
och själv skall du träffas av svår sjukdom, en sjukdom i dina inälvor, så svår att dina inälvor, efter år och dagar, skola falla ut i följd av sjukdomen.»
Och HERREN uppväckte mot Joram filistéernas ande och de arabers som bodde närmast etiopierna;
och de drogo upp mot Juda och bröto in där och förde bort allt gods som fanns i konungens hus, därtill ock hans söner och hustrur, så att han icke hade kvar någon av sina söner förutom Joahas, sin yngste son.
Och efter allt detta hemsökte HERREN honom med en obotlig sjukdom i inälvorna.
Och efter år och dagar, när två år voro förlidna, föllo hans inälvor ut i följd av sjukdomen, och han dog i svåra plågor; men hans folk anställde ingen förbränning till hans ära, såsom de hade gjort efter hans fäder.
Han var trettiotvå år gammal, när han blev konung, och han regerade åtta år i Jerusalem.
Och han gick bort utan att bliva saknad, och man begrov honom i Davids stad, men icke i konungagravarna.
Och Jerusalems invånare gjorde Ahasja, hans yngste son, till konung efter honom; ty alla de äldre hade blivit dräpta av den rövarskara som med araberna hade kommit till lägret.
Så blev då Ahasja, Jorams son, konung i Juda.
Fyrtiotvå år gammal var Ahasja, är han blev konung, ock han regerade ett år i Jerusalem.
Hans moder hette Atalja, Omris dotter.
Också han vandrade på Ahabs hus' vägar, ty hans moder var hans rådgiverska i ogudaktighet.
Han gjorde vad ont var i HERRENS ögon likasom Ahabs hus; ty därifrån tog han, efter sin faders död, sina rådgivare, till sitt eget fördärv.
Det var ock deras råd han följde, när han drog åstad med Joram, Ahabs son, Israels konung, och stridde mot Hasael, konungen i Aram, vid Ramot i Gilead.
Men Joram blev sårad av araméerna.
Då vände han tillbaka, för att i Jisreel låta hela sig från de sår som han hade fått vid Rama, i striden mot Hasael, konungen i Aram.
Och Asarja, Jorams son, Juda konung, for ned för att besöka Joram, Ahabs son, i Jisreel, eftersom denne låg sjuk.
Men till Ahasjas fördärv var det av Gud bestämt att han skulle komma till Joram.
Ty när han hade kommit dit, for han med Joram för att möta Jehu, Nimsis son, som HERREN hade smort till att utrota Ahabs hus.
Så hände sig att Jehu, när han utförde straffdomen över Ahabs hus, träffade på de Juda furstar och de brorsöner till Ahasja, som voro i Ahasjas tjänst, och dräpte dem.
Sedan sökte han efter Ahasja; och man grep denne, där han höll sig gömd i Samaria, och förde honom till Jehu och dödade honom.
Men därefter begrovo de honom, ty de sade: »Han var dock son till Josafat, som sökte HERREN av allt sitt hjärta.»
Och av Ahasjas hus fanns sedan ingen dom förmådde övertaga konungadömet.
När nu Atalja, Ahasjas moder, förnam att hennes son var död, stod hon upp och förgjorde hela konungasläkten i Juda hus.
Men just när konungabarnen skulle dödas, tog konungadottern Josabeat Joas, Ahasjas son, och skaffade honom hemligen undan, i det att han förde honom jämte hans amma in i sovkammaren; där höll Josabeat, konung Jorams dotter, prästen Jojadas hustru -- som ju ock var Ahasjas syster -- honom dold för Atalja, så att denna icke fick döda honom.
Sedan var han hos dem i Guds hus, där han förblev gömd i sex år, medan Atalja regerade i landet.
Men i det sjunde året tog Jojada mod till sig och förband sig med underhövitsmännen Asarja, Jerohams son, Ismael, Johanans son, Asarja, Obeds son, Maaseja, Adajas son, och Elisafat, Sikris son.
Dessa foro därefter omkring i Juda och församlade leviterna ur alla Juda städer, så ock huvudmännen för Israels familjer.
Och när de kommo till Jerusalem,
Slöt hela församlingen i Guds hus ett förbund med konungen.
Och Jojada sade till dem: »Konungens son skall nu vara konung, såsom HERREN har talat angående Davids söner.
Detta är alltså vad I skolen göra: en tredjedel av eder, nämligen de präster och leviter som hava att inträda i vakthållningen på sabbaten, skall stå på vakt vid trösklarna
och en tredjedel vid konungshuset och en tredjedel vid Jesodporten; och allt folket skall vara på förgårdarna till HERRENS hus.
Dock må ingen annan än prästerna och de tjänstgörande leviterna gå in i HERRENS hus; dessa må gå in, ty de äro heliga.
Men allt det övriga folket skall iakttaga vad HERREN har bjudit dem iakttaga.
Och leviterna skola ställa sig runt omkring konungen, var och en med sina vapen i handen; och om någon vill tränga sig in i huset, skall han dödas.
Och I skolen följa konungen, vare sig han går in eller ut.»
Leviterna och hela Juda gjorde allt vad prästen Jojada hade bjudit dem, var och en av dem tog sina män, både de som skulle inträda i vakthållningen på sabbaten och de som skulle avgå därifrån på sabbaten, ty prästen Jojada lät ingen avdelning vara fri ifrån tjänstgöring.
Och prästen Jojada gav åt underhövitsmännen de spjut och de sköldar av olika slag, som hade tillhört konung David, och som funnos i Guds hus.
Och han ställde upp allt folket, var och en med sitt vapen i handen, från husets södra sida till husets norra sida, mot altaret och mot huset, runt omkring konungen.
Därefter förde de ut konungasonen och satte på honom kronan och gåvo honom vittnesbördet och gjorde honom till konung; och Jojada och hans söner smorde honom och ropade: »Leve konungen!»
När Atalja nu hörde folkets rop, då de skyndade fram och hyllade konungen, gick hon in i HERRENS hus till folket.
Där fick hon då se konungen stå vid sin pelare, nära ingången, och hövitsmännen och trumpetblåsarna bredvid konungen, och fick höra huru hela folkmängden jublade och stötte i trumpeterna, och huru sångarna med sina instrumenter ledde hyllningssången.
Då rev Atalja sönder sina kläder och ropade: »Sammansvärjning!
Sammansvärjning!»
Men prästen Jojada lät underhövitsmännen som anförde skaran träda fram, och han sade till dem: »Fören henne ut mellan leden, och om någon följer henne, så må han dödas med svärd.»
Prästen förbjöd dem nämligen att döda henne i HERRENS hus.
Alltså grepo de henne, och när hon hade kommit fram dit där Hästporten för in i konungshuset, dödade de henne där.
Och Jojada slöt ett förbund mellan sig och allt folket och konungen, att de skulle vara ett HERRENS folk.
Och allt folket begav sig till Baals tempel och rev ned det och slog sönder dess altaren och bilder; och Mattan, Baals präst, dräpte de framför altarna.
Därefter ställde Jojada ut vakter vid HERRENS hus och betrodde detta värv åt de levitiska prästerna, dem som David hade indelat i klasser för tjänstgöringen i HERRENS hus, till att offra brännoffer åt HERREN, såsom det var föreskrivet i Moses lag, med jubel och sång, efter Davids anordning.
Och han ställde dörrvaktarna vid portarna till HERRENS hus, för att ingen skulle komma in, som på något sätt var oren.
Och han tog med sig underhövitsmännen och de förnämsta och mäktigaste bland folket och hela folkmängden och förde konungen ned från HERRENS hus, och de gingo in i konungshuset genom Övre porten; och de satte konungen på konungatronen.
Och hela folkmängden gladde sig, och staden förblev lugn.
Men Atalja hade de dödat med svärd.
Joas var sju år gammal, när han blev konung, och han regerade fyrtio år i Jerusalem.
Hans moder hette Sibja, från Beer-Seba.
Och Joas gjorde vad rätt var i HERRENS ögon, så länge prästen Jojada levde.
Och Jojada tog åt honom två hustrur, och han födde söner och döttrar.
Därefter blev Joas betänkt på att upphjälpa HERRENS hus.
Och han församlade prästerna och leviterna och sade till dem: »Faren vart år ut till Juda städer, och samlen från hela Israel in penningar till att sätta eder Guds hus i stånd; och I skolen bedriva denna sak med skyndsamhet.»
Men leviterna skyndade sig icke.
Då kallade konungen till sig översteprästen Jojada och sade till honom: »Varför har du icke tillhållit leviterna att från Juda och Jerusalem indriva den skatt som HERRENS tjänare Mose pålade, och som Israels församling skulle erlägga till vittnesbördets tabernakel?
Ty Ataljas, den ogudaktiga kvinnans, söner hava fördärvat Gud hus; ja, allt som var helgat till HERRENS hus hava de använt till Baalerna.»
På konungens befallning gjorde man därefter en kista och ställde den utanför porten till HERREN hus.
Och man lät utropa i Juda och Jerusalem att den skatt som Guds tjänare Mose hade pålagt Israel i öknen skulle erläggas åt HERREN.
Och alla furstarna och allt folket buro fram penningar med glädje och kastade dem i kistan, till dess att allt var insamlat.
Och när tid blev att genom leviternas försorg föra kistan till de granskningsmän som konungen hade förordnat, och dessa då märkte att mycket penningar fanns i den, då kommo konungens sekreterare och översteprästens tillsyningsman och tömde kistan och buro den sedan tillbaka till dess plats.
Så gjorde de gång efter annan och samlade in penningar i myckenhet.
Därefter lämnade konungen och Jojada dessa åt den som skulle utföra arbetet på HERRENS hus, och lejde stenhuggare och timmermän till att upphjälpa HERRENS hus, så ock järn- och kopparsmeder till att sätta HERRENS hus i stånd.
Och de som utförde arbetet bedrevo det så, att arbetet gick framåt under deras händer, Och de återställde Guds hus i dess förra skick och satte det i gott stånd.
Och när de hade slutat, buro de återstoden av penningarna till konungen och Jojada; och man gjorde därav kärl till HERRENS hus, kärl till gudstjänsten och offren, skålar och andra kärl av guld och silver Och man offrade brännoffer i HERRENS hus beständigt, så länge Jojada levde.
Men Jojada blev gammal och mätt på att leva och dog så; ett hundra trettio år gammal var han vid sin död.
Och man begrov honom i Davids stad bland konungarna, därför att han hade gjort vad gott var mot Israel och mot Gud och hans hus.
Men efter Jojadas död kommo Juda furstar och föllo ned för konungen; då lyssnade konungen till dem.
Och de övergåvo HERRENS, sina fäders Guds, hus och tjänade Aserorna och avgudarna.
Då kom förtörnelse över Juda och Jerusalem genom den skuld de så ådrogo sig.
Och profeter sändes ibland dem för att omvända dem till HERREN; och dessa varnade dem, men de lyssnade icke därtill.
Men Sakarja, prästen Jojadas son, hade blivit beklädd med Guds Andes kraft, och han trädde fram inför folket och sade till dem: »Så säger Gud: Varför överträden I HERRENS bud, eder själva till ingen fromma?
Eftersom I haven övergivit HERREN, har han ock övergivit eder.»
Då sammansvuro de sig mot honom och stenade honom, enligt konungens befallning, på förgården till HERRENS hus.
Ty konung Joas tänkte icke på den kärlek som Jojada, dennes fader, hade bevisat honom, utan dräpte hans son.
Men denne sade i sin dödsstund: »Må HERREN se detta och utkräva det.»
Och när året hade gått till ända, drog araméernas här upp mot honom, och de kommo till Juda och Jerusalem och utrotade ur folket alla folkets furstar.
Och allt byte som de togo sände de till konungen i Damaskus.
Ty fastän araméernas här som då ryckte an utgjorde allenast en ringa skara, gav HERREN likväl i deras hand en mycket talrik här, därför att folket hade övergivit HERREN, sina fäders Gud.
Så fingo de utföra straffdomen över Joas.
Och när dessa drogo bort ifrån honom -- ty de lämnade honom kvar illa sjuk -- sammansvuro sig hans tjänare mot honom, därför att han hade utgjutit prästen Jojadas söners blod, och dräpte honom på hans säng; detta blev hans död.
Och man begrov honom i Davids stad; dock begrov man honom icke i konungagravarna.
Och de som sammansvuro sig mot honom voro Sabad, son till ammonitiskan Simeat, och Josabad, son till moabitiskan Simrit.
Men om hans söner, och om de många profetior som förkunnades mot honom, och om huru Guds hus åter upprättades, härom är skrivet i »Utläggning av Konungaboken».
Och hans son Amasja blev konung efter honom.
Amasja var tjugufem år gammal, när han blev konung, och han regerade tjugunio år i Jerusalem.
Hans moder hette Joaddan, från Jerusalem.