Han gjorde vad rätt var i HERRENS ögon, dock icke av fullt hängivet hjärta.
Och sedan hans konungadöme hade blivit befäst, lät han dräpa dem av sina tjänare, som hade dödat hans fader, konungen.
Men deras barn dödade han icke, utan handlade i enlighet med vad föreskrivet var i Moses lagbok, där HERREN hade bjudit och sagt: »Föräldrarna skola icke dö för sina barns skull, och barnen skola icke dö för sina föräldrars skull, utan var och en skall dö genom sin egen synd.»
Och Amasja församlade Juda barn och lät dem ställa upp sig efter sina familjer, efter sina över- och under- hövitsmän, hela Juda och Benjamin.
Därefter inmönstrade han dem som voro tjugu år gamla eller därutöver, och fann dem utgöra tre hundra tusen utvalda stridbara män, som kunde föra spjut och sköld.
Därtill lejde han för hundra talenter silver ett hundra tusen tappra stridsmän ur Israel.
Men en gudsman kom till honom och sade: »O konung, låt icke Israels här draga åstad med dig, ty HERREN är icke med Israel, icke med hela hopen av Efraims barn;
utan du själv må allena draga åstad.
Grip verket an, gå frimodigt ut i striden.
Gud skall eljest låta dig komma på fall genom fienden; ty Gud förmår både att hjälpa och att stjälpa.»
Amasja sade till gudsmannen: »Men huru skall det då gå med de hundra talenterna som jag har givit åt skaran från Israel?»
Gudsmannen svarade: »HERREN kan väl giva dig mer än det.»
Då avskilde Amasja den skara som hade kommit till honom från Efraim och lät dem gå hem igen.
Häröver blevo dessa högeligen förgrymmade på Juda och vände tillbaka hem i vredesmod.
Men Amasja tog mod till sig och tågade ut med sitt folk och drog till Saltdalen och nedgjorde där av Seirs barn tio tusen.
Och Juda barn togo andra tio tusen till fånga levande; dem förde de upp på spetsen av en klippa och störtade dem ned från klippspetsen, så att de alla krossades.
Men de som tillhörde den skara som Amasja hade sänt tillbaka, och som icke hade fått gå med honom ut i striden, företogo plundringståg i Juda städer, från Samaria ända till Bet-Horon; och de nedgjorde tre tusen av invånarna och togo stort byte.
När sedan Amasja kom tillbaka från sin seger över edoméerna, förde han med sig Seirs barns gudar och ställde upp dem till gudar åt sig; och han tillbad inför dem och tände offereld åt dem.
Då upptändes HERRENS vrede mot Amasja, och han sände till honom en profet; denne sade till honom: »Varför söker du detta folks gudar, som ju icke hava kunnat rädda sitt eget folk ur din hand?»
När denne så talade till honom, svarade han honom: »Hava vi satt dig till konungens rådgivare?
Håll upp, om du icke vill att man skall dräpa dig.»
Då höll profeten upp och sade: »Jag förstår nu att Gud har beslutit att fördärva dig, eftersom du gör på detta sätt och icke vill höra på mitt råd.»
Och sedan Amasja, Juda konung, hade hållit rådplägning, sände han till Joas, son till Joahas, son till Jehu, Israels konung, och lät säga: »Kom, låt oss drabba samman med varandra.»
Men Joas, Israels konung, sände då till Amasja, Juda konung, och lät svara: »Törnbusken på Libanon sände en gång bud till cedern på Libanon och lät säga: 'Giv din dotter åt min son till hustru.'
Men sedan gingo markens djur på Libanon fram över törnbusken och trampade ned den.
Du tänker på huru du har slagit Edom, och däröver förhäver du dig ditt hjärta och vill vinna ännu mer ära.
Men stanna nu hemma.
Varför utmanar du olyckan, dig själv och Juda med dig till fall?»
Men Amasja ville icke höra härpå, ty Gud skickade det så, för att de skulle bliva givna i fiendehand, eftersom de hade sökt Edoms gudar.
Så drog då Joas, Israels konung, upp, och de drabbade samman med varandra, han och Amasja, Juda konung, vid det Bet-Semes som hör till Juda.
Och Juda män blevo slagna av Israels män och flydde, var och en till sin hydda.
Och Amasja, Juda konung, son till Joas, son till Joahas, blev tagen till fånga i Bet-Semes av Joas, Israels konung.
Och när denne hade fört honom till Jerusalem, bröt han ned ett stycke av Jerusalems mur, från Efraimsporten ända till Poneporten, fyra hundra alnar.
Och han tog allt guld och silver och alla kärl som funnos i Guds hus, hos Obed-Edom, och konungshusets skatter, därtill ock gisslan, och vände så tillbaka till Samaria.
Men Amasja, Joas' son, Juda konung, levde i femton år efter Joas', Joahas' sons, Israels konungs, död.
Vad nu mer är att säga om Amasja, om hans första tid såväl som om hans sista, det finnes upptecknat i boken om Judas och Israels konungar.
Och från den tid då Amasja vek av ifrån HERREN begynte man anstifta en sammansvärjning mot honom i Jerusalem, så att han måste fly till Lakis.
Då sändes män efter honom till Lakis, och dessa dödade honom där.
Sedan förde man honom därifrån på hästar och begrov honom hos hans fäder i Juda huvudstad.
Och allt folket i Juda tog Ussia, som då var sexton år gammal, och gjorde honom till konung i hans fader Amasjas ställe.
Det var han som befäste Elot, och han lade det åter under Juda, sedan konungen hade gått till vila hos sina fäder.
Ussia var sexton år gammal, när han blev konung, och han regerade femtiotvå år i Jerusalem.
Hans moder hette Jekilja, från Jerusalem.
Han gjorde vad rätt var i HERRENS ögon, alldeles såsom hans fader Amasja hade gjort.
Och han sökte Gud, så länge Sakarja levde, han som aktade på Guds syner.
Och så länge han sökte HERREN, lät Gud det gå honom väl.
Han drog ut och stridde mot filistéerna och bröt ned Gats, Jabnes och Asdods murar; och han byggde städer på Asdods område och annorstädes i filistéernas land.
Och Gud hjälpte honom mot filistéerna och mot de araber som bodde i Gur-Baal och mot maoniterna.
Och ammoniterna måste giva skänker åt Ussia, och ryktet om honom sträckte sig ända till Egypten, ty han blev övermåttan mäktig.
Och Ussia byggde torn i Jerusalem över Hörnporten och över Dalporten och över Vinkeln och befäste dem.
Han byggde ock torn i öknen och högg ut många brunnar, ty han hade mycken boskap, både i låglandet och på slätten.
Jordbruks- och vingårdsarbetare hade han i bergsbygden och på de bördiga fälten, ty han var en vän av åkerbruk.
Och Ussia hade en krigshär som drog ut till strid i avdelade skaror, med en mansstyrka som hade blivit fastställd vid mönstring genom sekreteraren Jeguel och tillsyningsmannen Maaseja, under överinseende av Hananja, en av konungens hövitsmän.
Hela antalet av de tappra stridsmän som voro huvudmän för familjerna var två tusen sex hundra.
Under deras befäl stod en krigshär av tre hundra sju tusen fem hundra män, som stridde med kraft och mod och voro konungens hjälp mot fienden.
Och Ussia försåg hela denna här med sköldar, spjut, hjälmar, pansar och bågar, så ock med slungstenar.
Och han lät i Jerusalem göra krigsredskap, konstmässigt uttänkta, till att sätta upp på tornen och på murarnas hörn, för att med dem avskjuta pilar och stora stenar.
Och ryktet om honom gick ut vida omkring, ty underbart hjälptes han fram till makt.
Men när han nu var så mäktig, blev hans hjärta högmodigt, så att han gjorde vad fördärvligt var; han förbröt sig trolöst mot HERREN, sin Gud, i det att han gick in i HERRENS tempel för att antända rökelse på rökelsealtaret.
Då gick prästen Asarja ditin efter honom, åtföljd av åttio HERRENS präster, oförskräckta män.
Dessa trädde fram mot konung Ussia och sade till honom: »Det hör icke dig till, Ussia, att antända rökelse åt HERREN, utan det tillhör prästerna, Arons söner, som är helgade till att antända rökelse.
Gå ut ur helgedomen, ty du har begått en förbrytelse, och HERREN Gud skall icke låta detta lända dig till ära.»
Då for Ussia ut i vrede, där han stod med ett rökelsekar i sin hand för att antända rökelse.
Men just som han for ut mot prästerna, slog spetälska ut på hans panna, i prästernas närvaro, inne i HERRENS hus, bredvid rökelsealtaret.
Och när översteprästen Asarja och alla prästerna vände sig till honom och fingo se att han var spetälsk i pannan, drevo de honom strax ut därifrån.
Själv skyndade han också ut, eftersom HERREN så hemsökte honom.
Sedan var konung Ussia spetälsk för hela sitt liv och bodde i ett särskilt hus såsom spetälsk, ty han var utesluten från HERRENS hus.
Hans son Jotam förestod då konungens hus och dömde folket i landet.
Vad nu mer är att säga om Ussia, om hans första tid såväl som om hans sista, det har profeten Jesaja, Amos' son, tecknat upp.
Och Ussia gick till vila hos sina fäder, och man begrov honom hos hans fäder, ute på konungagravens mark, detta med tanke därpå att han hade varit spetälsk.
Och hans son Jotam blev konung efter honom.
Jotam var tjugufem år gammal när han blev konung, och han regerade sexton år i Jerusalem.
Hans moder hette Jerusa, Sadoks dotter.
Han gjorde vad rätt var i HERRENS ögon, alldeles såsom hans fader Ussia hade gjort, vartill kom att han icke trängde in i HERRENS tempel; men folket gjorde ännu vad fördärvligt var.
Han byggde Övre porten till HERRENS hus, och på Ofelmuren utförde han stora byggnadsarbeten.
Därtill byggde han städer i Juda bergsbygd, och i skogarna byggde han borgar och torn.
Och när han så kom i strid med Ammons barns konung, blev han dem övermäktig, så att Ammons barn det året måste giva honom ett hundra talenter silver, tio tusen korer vete och tio tusen korer korn.
Lika mycket måste Ammons barn erlägga åt honom också nästa år och året därpå.
Så mäktig blev Jotam, därför att han vandrade ståndaktigt inför HERREN, sin Gud.
Vad nu mer är att säga om Jotam och om alla hans krig och andra företag, det finnes upptecknat i boken om Israels och Juda konungar.
Han var tjugufem år gammal, när han blev konung, och han regerade sexton år i Jerusalem.
Och Jotam gick till vila hos sina fäder, och man begrov honom i Davids stad.
Och hans son Ahas blev konung efter honom.
Ahas var tjugu år gammal när han blev konung, och han regerade sexton år i Jerusalem.
Han gjorde icke vad rätt var i HERRENS ögon, såsom hans fader David,
utan vandrade på Israels konungars väg; ja, han lät ock göra gjutna beläten åt Baalerna.
Och själv tände han offereld i Hinnoms sons dal och brände upp sina barn i eld, efter den styggeliga seden hos de folk som HERREN hade fördrivit för Israels barn.
Och han frambar offer och tände offereld på höjderna och kullarna och under alla gröna träd.
Därför gav HERREN, hans Gud, honom i den arameiske konungens hand; de slogo honom och togo av hans folk en stor hop fångar och förde dem till Damaskus.
Han blev ock given i Israels konungs hand, så att denne tillfogade honom ett stort nederlag.
Ty Peka, Remaljas son, dräpte av Juda ett hundra tjugu tusen man på en enda dag, allasammans stridbara män.
Detta skedde därför att de hade övergivit HERREN, sina fäders Gud.
Och Sikri, en tapper man från Efraim, dräpte Maaseja, konungasonen, och Asrikam, slottshövdingen, och Elkana, konungens närmaste man.
Och Israels barn bortförde från sina bröder två hundra tusen fångar, nämligen deras hustrur, söner och döttrar, och togo därjämte mycket byte från dem och förde bytet till Samaria.
Men där var en HERRENS profet som hette Oded; denne gick ut mot hären, när den kom till Samaria, och sade till dem: »Se, i sin vrede över Juda har HERREN, edra fäders Gud, givit dem i eder hand, men I haven dräpt dem med en hätskhet som har nått upp till himmelen.
Och nu tänken I göra Judas och Jerusalems barn till trälar och trälinnor åt eder.
Därmed dragen I ju allenast skuld över eder själva inför HERREN, eder Gud.
Så hören mig nu: Sänden tillbaka fångarna som I haven tagit från edra bröder; ty HERRENS vrede är upptänd mot eder.»
Några av huvudmännen bland Efraims barn, nämligen Asarja, Johanans son, Berekja, Mesillemots son, Hiskia, Sallums son, och Amasa, Hadlais son, stodo då upp och gingo emot dem som kommo från kriget
och sade till dem: »I skolen icke föra dessa fångar hitin; ty I förehaven något som drager skuld över oss inför HERREN, och varigenom I ytterligare föröken våra synder och vår skuld.
Vår skuld är ju redan stor nog, och vrede är upptänd mot Israel.»
Då lämnade krigsfolket ifrån sig fångarna och bytet inför de överste och hela församlingen.
Och de nämnda männen stodo upp och togo sig an fångarna.
Alla som voro nakna bland dem klädde de upp med vad de hade tagit såsom byte; de gåvo dem kläder och skor, mat och dryck, och smorde dem med olja, och alla som icke orkade gå läto de sätta sig upp på åsnor, och förde dem så till Jeriko, Palmstaden, till deras bröder där.
Sedan vände de tillbaka till Samaria.
Vid samma tid sände konung Ahas bud till konungarna i Assyrien, med begäran att de skulle hjälpa honom.
Ty förutom allt annat hade edoméerna kommit och slagit Juda och tagit fångar.
Och filistéerna hade fallit in i städerna i Juda lågland och sydland och hade intagit Bet-Semes, Ajalon och Gederot, så ock Soko med underlydande orter, Timna med underlydande orter och Gimso med underlydande orter, och hade bosatt sig i dem.
Ty HERREN ville förödmjuka Juda, för Ahas', den israelitiske konungens, skull, därför att denne hade vållat oordning i Juda och varit otrogen mot HERREN.
Men Tillegat-Pilneeser, konungen i Assyrien, drog emot honom och angrep honom, i stället för att understödja honom.
Ty fastän Ahas plundrade HERRENS hus och konungshuset och de överstes hus och gav allt åt konungen i Assyrien, så hjälpte det honom dock icke.
Och i sin nöd försyndade sig samme konung Ahas ännu mer genom otrohet mot HERREN.
Han offrade nämligen åt gudarna i Damaskus, som hade slagit honom; ty han tänkte: »Eftersom de arameiska konungarnas gudar hava förmått hjälpa dem, vill jag offra åt dessa gudar, för att de ock må hjälpa mig.»
Men i stället var det dessa som kommo honom och hela Israel på fall.
Ahas samlade ihop de kärl som funnos i Guds hus och bröt sönder kärlen i Guds hus och stängde igen dörrarna till HERRENS hus, och gjorde sig altaren i vart hörn i Jerusalem.
Och i var och en av Juda städer uppförde han offerhöjder för att där tända offereld åt andra gudar, och han förtörnade så HERREN, sina fäders Gud.
Vad nu mer är att säga om honom och om alla hans företag, under hans första tid såväl som under hans sista, det finnes upptecknat i boken om Judas och Israels konungar.
Och Ahas gick till vila hos sina fäder, och man begrov honom i Jerusalem, inne i själva staden; de lade honom nämligen icke i Israels konungars gravar.
Och hans son Hiskia blev konung efter honom.
Hiskia var tjugufem år gammal, när han blev konung, och han regerade tjugunio år i Jerusalem.
Hans moder hette Abia, Sakarjas dotter.
Han gjorde vad rätt var i HERRENS ögon, alldeles såsom hans fader David hade gjort.
I sitt första regeringsår, i första månaden, öppnade han dörrarna till HERRENS hus och satte dem i stånd
Och han lät hämta prästerna och leviterna och församlade dem på den öppna platsen mot öster.
Och han sade till dem: »Hören mig, I leviter.
Helgen nu eder själva, och helgen HERRENS, edra fäders Guds, hus, och skaffen orenheten ut ur helgedomen.
Ty våra fäder voro otrogna och gjorde vad ont var i HERRENS, vår Guds, ögon och övergåvo honom; de vände sitt ansikte bort ifrån HERRENS boning och vände honom ryggen.
De stängde ock igen dörrarna till förhuset, släckte ut lamporna, tände ingen rökelse och offrade inga brännoffer i helgedomen åt Israels Gud.
Därför har HERRENS förtörnelse kommit över Juda och Jerusalem, och han har gjort dem till en varnagel, till ett föremål för häpnad och begabberi, såsom I sen med egna ögon.
Ja, därför hava ock våra fäder fallit för svärd, och våra söner och döttrar och hustrur hava fördenskull kommit i fångenskap.
Men nu har jag i sinnet att sluta ett förbund med HERREN, Israels Gud, för att hans vredes glöd må vända sig ifrån oss.
Så varen nu icke försumliga, mina barn, ty eder har HERREN utvalt till att stå inför hans ansikte och göra tjänst inför honom, till att vara hans tjänare och antända rökelse åt honom.»
Då stodo leviterna upp: Mahat, Amasais son, och Joel, Asarjas son, av kehatiternas barn; av Meraris barn Kis, Abdis son, och Asarja, Jehallelels son; av gersoniterna Joa, Simmas son, och Eden, Joas son;
av Elisafans barn Simri och Jeguel; av Asafs barn Sakarja och Mattanja;
av Hemans barn Jehuel och Simei; av Jedutuns barn Semaja och Ussiel.
Dessa församlade nu sina bröder och helgade sig och gingo, såsom konungen hade bjudit i kraft av HERRENS ord, sedan in för att rena HERRENS hus.
Men prästerna gingo in i det inre av HERRENS hus för att rena det, och all orenhet som de funno i HERRENS tempel buro de ut på förgården till HERRENS hus; där togo leviterna emot den och buro ut den i Kidrons dal.
De begynte att helga templet på första dagen i första månaden, och på åttonde dagen i månaden hade de hunnit till HERRENS förhus och helgade sedan HERRENS hus under åtta dagar; och på sextonde dagen i första månaden hade de fullgjort sitt arbete.
Då gingo de in till konung Hiskia och sade: »Vi hava renat hela HERRENS hus och brännoffersaltaret med alla dess tillbehör och skådebrödsbordet med alla dess tillbehör.
Och alla de kärl som konung Ahas under sin regering i sin otrohet förkastade, dem hava vi återställt och helgat, och de stå nu framför HERRENS altare.»
Då lät konung Hiskia bittida om morgonen församla de överste i staden och gick upp i HERRENS hus.
Och man förde fram sju tjurar, sju vädurar och sju lamm, så ock sju bockar till syndoffer för riket och för helgedomen och för Juda; och han befallde Arons söner, prästerna, att offra detta på HERRENS altare.
Då slaktade de fäkreaturen, och prästerna togo upp blodet och stänkte det på altaret; därefter slaktade de vädurarna och stänkte blodet på altaret; sedan slaktade de lammen och stänkte blodet på altaret.
Därefter förde de syndoffersbockarna fram inför konungen och församlingen, och de lade sina händer på dem.
Och prästerna slaktade dem och läto deras blod såsom syndoffer komma på altaret, till försoning för hela Israel; ty konungen hade befallt att offra dessa brännoffer och syndoffer för hela Israel.
Och han lät leviterna ställa upp sig till tjänstgöring i HERRENS hus med cymbaler, psaltare och harpor, såsom David och Gad, konungens siare, och profeten Natan hade bjudit; ty budet härom var givet av HERREN genom hans profeter.
Och leviterna ställde upp sig med Davids instrumenter, och prästerna med trumpeterna.
Och Hiskia befallde att man skulle offra brännoffret på altaret; och på samma gång som offret begynte, begynte ock HERRENS sång ljuda jämte trumpeterna, och detta under ledning av Davids, Israels konungs, instrumenter.
Och hela församlingen föll ned, under det att sången sjöngs och trumpeterna skallade -- allt detta ända till dess brännoffret var fullbordat.
Och när de hade offrat brännoffret, knäböjde konungen och alla som voro där tillstädes med honom, och tillbådo.
Och konung Hiskia och de överste befallde leviterna att lova HERREN med Davids och siaren Asafs ord; och de sjöngo hans lov med glädje och böjde sig ned och tillbådo.
Och Hiskia tog till orda och sade: »I haven nu tagit handfyllning till HERRENS tjänst.
Så träden nu hit och fören fram slaktoffer och lovoffer till HERRENS hus.»
Då förde församlingen fram slaktoffer och lovoffer, och var och en som av sitt hjärta manades därtill offrade brännoffer.
Antalet av de brännoffersdjur som församlingen förde fram var sjuttio tjurar, ett hundra vädurar och två hundra lamm, alla dessa till brännoffer åt HERREN.
Och tackoffren utgjordes av sex hundra tjurar och tre tusen djur av småboskapen.
Men prästerna voro för få, så att de icke kunde draga av huden på alla brännoffersdjuren; därför understöddes de av sina bröder leviterna, till dess detta göromål var fullgjort, och till dess prästerna hade helgat sig.
Ty i fråga om att helga sig hade leviterna visat sig mer rättsinniga än prästerna.
Också var antalet stort av brännoffer, vartill kommo fettstyckena från tackoffren, så ock de drickoffer som hörde till brännoffren.
Så blev det ordnat med tjänstgöringen i HERRENS hus.
Och Hiskia och allt folket gladde sig över vad Gud hade berett åt folket; ty helt oväntat hade detta kommit till stånd.
Därefter sände Hiskia ut bud till hela Israel och Juda och skrev också brev till Efraim och Manasse, att de skulle komma till HERRENS hus i Jerusalem för att hålla HERRENS, Israels Guds, påskhögtid.
Och konungen och hans förnämsta män och hela församlingen i Jerusalem enade sig om att hålla påskhögtiden i andra månaden;
ty de kunde icke hålla den nu genast, eftersom prästerna ännu icke hade helgat sig i tillräckligt antal och folket icke hade hunnit församla sig till Jerusalem.
Därför syntes det konungen och hela församlingen rätt att göra så.
Och de beslöto att låta utropa i hela Israel, från Beer-Seba ända till Dan, att man skulle komma och hålla HERRENS, Israels Guds, påskhögtid i Jerusalem; ty man hade icke eljest hållit den samfällt, såsom föreskrivet var.
Så begåvo sig då ilbuden åstad med breven från konungen och hans förnämsta män och drogo genom hela Israel och Juda, enligt konungens befallning, och sade: »I Israels barn, vänden om till HERREN, Abrahams, Isaks och Israels Gud, på det att han må vända om till den kvarleva av eder, som har räddats undan de assyriska konungarnas hand.
Och varen icke såsom edra fäder och bröder, som voro otrogna mot HERREN, sina fäders Gud, så att han prisgav dem åt förödelse, såsom I själva haven sett.
Varen alltså nu icke hårdnackade såsom edra fäder, utan underkasten eder HERREN och kommen till hans helgedom, den som han har helgat för evig tid, och tjänen HERREN, eder Gud, på det att hans vredes glöd må vända sig ifrån eder.
Ty om I vänden om till HERREN, skola edra bröder och edra barn finna barmhärtighet inför dem som hålla dem fångna, så att de få vända tillbaka till detta land; ty HERREN, eder Gud, är nådig och barmhärtig, och han skall icke vända sitt ansikte ifrån eder, om I vänden om till honom.»
Och ilbuden foro ifrån stad till stad i Efraims och Manasse land och ända till Sebulon; men man gjorde spe av dem och bespottade dem.
Dock funnos några i Aser, Manasse och Sebulon, som ödmjukade sig och kommo till Jerusalem.
Också i Juda verkade Guds hand, så att han gav dem ett endräktigt hjärta till att göra efter vad konungen och de överste hade bjudit i kraft av HERRENS ord.
Och mycket folk kom tillhopa i Jerusalem för att hålla det osyrade brödets högtid i andra månaden, en mycket stor församling.
Och de stodo upp och skaffade bort de altaren som funnos i Jerusalem; också alla offereldsaltarna skaffade de bort och kastade dem i Kidrons dal.
Och de slaktade påskalammet på fjortonde dagen i andra månaden; prästerna och leviterna, som nu kände blygsel och därför hade helgat sig, förde därvid fram brännoffer till HERRENS hus.
Och de inställde sig till tjänstgöring på sina platser, såsom det var föreskrivet för dem, efter gudsmannen Moses lag; och prästerna stänkte med blodet, sedan de hade tagit emot det av leviterna.
Ty många funnos i församlingen, som icke hade helgat sig; därför måste leviterna slakta påskalammen för alla som icke voro rena, och så helga dem åt HERREN.
Det var nämligen en myckenhet av folket, många från Efraim och Manasse, Isaskar och Sebulon, som icke hade renat sig, utan åto påskalammet på annat sätt än föreskrivet var.
Men Hiskia hade bett för dem och sagt: »HERREN, den gode, förlåte var och en
som har vänt sitt hjärta till att söka Gud, HERREN, sina fäders Gud, om han än icke är ren efter helgedomens ordning.»
Och HERREN hörde Hiskia och skonade folket.
Så höllo Israels barn, de som då voro tillstädes i Jerusalem, det osyrade brödets högtid i sju dagar med stor glädje; och leviterna och prästerna lovade HERREN var dag med kraftiga instrumenter, HERREN till ära.
Och Hiskia talade vänligt till alla de leviter som voro väl förfarna i HERRENS tjänst.
Och de åto av högtidsoffren under de sju dagarna, i det att de offrade tackoffer och prisade HERREN, sina faders Gud.
Och hela församlingen enade sig om att hålla högtid under ännu sju dagar; och så höll man högtid med glädje också under de sju dagarna.
Ty Hiskia, Juda konung, hade såsom offergärd givit åt församlingen ett tusen tjurar och av småboskapen sju tusen djur, och de överste hade såsom offergärd givit åt församlingen ett tusen tjurar och av småboskapen tio tusen djur.
Och ett stort antal präster helgade sig.
Och hela Juda församling gladde sig med prästerna och leviterna, så ock hela församlingen av dem som hade kommit från Israel, ävensom de främlingar som hade kommit från Israels land, eller som bodde i Juda.
Och i Jerusalem var stor glädje; ty alltsedan Salomos, Davids sons, Israels konungs, tid hade icke något sådant som detta skett i Jerusalem.
Och de levitiska prästerna stodo upp och välsignade folket, och deras röst blev hörd, och deras bön kom till himmelen, hans heliga boning.
När nu allt detta var till ända, drogo alla israeliter som hade varit där tillstädes ut till Juda städer och slogo sönder stoderna, höggo ned Aserorna och bröto ned offerhöjderna och altarna i hela Juda och Benjamin och i Efraim och Manasse, till dess att de hade gjort ände på dem; sedan vände alla Israels barn tillbaka till sina städer, var och en till sin egendom.
Och Hiskia förordnade om prästernas och leviternas avdelningar, alltefter som de tillhörde den ena eller den andra avdelningen, så att var och en av såväl prästerna som leviterna fick sitt bestämda göromål, när brännoffer och tackoffer skulle offras, till att därvid göra tjänst och tacka och lovsjunga i portarna till HERRENS läger.
Och konungen anslog en del av sin egendom till brännoffren, nämligen till att offra brännoffer morgon och afton, och till att offra brännoffer på sabbaterna, vid nymånaderna och vid högtiderna, såsom det var föreskrivet i HERRENS lag.
Och han befallde folket som bodde i Jerusalem att giva prästerna och leviterna deras del, för att de skulle kunna hålla fast vid HERRENS lag.
Och när denna befallning blev känd, gåvo Israels barn rikligen en förstling av säd, vin, olja och honung och av all markens avkastning; och tionde av allt förde de fram i myckenhet.
Och de av Israels och Juda barn, som bodde i Juda städer, förde ock fram tionde av fäkreatur och små boskap, så ock tionde av de heliga gåvor som helgades åt HERRENS, deras Gud, och lade upp dem i särskilda högar.
I tredje månaden begynte de att lägga upp högarna, och i sjunde månaden hade de slutat därmed.
När då Hiskia och de överste kommo och sågo högarna, prisade de HERREN och hans folk Israel.
Och Hiskia frågade prästerna och leviterna om högarna.
Då svarade honom översteprästen Asarja, av Sadoks hus, och sade; »Alltsedan man begynte föra fram offergärden till HERRENS hus, hava vi ätit och blivit mätta och dock fått mycket kvar; ty HERREN har välsignat sitt folk, och vad som är kvar är denna stora rikedom.»
Och Hiskia befallde att man skulle inreda förrådskamrar i HERRENS hus, och man inredde sådana.
Och i dem förde man in offergärden och tionden och de heliga gåvorna, allt på heder och tro.
Och överuppsyningsman däröver var leviten Konanja, och hans närmaste man var hans broder Simei.
Men Jehiel, Asasja, Nahat, Asael, Jerimot, Josabad, Eliel, Jismakja, Mahat och Benaja voro tillsyningsmän under Konanja och hans broder Simei, efter förordnande av konung Hiskia och Asarja, fursten i Guds hus.
Och leviten Kore, Jimnas son, som var dörrvaktare på östra sidan, hade uppsikten över de frivilliga gåvorna åt Gud och skulle fördela HERRENS offergärd och det högheliga av offren.
Och under honom sattes Eden, Minjamin, Jesua, Semaja, Amarja och Sekanja till förtroendemän i präststäderna för att ombesörja utdelningen åt sina bröder, efter deras avdelningar, åt den minste såväl som åt den störste.
Härifrån voro undantagna alla sådana i sina släktregister upptecknade personer av mankön, från tre års ålder och därutöver, som skulle infinna sig i HERRENS hus, där var dag de för den dagen bestämda sysslorna skulle utföras genom dem som hade tjänstgöringen, med de särskilda åligganden de hade efter sina avdelningar.
Och vad angick prästernas släktregister, så var det uppgjort efter deras familjer; och av leviterna voro de upptagna, som voro tjugu år gamla eller därutöver, efter sina särskilda åligganden, alltefter sina avdelningar.
Och i släktregistret skulle de vara upptecknade jämte alla sina späda barn, hustrur, söner och döttrar, så många de voro.
Ty på heder och tro skulle de förvalta det heliga såsom heligt.
Och för dem av Arons söner, prästerna, som bodde på sina städers utmarker, voro i var särskild stad namngivna män tillsatta, som åt allt mankön bland prästerna och åt alla de leviter som voro upptecknade i släktregistret skulle utdela vad dem tillkom.
Så förfor Hiskia i hela Juda, och han gjorde inför HERREN, sin Gud, vad gott och rätt och sant var.
Och allt som han företog sig, när han nu sökte sin Gud, allt, vare sig det angick tjänstgöringen i Guds hus eller det angick lagen och budorden, det gjorde han av allt sitt hjärta, och det lyckades honom väl.
Sedan han hade utfört detta och bevisat sådan trohet, kom Sanherib, konungen i Assyrien, och drog in i Juda och belägrade dess befästa städer och tänkte erövra dem åt sig.
Då nu Hiskia såg att Sanherib kom, i avsikt att belägra Jerusalem,
rådförde han sig med sina förnämsta män och sina hjältar om att täppa för vattnet i de källor som lågo utom staden; och de hjälpte honom härmed.
Mycket folk församlades och täppte till alla källorna och dämde för bäcken som flöt mitt igenom trakten, ty de sade: »När de assyriska konungarna komma, böra de icke finna vatten i sådan myckenhet.»
Och han tog mod till sig och byggde upp muren överallt där den var nedbruten, och byggde tornen högre, och förde upp en annan mur därutanför, och befäste Millo i Davids stad, och lät göra skjutvapen i myckenhet, så ock sköldar.
Och han tillsatte krigshövitsmän över folket och församlade dem till sig på den öppna platsen vid stadsporten, och talade uppmuntrande till dem och sade:
»Varen frimodiga och oförfärade, frukten icke och varen icke förskräckta för konungen i Assyrien och för hela den hop han har med sig; ty med oss är en som är större än den som är med honom.
Med honom är en arm av kött, men med oss är HERREN, vår Gud, och han skall hjälpa oss och föra våra krig.
Och folket tryggade sig vid Hiskias, Juda konungs, ord.
Därefter sände Sanherib, konungen i Assyrien -- som nu med hela sin härsmakt låg framför Lakis -- sina tjänare till Jerusalem, till Hiskia, Juda konung, och till alla dem av Juda, som voro i Jerusalem, och lät säga:
»Så säger Sanherib, konungen i Assyrien: Varpå förtrösten I, eftersom I stannen kvar i det belägrade Jerusalem?
Se, Hiskia uppeggar eder, så att I kommen att dö genom hunger och törst; han säger: 'HERREN, vår Gud, skall rädda oss ur den assyriske konungens hand.'
Har icke denne samme Hiskia avskaffat hans offerhöjder och altaren och sagt till Juda och Jerusalem: 'Inför ett enda altare skolen I tillbedja, och på detta skolen I tända offereld'?
Veten I icke vad jag och mina fäder hava gjort med andra länders alla folk?
Hava väl de gudar som dyrkas av folken i dessa andra länder någonsin förmått rädda sina länder ur min hand?
Ja, vilket bland alla dessa folk som mina fäder hava givit till spillo har väl haft någon gud som har förmått rädda sitt folk ur min hand eftersom I menen att eder Gud förmår rädda eder ur min hand!»
Nej, låten nu icke Hiskia så bedraga och uppegga eder, och tron honom icke; ty ingen gud hos något folk eller i något rike har förmått rädda sitt folk ur min hand eller ur mina fäders hand.
Huru mycket mindre skall då eder Gud kunna rädda eder ur min hand!»
Och hans tjänare talade ännu mer mot HERREN Gud och mot hans tjänare Hiskia.
Han hade ock skrivit ett brev vari han smädade HERREN, Israels Gud, och talade mot honom så: »Lika litet som de gudar som dyrkas av folken i de andra länderna hava kunnat rädda sina folk ur min hand, lika litet skall Hiskias Gud kunna rädda sitt folk ur min hand.»
Och till Jerusalems folk, dem som stodo på muren, ropade de med hög röst på judiska för att göra dem modlösa och förskräckta, så att man sedan skulle kunna intaga staden.
Och de talade om Jerusalems Gud på samma sätt som om de främmande folkens gudar, vilka äro verk av människohänder.
Men vid allt detta bådo konung Hiskia och profeten Jesaja, Amos' son, och ropade till himmelen.
Då sände HERREN en ängel, som förgjorde alla de tappra stridsmännen och furstarna och hövitsmännen i den assyriske konungens läger, så att han med skam måste draga tillbaka till sitt land.
Och när han en gång gick in i sin guds hus, blev han där nedhuggen med svärd av sina egna söner.
Så frälste HERREN Hiskia och Jerusalems invånare ur Sanheribs, den assyriske konungens, hand och ur alla andras hand; och han beskyddade dem på alla sidor.
Och många förde skänker till HERREN i Jerusalem och dyrbara gåvor till Hiskia, Juda konung; och han blev härefter högt aktad av alla folk.
Vid den tiden blev Hiskia dödssjuk.
Då bad han till HERREN, och han svarade honom och gav honom ett undertecken.
Dock återgäldade Hiskia icke det goda som hade blivit honom bevisat, utan hans hjärta blev högmodigt; därför kom förtörnelse över honom och över Juda och Jerusalem.
Men då Hiskia ödmjukade sig, mitt i sitt hjärtas högmod, och Jerusalems invånare med honom, drabbade HERRENS förtörnelse dem icke, så länge Hiskia levde.
Och Hiskias rikedom och härlighet var mycket stor; han hade byggt sig skattkamrar för silver och guld och ädla stenar, och för välluktande kryddor, och för sköldar och för allahanda dyrbara håvor av andra slag,
så ock förrådshus för vad som kom in av säd, vin och olja, ävensom stall för allt slags boskap; och hjordar hade han skaffat för sina fållor.
Och han hade byggt sig städer och förvärvat sig stor rikedom på får och fäkreatur; ty Gud hade givit honom mycket stora ägodelar.
Det var ock Hiskia som täppte till Gihonsvattnets övre källa och ledde vattnet nedåt, väster om Davids stad.
Och Hiskia var lyckosam i allt vad han företog sig.
Jämväl när från Babels furstar de sändebud kommo, som voro skickade till honom för att fråga efter det under som hade skett i landet, övergav Gud honom allenast för att pröva honom, på det att han skulle förnimma allt vad som var i hans hjärta.
Vad nu mer är att säga om Hiskia och om hans fromma gärningar, det finnes upptecknat i »Profeten Jesajas, Amos' sons, syner», i boken om Judas och Israels konungar.
Och Hiskia gick till vila hos sina fäder, och han begrov honom på den plats där man går upp till Davids hus' gravar; och hela Juda och Jerusalems invånare bevisade honom ära vid hans död.
Och hans son Manasse blev konung efter honom.
Manasse var tolv år gammal, när han blev konung, och han regerade femtiofem år i Jerusalem.
Han gjorde vad ont var i HERRENS ögon, efter den styggeliga seden hos de folk som HERREN hade fördrivit för Israels barn.
Han byggde åter upp de offerhöjder som hans fader Hiskia hade brutit ned, och reste altaren åt Baalerna och gjorde Aseror, och tillbad och tjänade himmelens hela härskara.
Ja, han byggde altaren i HERRENS hus, det om vilket HERREN hade sagt: »I Jerusalem skall mitt namn vara till evig tid.»
Han byggde altaren åt himmelens hela härskara på de båda förgårdarna till HERRENS hus.
Han lät ock sina barn gå genom eld i Hinnoms sons dal och övade teckentyderi, svartkonst och trolldom och skaffade sig andebesvärjare och spåmän och gjorde mycket som var ont i HERRENS ögon, så att han förtörnade honom.
Och avgudabelätet som han hade låtit göra satte han i Guds hus, om vilket Gud hade sagt till David och till hans son Salomo: »Vid detta hus och vid Jerusalem, som jag har utvalt bland alla Israels stammar, vill jag fästa mitt namn för evig tid.
Och jag skall icke mer låta Israel vandra bort ifrån det land som jag har bestämt åt edra fäder, om de allenast hålla och göra allt vad jag har bjudit dem, alldeles efter den lag, de stadgar och rätter som de hava fått genom Mose.»
Men Manasse förförde Juda och Jerusalems invånare, så att de gjorde mer ont än de folk som HERREN hade förgjort för Israels barn.
Och HERREN talade till Manasse och hans folk, men de aktade icke därpå.
Då lät HERREN den assyriske konungens härhövitsmän komma över dem; de slogo Manasse i bojor och fängslade honom med kopparfjättrar och förde honom till Babel.
Men när han nu var i nöd, bön föll han inför HERREN, sin Gud, och ödmjukade sig storligen för sina fäders Gud.
Och när han så bad till honom, lät han beveka sig och hörde hans bön och lät honom komma tillbaka till Jerusalem såsom konung.
Och då besinnade Manasse att HERREN är Gud.
Därefter byggde han en yttre mur till Davids stad västerut mot Gihon i dalen, intill Fiskporten, och runt omkring Ofel, och gjorde den mycket hög.
Och han insatte krigshövitsmän i alla befästa städer i Juda.
Och han skaffade bort de främmande gudarna och avgudabelätet ur HERRENS hus, så ock alla de altaren som han hade byggt på det berg där HERRENS hus stod och i Jerusalem, och kastade dem utanför staden.
Och han upprättade HERRENS altare och offrade tackoffer och lovoffer därpå, och uppmanade Juda att tjäna HERREN, Israels Gud.
Men folket offrade ännu på höjderna, dock allenast åt HERREN, sin Gud.
Vad nu mer är att säga om Manasse och om hans bön till sin Gud och om de ord som siarna talade till honom i HERRENS, Israels Guds, namn, det står i Israels konungars krönika.
Och om hans bön och huru han blev bönhörd, och om all hans synd och otrohet, och om de platser på vilka han byggde offerhöjder och ställde upp sina Aseror och beläten, innan han ödmjukade sig, härom är skrivet i Hosais krönika.
Och Manasse gick till vila hos sina fäder, och man begrov honom där han bodde.
Och hans son Amon blev konung efter honom.
Amon var tjugutvå år gammal, när han blev konung, och han regerade två år i Jerusalem.
Han gjorde vad ont var i HERRENS ögon, såsom hans fader Manasse hade gjort; åt alla de beläten som hans fader Manasse hade låtit göra offrade Amon, och han tjänade dem.
Men han ödmjukade sig icke för HERREN, såsom hans fader Manasse hade gjort, utan denne Amon hopade skuld på skuld.
Och hans tjänare sammansvuro sig mot honom och dödade honom hemma i hans hus.
Men folket i landet dräpte alla som hade sammansvurit sig mot konung Amon.
Därefter gjorde folket i landet hans son Josia till konung efter honom.
Josia var åtta år gammal, när han blev konung, och han regerade trettioett år i Jerusalem.
Han gjorde vad rätt var i HERRENS ögon och vandrade på sin fader Davids vägar och vek icke av vare sig till höger eller till vänster.
I sitt åttonde regeringsår, medan han ännu var en yngling, begynte han att söka sin fader Davids Gud; och i det tolfte året begynte han att rena Juda och Jerusalem från offerhöjderna och Aserorna och från de skurna och gjutna belätena.
Men Baalsaltarna brötos ned i hans åsyn, och solstoderna som voro uppställda på dem högg han ned, och Aserorna och de skurna och gjutna belätena slog han sönder och krossade dem till stoft och strödde ut stoftet på de mäns gravar, som hade offrat åt dem.
Och prästernas ben brände han upp på deras altaren.
Så renade han Juda och Jerusalem.
Och i Manasses, Efraims och Simeons städer ända till Naftali genomsökte han överallt husen.
Och sedan han hade brutit ned altarna och krossat Aserorna och belätena sönder till stoft och huggit ned alla solstoder i hela Israels land, vände han tillbaka till Jerusalem.
Och i sitt adertonde regeringsår, medan han höll på med att rena landet och templet, sände han Safan, Asaljas son, och Maaseja, hövitsmannen i staden, och kansleren Joa, Joahas' son, för att sätta HERRENS, sin Guds, hus i stånd.
Och de gingo till översteprästen Hilkia och avlämnade de penningar som hade influtit till Guds hus, sedan de av de leviter som höllo vakt vid tröskeln hade blivit insamlade från Manasse, Efraim och hela det övriga Israel, så ock från hela Juda och Benjamin och från Jerusalems invånare;
de överlämnade dem åt de män som förrättade arbete såsom tillsyningsmän vid HERRENS hus.
Sedan gåvos penningarna av dessa män, som förrättade arbete och hade befattning vid HERRENS hus med att laga huset och sätta det i stånd,
de gåvos åt timmermännen och byggningsmännen, till att inköpa huggen sten och trävirke till stockar, för att man därmed skulle timra upp de hus som Juda konungar hade förstört.
Och männen fingo vid sitt arbete handla på heder och tro; och tillsyningsmän över dem och föreståndare för arbetet voro Jahat och Obadja, leviter av Meraris barn, och Sakarja och Mesullam, av kehatiternas barn, så ock alla de leviter som voro kunniga på musikinstrumenter.
De hade ock tillsynen över bärarna, så att föreståndare funnos för alla arbetarna vid de särskilda göromålen.
Av leviterna togos ock skrivare, uppsyningsmän och dörrvaktare.
När de nu togo ut penningarna som hade influtit till HERRENS hus, fann prästen Hilkia HERRENS lagbok, den som hade blivit given genom Mose
Då tog Hilkia till orda och sade till sekreteraren Safan: »Jag har funnit lagboken i HERRENS hus.»
Och Hilkia gav boken åt Safan.
Och Safan bar boken till konungen och avgav därjämte sin berättelse inför konungen och sade: »Allt vad dina tjänare hava fått i uppdrag att göra, det göra de.
Och de hava tömt ut de penningar som funnos i HERRENS hus, och hava överlämnat dem åt tillsyningsmännen och åt arbetarna.»
Vidare berättade sekreteraren Safan för konungen och sade: »Prästen Hilkia har givit mig en bok.»
Och Safan föreläste därur för konungen
När konungen nu hörde lagens ord, rev han sönder sina kläder.
Och konungen bjöd Hilkia och Ahikam, Safans son, och Abdon, Mikas son, och sekreteraren Safan och Asaja, konungens tjänare, och sade:
»Gån och frågen HERREN för mig och för dem som äro kvar av Israel och Juda, angående det som står i den bok som nu har blivit funnen.
Ty stor är HERRENS vrede, den som är utgjuten över oss, därför att våra fäder icke hava hållit HERRENS ord och icke hava gjort allt som är föreskrivet i denna bok.»
Då gick Hilkia, tillika med andra som konungen sände åstad, till profetissan Hulda, hustru åt Sallum, klädkammarvaktaren, som var son till Tokehat, Hasras son; hon bodde i Jerusalem, i Nya staden.
Och de talade med henne såsom dem bjudet var.
Då svarade hon dem: »Så säger HERREN, Israels Gud: Sägen till den man som har sänt eder till mig:
Så säger HERREN: Se, över denna plats och över dess invånare skall jag låta olycka komma, alla de förbannelser som äro skrivna i den bok som man har föreläst för Juda konung --
detta därför att de hava övergivit mig och tänt offereld åt andra gudar, och så hava förtörnat mig med alla sina händers verk.
Min vrede skall utgjutas över denna plats och skall icke bliva utsläckt.
Men till Juda konung, som har sänt eder för att fråga HERREN, till honom skolen I säga så: Så säger HERREN, Israels Gud, angående de ord som du har hört:
Eftersom ditt hjärta blev bevekt och du ödmjukade dig inför Gud, när du hörde hans ord mot denna plats och mot dess invånare, ja, ödmjukade dig inför mig och rev sönder dina kläder och grät inför mig, fördenskull har jag ock hört dig, säger HERREN.
Se, jag vill samla dig till dina fäder, så att du får samlas till dem i din grav med frid, och dina ögon skola slippa att se all den olycka som jag skall låta komma över denna plats och dess invånare.»
Och de vände tillbaka till konungen med detta svar.
Då sände konungen åstad och lät församla alla de äldste i Juda och Jerusalem.
Och konungen gick upp i HERRENS hus med alla Juda män och Jerusalems invånare, också prästerna och leviterna, ja, allt folket, ifrån den störste till den minste.
Och han läste upp för dem allt vad som stod i förbundsboken, som hade blivit funnen i HERRENS hus.
Och konungen trädde fram på sin plats och slöt inför HERRENS ansikte det förbundet, att de skulle följa efter HERREN och hålla hans bud, hans vittnesbörd och hans stadgar, av allt sitt hjärta och av all sin själ, och göra efter förbundets ord, dem som voro skrivna i denna bok.
Och han lät alla som funnos i Jerusalem och Benjamin träda in i förbundet Och Jerusalems invånare gjorde efter Guds, sina fäders Guds, förbund.
Och Josia skaffade bort alla styggelser ur Israels barns alla landområden, och tillhöll alla dem som funnos i Israel att tjäna HERREN, sin Gud.
Så länge han levde, veko de icke av ifrån HERREN, sina fäders Gud.
Därefter höll Josia HERRENS påskhögtid i Jerusalem; man slaktade påskalammet på fjortonde dagen i första månaden.
Och han fastställde prästernas åligganden och styrkte dem till tjänstgöringen i HERRENS hus.
Och han sade till leviterna som undervisade hela Israel, och som voro helgade åt HERREN: »Sätten den heliga arken i det hus som Salomo, Davids son, Israels konung, har byggt.
Den skall icke mer vara en börda på edra axlar.
Tjänen nu HERREN, eder Gud, och hans folk Israel.
Gören eder redo efter edra familjer, i edra avdelningar, enligt vad David, Israels konung, har föreskrivit, och enligt hans son Salomos föreskrifter,
och inställen eder i helgedomen, ordnade efter edra bröders, det meniga folkets, familjeskiften, så att en avdelning av en levitisk familj kommer på vart skifte.
Och slakten påskalammet och helgen eder och reden till det för edra bröder, så att I gören efter HERRENS ord genom Mose.»
Och Josia gav åt det meniga folket såsom offergärd småboskap, dels lamm och dels killingar, till ett antal av trettio tusen, alltsammans till påskoffer, åt alla som voro där tillstädes, så ock tre tusen fäkreatur, detta allt av konungens enskilda egendom.
Och hans förnämsta män gåvo efter sin fria vilja offergåvor åt folket, åt prästerna och leviterna.
Hilkia, Sakarja och Jehiel, furstarna i Guds hus, gåvo åt prästerna två tusen sex hundra lamm och killingar till påskoffer, så ock tre hundra fäkreatur.
Men Konanja och hans bröder, Semaja och Netanel, jämte Hasabja, Jegiel och Josabad, de översta bland leviterna, gåvo åt leviterna såsom offergärd fem tusen lamm och killingar till påskoffer, så ock fem hundra fäkreatur.
Så blev det då ordnat för gudstjänsten; och prästerna inställde sig till tjänstgöring på sina platser och likaledes leviterna, efter sina avdelningar, såsom konungen hade bjudit.
Därefter slaktade de påskalammet, och prästerna stänkte med blodet som de togo emot av leviterna; och dessa drogo av huden.
Och de avskilde brännoffersstyckena och delade ut dem åt det meniga folket, efter deras familjeskiften, för att de skulle offra dem åt HERREN, såsom det var föreskrivet i Moses bok.
På samma sätt gjorde de ock med fäkreaturen.
Och de stekte påskalammet på eld, på föreskrivet sätt; men tackoffersköttet kokade de i grytor, pannor och kittlar och delade ut det med hast åt allt det meniga folket.
Sedan redde de till åt sig själva och åt prästerna; ty prästerna, Arons söner, voro upptagna ända till natten med att offra brännoffret och fettstyckena; därför måste leviterna reda till både åt sig och åt prästerna, Arons söner.
Och sångarna, Asafs barn, stodo på sin plats, såsom David och Asaf och Heman och konungens siare Jedutun hade bjudit, och dörrvaktarna stodo var och en vid sin port; de behövde icke gå ifrån sin tjänstgöring, ty deras bröder, de andra leviterna, redde till åt dem.
Så blev allt ordnat för HERRENS tjänst på den dagen, i det att man höll påskhögtid och offrade brännoffer på HERRENS altare, såsom konung Josia hade bjudit.
De israeliter som voro där tillstädes höllo nu påskhögtid och firade det osyrade brödets högtid i sju dagar.
En påskhögtid lik denna hade icke blivit hållen i Israel sedan profeten Samuels tid; ty ingen av Israels konungar hade hållit en sådan påskhögtid som den vilken nu hölls av Josia jämte prästerna och leviterna och hela Juda och dem av Israel, som voro där tillstädes, jämväl Jerusalems invånare.
I Josias adertonde regeringsår hölls denna påskhögtid.
Efter allt detta, sedan Josia hade försatt templet i gott stånd, drog Neko, konungen i Egypten, upp för att strida vid Karkemis, som ligger vid Frat; och Josia drog ut mot honom.
Då skickade denne sändebud till honom och lät säga: »Vad har du med mig att göra, du Juda konung?
Det är icke mot dig jag nu kommer, utan mot min arvfiende, och Gud har befallt mig att skynda.
Hör upp att trotsa Gud, som är med mig, och tag dig till vara, så att han icke fördärvar dig.»
Men i stället för att vända om och lämna honom i fred förklädde Josia sig och gick att strida mot honom, utan att höra på Nekos ord, som dock kommo från Guds mun.
Och det kom till strid på Megiddos slätt.
Men skyttarnas skott träffade konung Josia; och konungen sade till sina tjänare: »Bären mig undan, ty jag är svårt sårad.»
Då buro hans tjänare honom från stridsvagnen och satte honom i hans andra vagn och förde honom till Jerusalem; och han gav upp andan och blev begraven där hans fäder voro begravna.
Och hela Juda och Jerusalem sörjde Josia.
Och Jeremia sjöng en klagosång över Josia.
Och alla sångare och sångerskor talade sedan i sina klagosånger om Josia, såsom man gör ännu i dag; och dessa sånger blevo allmänt gängse i Israel.
De finnas upptecknade bland »Klagosångerna».
Vad nu mer är att säga om Josia och om de fromma gärningar han gjorde, efter vad föreskrivet var i HERRENS lag,
och om annat som han företog sig under sin första tid såväl som under sin sista, det finnes upptecknat i boken om Israels och Juda konungar
Och folket i landet tog Josias son Joahas och gjorde honom till konung i Jerusalem efter hans fader.
Joahas var tjugutre år gammal, när han blev konung, och han regerade tre månader i Jerusalem.
Konungen i Egypten avsatte honom i Jerusalem och pålade landet en skatt av ett hundra talenter silver och en talent guld.
Och konungen i Egypten gjorde hans broder Eljakim till konung över Juda och Jerusalem och förändrade hans namn till Jojakim men hans broder Joahas, honom tog Neko med sig, och han förde honom till Egypten.
Jojakim var tjugufem år gammal när han blev konung, och han regerade elva år i Jerusalem.
Han gjorde vad ont var i HERRENS, sin Guds, ögon.
Och Nebukadnessar, konungen i Babel, drog upp mot honom och fängslade honom med kopparfjättrar och förde honom bort till Babel.
Och en del av kärlen i HERRENS hus förde Nebukadnessar till Babel, och han satte in dem i sitt tempel i Babel.
Vad nu mer är att säga om Jojakim och om de styggelser som han gjorde, och om vad han eljest har befunnits vara skyldig till, det finnes upptecknat i boken om Israels och Juda konungar.
Och hans son Jojakin blev konung efter honom.
Jojakin var åtta år gammal, när han blev konung, och han regerade tre månader och tio dagar i Jerusalem.
Han gjorde vad ont var i HERRENS ögon.
Och vid följande års början sände konung Nebukadnessar och lät hämta honom till Babel, tillika med de dyrbara kärlen i HERRENS hus; och han gjorde hans broder Sidkia till konung över Juda och Jerusalem.
Sidkia var tjuguett år gammal, när han blev konung, och han regerade elva år i Jerusalem.
Han gjorde vad ont var i HERRENS, sin Guds, ögon; han ödmjukade sig icke för profeten Jeremia, som talade HERRENS ord.
Han avföll från konung Nebukadnessar, som hade tagit ed av honom vid Gud.
Och han var hårdnackad och förstockade sitt hjärta, så att han icke omvände sig till HERREN, Israels Gud.
Alla de översta bland prästerna och folket försyndade sig ock storligen i otrohet mot Gud med hedningarnas alla styggelser och orenade HERRENS hus, som han hade helgat i Jerusalem.
Och HERREN, deras faders Gud, skickade sina budskap till dem titt och ofta genom sina sändebud, ty han ömkade sig över sitt folk och sin boning.
Men de begabbade Guds sändebud och föraktade hans ord och bespottade hans profeter, till dess HERRENS vrede över hans folk växte så, att ingen bot mer fanns.
Då sände han emot dem kaldéernas konung, och denne dräpte deras unga män med svärd i deras helgedomshus och skonade varken ynglingar eller jungfrur, ej heller gamla och gråhårsmän; allt blev givet i hans hand.
Och alla kärl i Guds hus, både stora och små, och skatterna i HERRENS hus, så ock konungens och hans förnämsta mäns skatter, allt förde han till Babel.
Och man brände upp Guds hus och bröt ned Jerusalems mur, och alla dess palats brände man upp i eld och förstörde alla de dyrbara föremål som funnos där.
Och dem som hade undsluppit svärdet förde han bort i fångenskap till Babel, och de blevo tjänare åt honom och åt hans söner, till dess att perserna kommo till väldet --
för att HERRENS ord genom Jeremias mun skulle uppfyllas -- alltså till dess att landet hade fått gottgörelse för sina sabbater.
Ty medan det låg öde, hade det sabbat -- till dess att sjuttio år hade gått till ända.
Men i den persiske konungens Kores' första regeringsår uppväckte HERREN -- för att HERRENS ord genom Jeremias mun skulle fullbordas -- den persiske konungen Kores' ande, så att denne lät utropa över hela sitt rike och tillika skriftligen kungöra följande:
»Så säger Kores, konungen i Persien: Alla riken på jorden har HERREN, himmelens Gud, givit mig; och han har anbefallt mig att bygga honom ett hus i Jerusalem i Juda.
Vemhelst nu bland eder, som tillhör hans folk, med honom vare HERREN, hans Gud, och han drage ditupp.»
Men i den persiske konungen Kores' första regeringsår uppväckte HERREN -- för att HERRENS ord från Jeremias mun skulle fullbordas -- den persiske konungen Kores' ande, så att denne lät utropa över hela sitt rike och tillika skriftligen kungöra följande:
»Så säger Kores, konungen i Persien: Alla riken på jorden har HERREN, himmelens Gud, givit mig; och han har anbefallt mig att bygga honom ett hus i Jerusalem i Juda.
Vemhelst nu bland eder, som tillhör hans folk, med honom vare hans Gud, och han drage upp till Jerusalem i Juda för att bygga på HERRENS, Israels Guds, hus; han är den Gud som bor i Jerusalem.
Och varhelst någon ännu finnes kvar, må han av folket på den ort där han bor såsom främling få hjälp med silver och guld, med gods och boskap, detta jämte vad som frivilligt gives till Guds hus i Jerusalem.»
Då stodo huvudmännen för Judas och Benjamins familjer upp, ävensom prästerna och leviterna, alla de vilkas ande Gud uppväckte till att draga upp och bygga på HERRENS hus i Jerusalem.
Och alla de som bodde i deras grannskap understödde dem med silverkärl, med guld, med gods och boskap och med dyrbara skänker, detta förutom allt vad man eljest frivilligt gav.
Och konung Kores utlämnade de kärl till HERRENS hus, som Nebukadnessar hade fört bort ifrån Jerusalem och låtit sätta in i sin guds hus.
Dem utlämnade nu Kores, konungen i Persien, åt skattmästaren Mitredat, och denne räknade upp den åt Sesbassar, hövdingen för Juda.
Och detta var antalet av dem: trettio bäcken av guld, ett tusen bäcken av silver, tjugunio andra offerkärl,
trettio bägare av guld, fyra hundra tio silverbägare av ringare slag, därtill ett tusen andra kärl.
Kärlen av guld och silver utgjorde tillsammans fem tusen fyra hundra.
Allt detta förde Sesbassar med sig, när de som hade varit i fångenskapen drogo upp från Babel till Jerusalem.
Och dessa voro de män från hövdingdömet, som drogo upp ur den landsflykt och fångenskap i Babel, till vilken de hade blivit bortförda av Nebukadnessar, konungen i Babel, och som vände tillbaka till Jerusalem och Juda, var och en till sin stad,
i det att de följde med Serubbabel, Jesua, Nehemja, Seraja, Reelaja, Mordokai, Bilsan, Mispar, Bigvai, Rehum och Baana.
Detta var antalet män av Israels meniga folk:
Pareos' barn: två tusen ett hundra sjuttiotvå;
Sefatjas barn: tre hundra sjuttiotvå;
Aras barn: sju hundra sjuttiofem;
Pahat-Moabs barn, av Jesuas och Joabs barn: två tusen åtta hundra tolv;
Elams barn: ett tusen två hundra femtiofyra;
Sattus barn: nio hundra fyrtiofem;
Sackais barn: sju hundra sextio;
Banis barn: sex hundra fyrtiotvå;
Bebais barn: sex hundra tjugutre;
Asgads barn: ett tusen två hundra tjugutvå;
Adonikams barn: sex hundra sextiosex;
Bigvais barn: två tusen femtiosex;
Adins barn: fyra hundra femtiofyra;
Aters barn av Hiskia: nittioåtta;
Besais barn: tre hundra tjugutre;
Joras barn: ett hundra tolv;
Hasums barn: två hundra tjugutre;
Gibbars barn: nittiofem;
Bet-Lehems barn: ett hundra tjugutre;
männen från Netofa: femtiosex;
männen från Anatot: ett hundra tjuguåtta;
Asmavets barn: fyrtiotvå;
Kirjat-Arims, Kefiras och Beerots barn: sju hundra fyrtiotre;
Ramas och Gebas barn: sex hundra tjuguen;
männen från Mikmas: ett hundra tjugutvå;
männen från Betel och Ai: två hundra tjugutre;
Nebos barn: femtiotvå;
Magbis' barn: ett hundra femtiosex;
den andre Elams barn: ett tusen två hundra femtiofyra;
Harims barn: tre hundra tjugu;
Lods, Hadids och Onos barn: sju hundra tjugufem;
Jerikos barn: tre hundra fyrtiofem;
Senaas barn: tre tusen sex hundra trettio.
Av prästerna: Jedajas barn av Jesuas hus: nio hundra sjuttiotre;
Immers barn: ett tusen femtiotvå;
Pashurs barn: ett tusen två hundra fyrtiosju;
Harims barn: ett tusen sjutton.
Av leviterna: Jesuas och Kadmiels barn, av Hodaujas barn: sjuttiofyra;
av sångarna: Asafs barn: ett hundra tjuguåtta;
av dörrvaktarnas barn: Sallums barn, Aters barn, Talmons barn, Ackubs barn, Hatitas barn, Sobais barn: alla tillsammans ett hundra trettionio.
Av tempelträlarna: Sihas barn, Hasufas barn, Tabbaots barn,
Keros' barn, Siahas barn, Padons barn,
Lebanas barn, Hagabas barn, Ackubs barn,
Hagabs barn, Samlais barn, Hanans barn,
Giddels barn, Gahars barn, Reajas barn,
Resins barn, Nekodas barn, Gassams barn,
Ussas barn, Paseas barn, Besais barn,
Asnas barn, Meunims barn, Nefisims barn,
Bakbuks barn, Hakufas barn, Harhurs barn,
Basluts barn, Mehidas barn, Harsas barn,
Barkos' barn, Siseras barn, Temas barn,
Nesias barn, Hatifas barn.
Av Salomos tjänares barn: Sotais barn, Hassoferets barn, Perudas barn,
Jaalas barn, Darkons barn, Giddels barn,
Sefatjas barn, Hattils barn, Pokeret-Hassebaims barn, Amis barn.
Tempelträlarna och Salomos tjänares barn utgjorde tillsammans tre hundra nittiotvå.
Och dessa voro de som drogo åstad från Tel-Mela, Tel-Harsa, Kerub, Addan och Immer, men som icke kunde uppgiva sina familjer och sin släkt och huruvida de voro av Israel:
Delajas barn, Tobias barn, Nekodas barn, sex hundra femtiotvå.
Och av prästernas barn: Habajas barn, Hackos' barn, Barsillais barn, hans som tog en av gileaditen Barsillais döttrar till hustru och blev uppkallad efter deras namn.
Dessa sökte efter sina släktregister, men kunde icke finna dem; därför blevo de såsom ovärdiga uteslutna från prästadömet.
Och ståthållaren tillsade dem att de icke skulle få äta av det högheliga, förrän en präst uppstode med urim och tummim.
Hela församlingen utgjorde sammanräknad fyrtiotvå tusen tre hundra sextio,
förutom deras tjänare och tjänarinnor, som voro sju tusen tre hundra trettiosju.
Och till dem hörde två hundra sångare och sångerskor.
De hade sju hundra trettiosex hästar, två hundra fyrtiofem mulåsnor,
fyra hundra trettiofem kameler och sex tusen sju hundra tjugu åsnor.
Och somliga av huvudmännen för familjerna gåvo, när de kommo till HERRENS hus i Jerusalem, frivilliga gåvor till Guds hus, för att det åter skulle byggas upp på samma plats.
De gåvo, efter som var och en förmådde, till arbetskassan i guld sextioett tusen dariker och i silver fem tusen minor, så ock ett hundra prästerliga livklädnader.
Och prästerna, leviterna, en del av meniga folket, sångarna, dörrvaktarna och tempelträlarna bosatte sig i sina städer: hela Israel i sina städer.
När sjunde månaden nalkades och Israels barn nu voro bosatta i sina städer, församlade sig folket såsom en man till Jerusalem.
Och Jesua, Josadaks son, och hans bröder, prästerna, och Serubbabel, Sealtiels son, och hans bröder stodo upp och byggde Israels Guds altare för att offra brännoffer därpå, såsom det var föreskrivet i gudsmannen Moses lag.
De uppförde altaret på dess plats, ty en förskräckelse hade kommit över dem för de främmande folken; och de offrade åt HERREN brännoffer därpå, morgonens och aftonens brännoffer.
Och de höllo lövhyddohögtiden, såsom det var föreskrivet, och offrade brännoffer för var dag till bestämt antal, på stadgat sätt, var dag det för den dagen bestämda antalet,
och därefter det dagliga brännoffret och de offer som hörde till nymånaderna och till alla HERRENS övriga helgade högtider, så ock alla de offer som man frivilligt frambar åt HERREN.
På första dagen i sjunde månaden begynte de att offra brännoffer åt HERREN, innan grunden till HERRENS tempel ännu var lagd.
Och de gåvo penningar åt stenhuggare och timmermän, så ock matvaror, dryckesvaror och olja åt sidonierna och tyrierna, för att dessa sjöledes skulle föra cederträ från Libanon till Jafo, i enlighet med den tillåtelse som Kores, konungen i Persien, hade givit dem.
Och året näst efter det då de hade kommit till Guds hus i Jerusalem, i andra månaden, begyntes verket av Serubbabel, Sealtiels son, och Jesua, Josadaks son, och deras övriga bröder, prästerna och leviterna, och av alla dem som ur fångenskapen hade kommit till Jerusalem; det begyntes därmed att de anställde leviterna, dem som voro tjugu år gamla eller därutöver, till att förestå arbetet på HERRENS hus.
Och Jesua med sina söner och bröder och Kadmiel med sina söner, Judas söner, allasammans, blevo anställda till att hava uppsikt över dem som utförde arbetet på Guds hus, sammaledes ock Henadads söner med sina söner och bröder, leviterna.
Och när byggningsmännen lade grunden till HERRENS tempel, ställdes prästerna upp i ämbetsskrud med trumpeter, så ock leviterna, Asafs barn, med cymbaler, till att lova HERREN, efter Davids, Israels konungs, anordning.
Och de sjöngo, under lov och tack till HERREN, därför att han är god, och därför att hans nåd varar evinnerligen över Israel.
Och allt folket jublade högt till HERRENS lov, därför att grunden till HERRENS hus var lagd.
Men många av prästerna och leviterna och huvudmännen för familjerna, de gamle som hade sett det förra huset, gräto högljutt, när de sågo grunden läggas till detta hus, många åter jublade och voro så glada att de ropade med hög röst.
Och man kunde icke skilja mellan det högljudda, glada jubelropet och folkets högljudda gråt; ty folket ropade så högt att ljudet därav hördes vida omkring.
Men när ovännerna till Juda och Benjamin fingo höra att de som hade återkommit ifrån fångenskapen höllo på att bygga ett tempel åt HERREN, Israels Gud,
gingo de till Serubbabel och till huvudmännen för familjerna och sade till dem: »Vi vilja bygga tillsammans med eder, ty vi söka eder Gud, likasom I, och åt honom offra vi alltsedan den tid då den assyriske konungen Esarhaddon lät föra oss hit.»
Men Serubbabel och Jesua och de övriga huvudmännen för Israels familjer sade till dem: »Det är icke tillbörligt att I tillsammans med oss byggen ett hus åt vår Gud, utan vi vilja för oss själva med varandra bygga huset åt HERREN, Israels Gud, såsom konung Kores, konungen i Persien, har bjudit oss.»
Men folket i landet bedrev det så, att judafolkets mod föll och de avskräcktes från att bygga vidare.
Och de lejde mot dem män som genom sina råd gjorde deras rådslag om intet, så länge Kores, konungen i Persien, levde, och sedan ända till dess att Darejaves, konungen i Persien, kom till regeringen.
(Sedermera, under Ahasveros' regering, redan i begynnelsen av hans regering, skrev man en anklagelseskrift mot dem som bodde i Juda och Jerusalem.
Och i Artasastas tid skrevo Bislam, Mitredat och Tabeel samt dennes övriga medbröder till Artasasta, konungen i Persien.
Och det som stod i skrivelsen var skrivet med arameiska bokstäver och avfattat på arameiska.
Likaledes skrevo rådsherren Rehum och sekreteraren Simsai ett brev om Jerusalem till konung Artasasta av följande innehåll.
De skrevo då, rådsherren Rehum och sekreteraren Simsai och de andra, deras medbröder: diniterna och afaresatkiterna, tarpeliterna, afaresiterna, arkeviterna, babylonierna, susaniterna, dehaviterna, elamiterna
och de andra folk som den store och mäktige Asenappar hade fört bort och låtit bosätta sig i staden Samaria och annorstädes i landet på andra sidan floden o. s. v.
Och detta är vad som stod skrivet i det brev som de sände till konung Artasasta: »Dina tjänare, männen på andra sidan floden o. s. v.
Det vare veterligt för konungen att de judar som drogo upp från dig hava kommit hit till oss i Jerusalem, och de hålla nu på att bygga upp den upproriska och onda staden, att sätta murarna i stånd och att förbättra grundvalarna.
Så må nu konungen veta, att om denna stad bliver uppbyggd och murarna bliva satta i stånd, skola de varken giva skatt eller tull eller vägpenningar, och sådant skall bliva till men för konungarnas inkomster.
Alldenstund vi nu äta palatsets salt, och det icke är tillbörligt att vi åse huru skada tillskyndas konungen, därför sända vi nu och låta konungen veta detta,
för att man må göra efterforskningar i dina fäders krönikor; ty av dessa krönikor skall du finna och erfara att denna stad har varit en upprorisk stad, till förfång för konungar och länder, och att man i den har anstiftat oroligheter ända ifrån äldsta tider, varför ock denna stad har blivit förstörd.
Så låta vi nu konungen veta, att om denna stad bliver uppbyggd och dess murar bliva satta i stånd, så skall du i följd härav icke mer hava någon del i landet på andra sidan floden.»
Då sände konungen följande svar till rådsherren Rehum och sekreteraren Simsai och de andra, deras medbröder, som bodde i Samaria och i det övriga landet på andra sidan floden: »Frid o. s. v.
Den skrivelse som I haven sänt till oss har noggrant blivit uppläst för mig.
Och sedan jag hade givit befallning att man skulle göra efterforskningar, fann man att denna stad ända ifrån äldsta tider har plägat sätta sig upp mot konungar, och att uppror och oroligheter där hava anstiftats.
I Jerusalem hava ock funnits mäktiga konungar, som hava varit herrar över allt land som ligger på andra sidan floden, och skatt, tull och vägpenningar hava blivit dem givna.
Så utfärden nu en befallning att man förhindrar dessa män att bygga upp denna stad, till dess jag giver befallning därom.
Och sen till, att I icke handlen försumligt i denna sak, så att skadan icke växer, konungarna till förfång.»
Så snart nu vad som stod i konung Artasastas skrivelse hade blivit läst för Rehum och sekreteraren Simsai och deras medbröder, gingo de med hast till judarna i Jerusalem och hindrade dem med våld och makt.)
Så förhindrades nu arbetet på Guds hus i Jerusalem.
Och det blev förhindrat ända till den persiske konungen Darejaves' andra regeringsår.
Men profeten Haggai och Sakarja, Iddos son, profeterna, profeterade för judarna i Juda och Jerusalem, i Israels Guds namn, efter vilket de voro uppkallade.
Och Serubbabel, Sealtiels son, och Jesua, Josadaks son, stodo då upp och begynte bygga på Guds hus i Jerusalem, och med dem Guds profeter, som understödde dem.
Vid samma tid kommo till dem Tattenai, ståthållaren i landet på andra sidan floden, och Setar-Bosenai och dessas medbröder, och sade så till dem: »Vem har givit eder tillåtelse att bygga detta hus och att sätta denna mur i stånd?»
Då sade vi dem vad de män hette, som uppförde byggnaden.
Och över judarnas äldste vakade deras Guds öga, så att man lovade att icke lägga något hinder i vägen för dem, till dess saken hade kommit inför Darejaves; sedan skulle man sända dem en skrivelse härom.
Detta är nu vad som stod skrivet i det brev som Tattenai, ståthållaren i landet på andra sidan floden, och Setar-Bosenai och hans medbröder, afarsekiterna, som bodde på andra sidan floden, sände till konung Darejaves;
de sände nämligen till honom en berättelse, och däri var så skrivet: »Frid vare i allo med konung Darejaves.
Det vare veterligt för konungen att vi kommo till det judiska hövdingdömet, till den store Gudens hus.
Detta håller man nu på att bygga upp med stora stenar, och i väggarna lägger man in trävirke; och arbetet bedrives med omsorg och har god framgång under deras händer.
Då frågade vi de äldste där och sade till dem så: 'Vem har givit eder tillåtelse att bygga detta hus och att sätta denna mur i stånd?'
Vi frågade dem ock huru de hette, för att kunna underrätta dig därom, och för att teckna upp namnen på de män som stodo i spetsen för dem.
Och detta var det svar som de gåvo oss: 'Vi äro himmelens och jordens Guds tjänare, och vi bygga nu upp det hus som fordom, för många år sedan, var uppbyggt här, och som en stor konung i Israel hade byggt och fulländat.
Men eftersom våra fäder förtörnade himmelens Gud, gav han dem i kaldéen Nebukadnessars, den babyloniske konungens, hand; och han förstörde detta hus och förde folket bort till Babel.
Men i den babyloniske konungen Kores' första regeringsår gav konung Kores befallning att man åter skulle bygga upp detta Guds hus.
Och tillika tog konung Kores ur templet i Babel de kärl av guld och silver, som hade tillhört Guds hus, men som Nebukadnessar hade tagit ur templet i Jerusalem och fört till templet i Babel; och de överlämnades åt en man vid namn Sesbassar, som han hade satt till ståthållare.
Och till honom sade han: Tag dessa kärl och far åstad och sätt in dem i templet i Jerusalem; ty Guds hus skall åter byggas upp på sin plats.
Så kom då denne Sesbassar hit och lade grunden till Guds hus i Jerusalem.
Och från den tiden och intill nu har man byggt därpå, och det är ännu icke färdigt.'
Om det nu täckes konungen, må man göra efterforskningar i konungens skattkammare därborta i Babel om det är så, att konung Kores har givit tillåtelse att bygga detta Guds hus i Jerusalem; därefter må konungen meddela oss sin vilja härom.»
Då gav konung Darejaves befallning att man skulle göra efterforskningar i kansliet i Babel, där skatterna nedlades.
Och i Ametas borg, i hövdingdömet Medien, fann man en bokrulle i vilken följande var upptecknat till hågkomst:
»I konung Kores' första regeringsår gav konung Kores denna befallning: 'Guds hus i Jerusalem, det huset skall byggas upp till att vara en plats där man frambär offer; och dess grundvalar skola göras fasta.
Det skall byggas sextio alnar högt och sextio alnar brett,
med tre varv stora stenar och med ett varv nytt trävirke; och vad som fordras för omkostnaderna skall utgivas från konungens hus.
De kärl av guld och silver i Guds hus, som Nebukadnessar tog ur templet i Jerusalem och förde till Babel, skall man ock giva tillbaka, så att de komma åter till sin plats i templet i Jerusalem, och man skall sätta in dem i Guds hus.' --
Alltså, du Tattenai, som är ståthållare i landet på andra sidan floden, och du Setar-Bosenai, och I afarsekiter, de nämndas medbröder på andra sidan floden: hållen eder fjärran därifrån.
Lämnen arbetet på detta Guds hus ostört.
Judarnas ståthållare och judarnas äldste må bygga detta Guds hus på dess plats.
Och härmed giver jag befallning om huru I skolen förfara med dessa judarnas äldste, när de bygga på detta Guds hus.
Av de penningar som givas åt konungen i skatt från landet på andra sidan floden skall vad som fordras för omkostnaderna redligt utgivas åt dessa män, så att hinder icke uppstår i arbetet.
Och vad de behöva, ungtjurar, vädurar och lamm till brännoffer åt himmelens Gud, så och vete, salt, vin och olja, det skall, efter uppgift av prästerna i Jerusalem, utgivas åt dem dag för dag utan någon försummelse,
för att de må kunna frambära offer, till en välbehaglig lukt åt himmelens Gud, och för att de må bedja för konungens och hans söners liv.
Och härmed giver jag befallning, att om någon överträder denna förordning, så skall en bjälke brytas ut ur hans hus, och på den skall man upphänga och fästa honom, och hans hus skall göras till en plats för orenlighet, därför att han har så gjort.
Och må den Gud som har låtit sitt namn bo där slå ned alla konungar och folk som uträcka sin hand till att överträda denna förordning, och till att förstöra detta Guds hus i Jerusalem.
Jag, Darejaves, giver denna befallning.
Blive den redligt fullgjord!»
Alldenstund nu konung Darejaves hade sänt ett sådant bud, blev detta redligt fullgjort av Tattenai, ståthållaren i landet på andra sidan floden, och av Setar-Bosenai, så ock av deras medbröder.
Och judarnas äldste byggde vidare och hade god framgång i arbetet genom profeten Haggais och Sakarjas, Iddos sons, profetiska tal; man byggde och fullbordade det såsom Israels Gud hade befallt, och såsom Kores och Darejaves och Artasasta, den persiske konungen, hade befallt.
Och huset blev färdigt till den tredje dagen i månaden Adar, i konung Darejaves' sjätte regeringsår.
Och Israels barn, prästerna och leviterna och de övriga som hade återkommit ifrån fångenskapen, firade invigningen av detta Guds hus med glädje.
Och till invigningen av detta Guds hus offrade de ett hundra tjurar, två hundra vädurar och fyra hundra lamm, så ock till syndoffer för hela Israel tolv bockar, efter antalet av Israels stammar.
Och man anställde prästerna, efter deras skiften, och leviterna, efter deras avdelningar, till att förrätta Guds tjänst i Jerusalem, såsom det var föreskrivet i Moses bok.
Och de som hade återkommit ifrån fångenskapen höllo påskhögtid på fjortonde dagen i första månaden.
Ty prästerna och leviterna hade då allasammans renat sig, så att de alla voro rena; och de slaktade påskalammet för alla dem som hade återkommit ifrån fångenskapen, också för sina bröder, prästerna, likasåväl som för sig själva.
Och de israeliter som hade återvänt ifrån fångenskapen åto därav, jämte alla sådana som hade avskilt sig från den hedniska landsbefolkningens orenhet och slutit sig till dem för att söka HERREN, Israels Gud.
Och de höllo det osyrade brödets högtid i sju dagar med glädje; ty HERREN hade berett dem glädje, i det att han hade vänt den assyriske konungens hjärta till dem, så att han understödde dem i arbetet på Guds, Israels Guds, hus.
Efter en tids förlopp, under den persiske konungen Artasastas regering, hände sig att Esra, son till Seraja, son till Asarja, son till Hilkia,
son till Sallum, son till Sadok, son till Ahitub,
son till Amarja, son till Asarja, son till Merajot,
son till Seraja, son till Ussi, son till Bucki,
son till Abisua, son till Pinehas, son till Eleasar, son till Aron, översteprästen --
det hände sig att denne Esra drog upp från Babel; han var en skriftlärd, väl förfaren i Moses lag, den som HERREN, Israels Gud, hade utgivit.
Och konungen gav honom allt vad han begärde, eftersom HERRENS, hans Guds, hand var över honom.
Också en del av Israels barn och av prästerna, leviterna, sångarna, dörrvaktarna och tempelträlarna drog upp till Jerusalem i Artasastas sjunde regeringsår.
Och han kom till Jerusalem i femte månaden, i konungens sjunde regeringsår.
Ty på första dagen i första månaden blev det bestämt att man skulle draga upp från Babel; och på första dagen i femte månaden kom han till Jerusalem, eftersom Guds goda hand var över honom.
Ty Esra hade vänt sitt hjärta till att begrunda HERRENS lag och göra efter den, och till att i Israel undervisa i lag och rätt.
Så stod nu skrivet i den skrivelse som konung Artasasta gav åt prästen Esra, den skriftlärde, som var lärd i det som HERREN hade bjudit och stadgat för Israel:
»Artasasta, konungarnas konung, till prästen Esra, den i himmelens Guds lag lärde, o. s. v. med övlig fortsättning.
Jag giver härmed befallning att var och en i mitt rike av Israels folk och av dess präster och leviter, som är villig att fara till Jerusalem, må fara med dig,
alldenstund du är sänd av konungen och hans sju rådgivare till att hålla undersökning om Juda och Jerusalem efter din Guds lag, som är i din hand,
och till att föra dit det silver och guld som konungen och hans rådgivare av fritt beslut hava givit åt Israels Gud, vilken har sin boning i Jerusalem,
så ock allt det silver och guld som du kan få i hela Babels hövdingdöme, tillika med de frivilliga gåvor som folket och prästerna giva till sin Guds hus i Jerusalem.
Alltså skall du nu för dessa penningar såsom en redlig man köpa tjurar, vädurar och lamm, jämte sådant som behöves till dithörande spisoffer och drickoffer; och detta skall du offra på altaret i eder Guds hus i Jerusalem.
Och vad du och dina bröder finnen för gott att göra med det silver och guld som bliver över, det mån I göra efter eder Guds vilja.
Och alla de kärl som givas dig till tempeltjänsten i din Guds hus skall du avlämna inför Jerusalems Gud.
Och vad du måste utbetala för det som härutöver behöves till din Guds hus, det må du låta utbetala ur konungens skattkammare.
Och jag, konung Artasasta, giver härmed befallning till alla skattmästare i landet på andra sidan floden att allt vad prästen Esra, den i himmelens Guds lag lärde, begär av eder, det skall redligt göras och givas,
ända till hundra talenter silver, hundra korer vete, hundra bat vin och hundra bat olja, så ock salt utan särskild föreskrift.
Allt vad himmelens Gud befaller skall noggrant göras och givas till himmelens Guds hus, för att icke vrede må komma över konungens och hans söners rike.
Och vi göra eder veterligt att ingen skall hava makt att lägga skatt, tull eller vägpenningar på någon präst eller levit, sångare, dörrvaktare, tempelträl eller annan tjänare i detta Guds hus.
Och du, Esra, må, efter din Guds vishet, den som har blivit dig betrodd, förordna domare och lagkloke till att döma allt folket i landet på andra sidan floden, alla dem som känna din Guds lagar; och om någon icke känner dessa, skolen I lära honom dem.
Och var och en som icke gör efter din Guds lag och konungens lag, över honom skall dom fällas med rättvisa, vare sig till död eller till landsförvisning eller till penningböter eller till fängelse.»
Lovad vare HERREN, våra fäders Gud, som ingav konungen sådant i hjärtat, nämligen att han skulle förhärliga HERRENS hus i Jerusalem,
och som lät mig finna nåd inför konungen och hans rådgivare och inför alla konungens mäktiga hövdingar!
Och jag kände mig frimodig, eftersom HERRENS, min Guds, hand var över mig, och jag församlade en del av huvudmännen i Israel till att draga upp med mig.
Och dessa voro de huvudmän för familjerna, som under konung Artasastas regering med mig drogo upp från Babel, och så förhöll det sig med deras släkter:
Av Pinehas' barn Gersom; av Itamars barn Daniel; av Davids barn Hattus;
av Sekanjas barn, av Pareos' barn, Sakarja och med honom i släktregistret upptagna män, ett hundra femtio;
av Pahat-Moabs barn Eljoenai, Serajas son, och med honom två hundra män;
av Sekanjas barn Jahasiels son och med honom tre hundra män;
av Adins barn Ebed, Jonatans son, och med honom femtio män;
av Elams barn Jesaja, Ataljas son, och med honom sjuttio män;
av Sefatjas barn Sebadja, Mikaels son, och med honom åttio män;
av Joabs barn Obadja, Jehiels son och med honom två hundra aderton män;
av Selomits barn Josifjas son och med honom ett hundra sextio män;
av Bebais barn Sakarja, Bebais son, och med honom tjuguåtta män;
av Asgads barn Johanan, Hackatans son, och med honom ett hundra tio män;
av Adonikams barn de sistkomna, vilka hette Elifelet, Jegiel och Semaja, och med dem sextio män;
av Bigvais barn Utai och Sabbud och med dem sjuttio män.
Och jag församlade dessa till den ström som flyter till Ahava, och vi voro lägrade där i tre dagar.
Men när jag närmare gav akt på folket och prästerna, fann jag där ingen av Levi barn.
Då sände jag åstad huvudmännen Elieser, Ariel, Semaja, Elnatan, Jarib, Elnatan, Natan, Sakarja och Mesullam och lärarna Jojarib och Elnatan;
jag bjöd dem gå till Iddo, huvudmannen i Kasifja, och jag lade dem i munnen de ord som de skulle tala till Iddo och hans broder och till tempelträlarna i Kasifja, på det att man skulle sända till oss tjänare för vår Guds hus.
Och eftersom vår Guds goda hand var över oss, sände de till oss en förståndig man av Mahelis, Levis sons, Israels sons, barn, ävensom Serebja med hans söner och bröder, aderton män,
vidare Hasabja och med honom Jesaja, av Meraris barn, med dennes bröder och deras söner, tjugu män,
så ock två hundra tjugu tempelträlar, alla namngivna, av de tempelträlar som David och hans förnämsta män hade givit till leviternas tjänst.
Och jag lät där, vid Ahavaströmmen, lysa ut en fasta, för att vi skulle ödmjuka oss inför vår Gud, till att av honom utbedja oss en lyckosam resa för oss och våra kvinnor och barn och all vår egendom.
Ty jag blygdes för att av konungen begära krigsfolk och ryttare till att hjälpa oss mot fiender på vägen, eftersom vi hade sagt till konungen: »Vår Guds hand är över alla dem som söka honom, och så går det dem väl, men hans makt och hans vrede äro emot alla dem som övergiva honom.»
Därför fastade vi och sökte hjälp av vår Gud, och han bönhörde oss.
Och jag avskilde tolv av de översta bland prästerna, så ock Serebja och Hasabja och med dem tio av deras bröder.
Och jag vägde upp åt dem silvret och guldet och kärlen, den gärd till vår Guds hus, som hade blivit given av konungen och hans rådgivare och hövdingar och av alla de israeliter som voro där.
Jag vägde upp åt dem sex hundra femtio talenter silver jämte silverkärl till ett värde av ett hundra talenter, så ock ett hundra talenter guld,
därtill tjugu bägare av guld, till ett värde av tusen dariker, samt två kärl av fin, glänsande koppar, dyrbara såsom guld.
Och jag sade till dem: »I ären helgade åt HERREN, och kärlen äro helgade, och silvret och guldet är en frivillig gåva åt HERREN, edra fäders Gud.
Så vaken däröver och bevaren det, till dess I fån väga upp det i Jerusalem inför de översta bland prästerna och leviterna och de översta inom Israels familjer, i kamrarna i HERRENS hus.»
Då togo prästerna och leviterna emot det uppvägda, silvret och guldet och kärlen, för att de skulle föra det till Jerusalem, till vår Guds hus.
Och vi bröto upp från Ahavaströmmen på tolfte dagen i första månaden för att draga till Jerusalem; och vår Guds hand var över oss och räddade oss undan fiender och försåt på vägen.
Och vi kommo till Jerusalem och blevo stilla där i tre dagar.
Men på fjärde dagen uppvägdes silvret och guldet och kärlen i vår Guds hus, och överlämnades åt prästen Meremot, Urias son, och jämte honom åt Eleasar, Pinehas' son, och jämte dessa åt leviterna Josabad, Jesuas son, och Noadja, Binnuis som --
alltsammans efter antal och vikt, och hela vikten blev då upptecknad.
De landsflyktiga som hade återkommit ifrån fångenskapen offrade nu till brännoffer åt Israels Gud tolv tjurar för hela Israel, nittiosex vädurar, sjuttiosju lamm och tolv syndoffersbockar, alltsammans till brännoffer åt HERREN.
Och de överlämnade konungens påbud åt konungens satraper och åt ståthållarna i landet på andra sidan floden, och dessa gåvo understöd åt folket och åt Guds hus.
Sedan allt detta hade skett, trädde några av furstarna fram till mig och sade: »Varken folket i Israel eller prästerna och leviterna hava hållit sig avskilda från de främmande folken, såsom tillbörligt hade varit för de styggelsers skull som hava bedrivits av dem, av kananéerna, hetiterna, perisséerna, jebuséerna, ammoniterna, moabiterna, egyptierna och amoréerna.
Ty av deras döttrar hava de tagit hustrur åt sig och åt sina söner, och så har det heliga släktet blandat sig med de främmande folken; och furstarna och föreståndarna hava varit de första att begå sådan otrohet.»
När jag nu hörde detta, rev jag sönder min livrock och min kåpa och ryckte av mig huvudhår och skägg och blev sittande i djup sorg.
Och alla de som fruktade för vad Israels Gud hade talat mot sådan otrohet som den de återkomna fångarna hade begått, de församlade sig till mig, under det att jag förblev sittande i min djupa sorg ända till tiden för aftonoffret.
Men vid tiden för aftonoffret stod jag upp från min bedrövelse och rev sönder min livrock och min kåpa; därefter föll jag ned på mina knän och uträckte mina händer till HERREN, min Gud,
och sade: »Min Gud, jag skämmes och blyges för att upplyfta mitt ansikte till dig, min Gud, ty våra missgärningar hava växt oss över huvudet, och vår skuld är stor allt upp till himmelen.
Från våra fäders dagar ända till denna dag hava vi varit i stor skuld, och genom våra missgärningar hava vi, med våra konungar och präster, blivit givna i främmande konungars hand, och hava drabbats av svärd, fångenskap, plundring och skam, såsom det går oss ännu i dag.
Men nu har ett litet ögonblick nåd vederfarits oss från HERREN, vår Gud, så att han har låtit en räddad skara bliva kvar av oss, och givit oss fotfäste på sin heliga plats, för att han, vår Gud, så skulle låta ljus gå upp för våra ögon och giva oss något litet andrum i vår träldom.
Ty trälar äro vi, men i vår träldom har vår Gud icke övergivit oss, utan han har låtit oss finna nåd inför Persiens konungar, så att de hava givit oss andrum till att upprätta vår Guds hus och bygga upp dess ruiner och bereda oss en hägnad plats i Juda och Jerusalem.
Och vad skola vi nu säga, o vår Gud, efter allt detta?
Vi hava ju övergivit dina bud,
dem som du gav genom dina tjänare profeterna, i det du sade: 'Det land dit I nu kommen, för att taga det i besittning, är ett besmittat land, genom de främmande folkens besmittelse, och genom de styggelser med vilka de i sin orenhet hava uppfyllt det från den ena ändan till den andra.
Så given nu icke edra döttrar åt deras söner, och tagen icke deras döttrar till hustrur åt edra söner.
Ja, I skolen aldrig fråga efter deras välfärd och lycka -- detta på det att I mån bliva starka, så att I fån äta av landets goda och lämna det till besittning åt edra barn för evärdlig tid.'
Skulle vi väl nu, efter allt vad som har kommit över oss genom våra onda gärningar och genom den stora skuld vi hava ådragit oss, och sedan du, vår Gud, har skonat oss mer än våra missgärningar förtjänade, och låtit en skara av oss, sådan som denna, bliva räddad --
skulle vi väl nu på nytt bryta mot dina bud och befrynda oss med folk som bedriva sådana styggelser?
Skulle du då icke vredgas på oss, ända därhän att du förgjorde oss, så att intet mer vore kvar och ingen räddning funnes?
HERRE, Israels Gud, du är rättfärdig, ty av oss har allenast blivit kvar en räddad skara, såsom i dag nogsamt synes.
Och se, nu ligga vi här i vår skuld inför dig, ty vid sådant kan ingen bestå inför dig.»
Då nu Esra så bad och bekände, där han låg gråtande framför Guds hus, församlade sig till honom av Israel en mycket stor skara, män, kvinnor och barn; ty också folket grät bitterligen.
Och Sekanja, Jehiels son, av Ulams barn, tog till orda och sade till Esra: »Ja, vi hava varit otrogna mot vår Gud, i det att vi hava tagit till oss främmande kvinnor från de andra folken här i landet.
Dock finnes ännu hopp för Israel.
Så låt oss nu sluta ett förbund med vår Gud, att vi, i kraft av Herrens rådslut och de mäns som frukta för vår Guds bud, vilja avlägsna ifrån oss alla sådana kvinnor jämte deras barn; så bör ju ske efter lagen.
Stå upp, ty dig åligger denna sak, och vi vilja vara med dig.
Var frimodig och grip verket an.»
Då stod Esra upp och tog en ed av de översta bland prästerna, leviterna och hela Israel, att de skulle göra såsom det var sagt; och de gingo eden.
Och Esra stod upp från platsen framför Guds hus och gick in i Johanans, Eljasibs sons, tempelkammare.
Och när han hade kommit dit, kunde han varken äta eller dricka; så sörjde han över den otrohet som de återkomna fångarna hade begått.
Och man lät utropa i Juda och Jerusalem, bland alla dem som hade återkommit ifrån fångenskapen, att de skulle församla sig i Jerusalem;
och vilken som icke komme till den tredje dagen därefter, i enlighet med furstarnas och de äldstes beslut, hans hela egendom skulle givas till spillo, och han själv skulle avskiljas från de återkomna fångarnas församling.
Så församlade sig då alla Judas och Benjamins män i Jerusalem till den tredje dagen, det är på tjugonde dagen i nionde månaden; och allt folket stannade på den öppna platsen vid Guds hus, skälvande både på grund av den sak som förelåg och på grund av det starka regnet.
Och prästen Esra stod upp och sade till dem: »I haven varit otrogna, i det att I haven tagit till eder främmande kvinnor och därigenom ökat Israels skuld.
Men bekännen det nu, HERREN, edra fäders Gud, till pris, och gören hans vilja: skiljen eder från de andra folken här i landet och från de främmande kvinnorna.»
Då svarade hela församlingen och sade med hög röst: »Såsom du har sagt, så tillkommer det oss att göra.
Men folket är talrikt, och regntiden är nu inne, och man kan icke stå härute; detta ärende kan ej heller avslutas på en dag eller två, ty vi hava mycket förbrutit oss härutinnan.
Må därför våra furstar stå redo för hela församlingen, och må alla i våra städer, som hava tagit till sig främmande kvinnor, infinna sig på bestämda tider, och med dem de äldste i var stad och domarna där, till dess att vi hava avvänt ifrån oss vår Guds vredes glöd i denna sak.»
Allenast Jonatan, Asaels son, och Jaseja, Tikvas son, trädde upp häremot, och Mesullam jämte leviten Sabbetai understödde dem.
Men de som hade återkommit ifrån fångenskapen gjorde såsom det var sagt.
Och man utsåg prästen Esra och några av huvudmännen för familjerna, efter de särskilda familjerna, alla namngivna; och på första dagen i tionde månaden satte de sig att rannsaka härom.
Och till första dagen i första månaden hade de avslutat rannsakningen om allt som angick de män vilka hade tagit till sig främmande kvinnor.
Bland prästernas söner befunnos följande hava tagit till sig främmande kvinnor: Av Jesuas, Josadaks sons, barn och hans bröder: Maaseja, Elieser, Jarib och Gedalja,
vilka nu gåvo sin hand därpå att de skulle avlägsna ifrån sig sina kvinnor; och de skulle frambära en vädur såsom skuldoffer för den skuld de hade ådragit sig;
av Immers barn: Hanani och Sebadja;
av Harims barn: Maaseja, Elia, Semaja, Jehiel och Ussia;
av Pashurs barn: Eljoenai, Maaseja, Ismael, Netanel, Josabad och Eleasa.
Av leviterna: Josabad, Simei och Kelaja, som ock hette Kelita, Petaja, Juda och Elieser;
av sångarna: Eljasib; av dörrvaktarna: Sallum, Telem och Uri.
Av det övriga Israel: av Pareos' barn: Ramja, Issia, Malkia Mijamin, Eleasar, Malkia och Benaja;
av Elams barn: Mattanja, Sakarja, Jehiel, Abdi, Jeremot och Elia;
av Sattus barn: Eljoenai, Eljasib, Mattanja, Jeremot, Sabad och Asisa;
av Bebais barn: Johanan, Hananja, Sabbai, Atlai;
av Banis barn: Mesullam, Malluk, Adaja, Jasub, Seal och Jeremot;
av Pahat-Moabs barn: Adna och Kelal, Benaja, Maaseja, Mattanja, Besalel, Binnui och Manasse;
vidare Harims barn: Elieser, Issia, Malkia, Semaja, Simeon,
Benjamin, Malluk, Semarja;
av Hasums barn: Mattenai, Mattatta, Sabad, Elifelet, Jeremai, Manasse, Simei;
av Banis barn: Maadai, Amram och Uel,
Benaja, Bedeja, Keluhi,
Vanja, Meremot, Eljasib,
Mattanja, Mattenai och Jaasu,
vidare Bani, Binnui, Simei,
vidare Selemja, Natan och Adaja,
Maknaddebai, Sasai, Sarai,
Asarel, Selemja, Semarja,
Sallum, Amarja, Josef;
av Nebos barn: Jegiel, Mattitja, Sabad, Sebina, Jaddu, Joel och Benaja.
Alla dessa hade tagit främmande kvinnor till hustrur; och bland dessa funnos kvinnor som hade fött barn.
Nehemjas, Hakaljas sons, berättelse.
I månaden Kisleu, i det tjugonde året, när jag var i Susans borg,
hände sig att Hanani, en av mina bröder, och några andra män kommo från Juda.
Och jag frågade dem om judarna, den räddade skara som fanns kvar efter fångenskapen, och om Jerusalem.
De sade till mig: »De kvarblivna, de som efter fångenskapen finnas kvar i hövdingdömet, lida stor nöd och smälek, och Jerusalems mur är nedbruten, och dess portar äro uppbrända i eld.»
När jag hade hört detta, satt jag gråtande och sörjande i flera dagar och fastade och bad inför himmelens Gud.
Och jag sade: »Ack HERRE, himmelens Gud, du store och fruktansvärde Gud, du som håller förbund och bevarar nåd mot dem som älska dig och hålla dina bud,
låt ditt öra akta härpå, och låt dina ögon vara öppna, och hör din tjänares bön, den som jag nu beder inför dig både dag och natt, för Israels barn, dina tjänare, i det att jag bekänner Israels barns synder, dem som vi hava begått mot dig; ty också jag och min faders hus hava syndat.
Vi hava svårt förbrutit oss mot dig; vi hava icke hållit de bud och stadgar och rätter som du gav din tjänare Mose.
Men tänk på det ord som du gav din tjänare Mose, när du sade: 'Om I ären otrogna, så skall jag förströ eder bland folken;
men om I vänden om till mig och hållen mina bud och gören efter dem, då vill jag, om än edra fördrivna vore vid himmelens ända, likväl församla dem därifrån och låta dem komma till den plats som jag har utvalt till boning åt mitt namn.'
De äro ju dina tjänare och ditt folk, som du har förlossat genom din stora kraft och din starka hand.
Ack Herre, låt ditt öra akta på din tjänares bön, ja, på vad dina tjänare bedja, de som vilja frukta ditt namn; låt nu din tjänare vara lyckosam och låt honom finna barmhärtighet inför denne man.»
Jag var då munskänk hos konungen.
I månaden Nisan, i Artasastas tjugonde regeringsår, vid ett tillfälle då vin stod framsatt för konungen, tog jag vinet och gav det åt honom.
Och jag hade icke förr visat mig sorgsen inför honom;
men nu sade konungen till mig: »Varför ser du så sorgsen ut?
Du är ju icke sjuk; du måste hava någon hjärtesorg.»
Då blev jag övermåttan häpen.
Och jag sade till konungen: »Må konungen leva evinnerligen!
Skulle jag icke se sorgsen ut, då den stad där mina fäders gravar äro ligger öde och dess portar äro förtärda av eld?»
Konungen sade till mig: »Vad är det då du begär?»
Då bad jag en bön till himmelens Gud
och sade till konungen: »Om det så täckes konungen, och om du finner behag i din tjänare, så beder jag att du ville låta mig fara till Juda, till den stad där mina fäders gravar äro, på det att jag åter må bygga upp den.»
Då frågade konungen mig, allt under det att drottningen satt vid hans sida: »Huru länge kan din resa räcka, och när kan du komma tillbaka?»
Då det nu alltså täcktes konungen att låta mig fara, uppgav jag för honom en bestämd tid.
Och jag sade till konungen: »Om det så täckes konungen, så må brev givas mig till ståthållarna i landet på andra sidan floden, att de låta mig fara därigenom, till dess jag kommer till Juda,
så ock ett brev till Asaf, uppsyningsmannen över den kungliga skogsparken, att han låter mig få virke för att därmed timra upp portarna till borgen som hör till templet, ävensom virke till stadsmuren, så ock till det hus där jag själv skall hava min bostad.»
Och konungen beviljade mig detta, eftersom min Guds goda hand var över mig.
När jag så kom till ståthållarna i landet på andra sidan floden, gav jag dem konungens brev.
Och konungen hade sänt med mig härhövitsmän och ryttare.
Men då horoniten Sanballat och Tobia, den ammonitiske tjänstemannen, hörde detta, förtröt det dem högeligen att någon hade kommit för att se Israels barn till godo.
När jag sedan hade kommit till Jerusalem och varit där i tre dagar,
stod jag upp om natten jämte några få män, utan att hava omtalat för någon människa vad min Gud ingav mig i hjärtat att göra för Jerusalem; och det djur som jag red på var det enda jag hade med mig.
Och jag drog om natten ut genom Dalporten fram emot Drakkällan och Dyngporten och besåg Jerusalems murar, huru de voro nedbrutna, och huru dess portar voro förtärda av eld.
Och jag drog vidare till Källporten och till Konungsdammen, men där var det icke möjligt för djuret att komma fram med mig.
Då begav jag mig uppför dalen om natten och besåg muren och vände sedan åter in genom Dalporten och kom så tillbaka.
Och föreståndarna hade icke fått veta vart jag hade gått, och vad jag ville göra, ty jag hade ännu icke omtalat något för judarna, prästerna, ädlingarna, föreståndarna och de övriga, som skulle få med arbetet att göra.
Men nu sade jag till dem: »I sen själva i vilken nöd vi äro, huru Jerusalem ligger öde, och huru dess portar äro uppbrända i eld.
Välan då, låt oss bygga upp Jerusalems mur, för att vi icke längre må vara till smälek.»
Och jag omtalade för dem huru min Guds hand hade varit mig nådig, så ock vad konungen hade lovat mig.
Då sade de: »Vi vilja stå upp och bygga.»
Och de togo mod till sig för det goda verket.
Men när horoniten Sanballat och Tobia, den ammonitiske tjänstemannen, och araben Gesem hörde detta, bespottade de oss och visade förakt för oss; och de sade: »Vad är det I gören?
Viljen I sätta eder upp mot konungen?»
Då gav jag dem detta svar: »Himmelens Gud skall låta det gå oss väl, och vi, hans tjänare, vilja stå upp och bygga; men I haven ingen del eller rätt eller åminnelse i Jerusalem.»
Och översteprästen Eljasib och hans bröder, prästerna, stodo upp och byggde Fårporten, vilken de helgade, och i vilken de sedan satte in dörrarna.
Vidare byggde de ända fram till Hammeatornet, som de helgade, och vidare fram till Hananeltornet.
Därbredvid byggde Jerikos män; och därbredvid byggde Sackur, Imris son.
Fiskporten byggdes av Hassenaas barn; de timrade upp den och satte in dess dörrar, dess riglar och bommar.
Därbredvid arbetade Meremot, son till Uria, son till Hackos, på att sätta muren i stånd; därbredvid arbetade Mesullam, son till Berekja, son till Mesesabel; och därbredvid arbetade Sadok, Baanas son.
Därbredvid arbetade tekoaiterna, men de förnämsta bland dem ville icke böja sin hals till att tjäna sin Herre.
Gamla porten sattes i stånd av Jojada, Paseas son, och Mesullam, Besodjas son; de timrade upp den och satte in dess dörrar, dess riglar och bommar.
Därbredvid arbetade gibeoniten Melatja och meronotiten Jadon jämte männen från Gibeon och Mispa, som lydde under ståthållaren i landet på andra sidan floden.
Därbredvid arbetade Ussiel, Harhajas son, jämte guldsmederna; och därbredvid arbetade Hananja, en av salvoberedarna.
Det nästföljande stycket av Jerusalem lät man vara, ända till Breda muren.
Därbredvid arbetade Refaja, Hurs son, hövdingen över ena hälften av Jerusalems område.
Därbredvid arbetade Jedaja, Harumafs son, mitt emot sitt eget hus; och därbredvid arbetade Hattus, Hasabnejas son.
En annan sträcka sattes i stånd av Malkia, Harims son, och av Hassub, Pahat-Moabs son, och därjämte Ugnstornet.
Därbredvid arbetade Sallum, Hallohes' son, hövdingen över andra hälften av Jerusalems område, han själv med sina döttrar.
Dalporten sattes i stånd av Hanun och Sanoas invånare; de byggde upp den och satte in dess dörrar, dess riglar och bommar.
De byggde ock ett tusen alnar på muren, ända fram till Dyngporten.
Och Dyngporten sattes i stånd av Malkia, Rekabs son, hövdingen över Bet-Hackerems område; han byggde upp den och satte in dess dörrar, dess riglar och bommar.
Och Källporten sattes i stånd av Sallun, Kol-Hoses son, hövdingen över Mispas område; han byggde upp den och lade tak därpå och satte in dess dörrar, dess riglar och bommar.
Han byggde ock muren vid Vattenledningsdammen, invid den kungliga trädgården, ända fram till trapporna som föra ned från Davids stad.
Därnäst sattes ett stycke i stånd av Nehemja, Asbuks son, hövdingen över ena hälften av Bet-Surs område, nämligen stycket ända fram till platsen mitt emot Davidsgravarna och vidare fram till den grävda dammen och till Hjältehuset.
Därnäst arbetade leviterna under Rehum, Banis son; därbredvid arbetade Hasabja, hövdingen över ena hälften av Kegilas område, för sitt område.
Därnäst arbetade deras bröder under Bavai, Henadads son, hövdingen över andra hälften av Kegilas område.
Därbredvid sattes en annan sträcka i stånd av Eser, Jesuas son, hövdingen över Mispa, nämligen från platsen mitt emot uppgången till tyghuset i Vinkeln.
Därnäst sattes, under ivrigt arbete, en annan sträcka i stånd av Baruk, Sabbais son, från Vinkeln ända fram till ingången till översteprästen Eljasibs hus.
Därnäst sattes en annan sträcka i stånd av Meremot, son till Uria, son till Hackos, från ingången till Eljasibs hus ända dit där Eljasibs hus slutar.
Därnäst arbetade prästerna, männen från Jordanslätten.
Därnäst arbetade Benjamin och Hassub, mitt emot sitt eget hus; därnäst arbetade Asarja, son till Maaseja, son till Ananja, utmed sitt eget hus.
Därnäst sattes en annan sträcka i stånd av Binnui, Henadads son, från Asarjas hus ända fram till Vinkeln och vidare fram till Hörnet.
Palal, Usais son, satte i stånd stycket från platsen mitt emot Vinkeln och det torn som skjuter ut från det övre konungshuset, vid fängelsegården; därnäst kom Pedaja, Pareos' son.
(Men tempelträlarna bodde på Ofel ända fram till platsen mitt emot Vattenporten mot öster och det utskjutande tornet.)
Därnäst sattes en annan sträcka i stånd av tekoaiterna, från platsen mitt emot det stora utskjutande tornet ända fram till Ofelmuren.
Ovanför Hästporten arbetade prästerna, var och en mitt emot sitt eget hus.
Därnäst arbetade Sadok, Immers son, mitt emot sitt eget hus; och därnäst arbetade Semaja, Sekanjas son, som hade vakten vid Östra porten.
Därnäst sattes en annan sträcka i stånd av Hananja, Selemjas son, och Hanun, Salafs sjätte son; därnäst arbetade Mesullam, Berekjas son, mitt emot sin tempelkammare.
Därnäst sattes ett stycke i stånd av Malkia, en av guldsmederna, ända fram till tempelträlarnas och köpmännens hus, mitt emot Mönstringsporten och vidare fram till Hörnsalen.
Och mellan Hörnsalen och Fårporten arbetade guldsmederna och köpmännen på att sätta muren i stånd.
När nu Sanballat hörde att vi höllo på att bygga upp muren, vredgades han och blev högeligen förtörnad.
Och han bespottade judarna
och talade så inför sina bröder och inför Samariens krigsfolk: »Vad är det dessa vanmäktiga judar göra?
Skall man låta dem hållas?
Skola de få offra?
Skola de kanhända i sinom tid fullborda sitt verk?
Skola de kunna giva liv åt stenarna i grushögarna, där de ligga förbrända?»
Och ammoniten Tobia, som stod bredvid honom sade: »Huru de än bygga, skall dock en räv komma deras stenmur att rämna, blott han hoppar upp på den.»
Hör, vår Gud, huru föraktade vi äro.
Låt deras smädelser falla tillbaka på deras egna huvuden.
Ja, låt dem bliva utplundrade i ett land dit de föras såsom fångar.
Överskyl icke deras missgärningar, och låt deras synd icke varda utplånad ur din åsyn, eftersom de hava varit de byggande till förargelse.
Och vi byggde på muren, och hela muren blev hopfogad till sin halva höjd; och folket arbetade med gott mod.
Men när Sanballat och Tobia och araberna, ammoniterna och asdoditerna hörde att man alltjämt höll på med att laga upp Jerusalems murar, och att rämnorna begynte igentäppas, då blevo de mycket vreda.
Och de sammansvuro sig allasammans att gå åstad och angripa Jerusalem och störa folket i deras arbete.
Då bådo vi till vår Gud; och vi läto hålla vakt mot dem både dag och natt för att skydda oss mot dem.
Men judarna sade: »Bärarnas kraft sviker, och gruset är alltför mycket; vi förmå icke mer att bygga på muren.»
Våra ovänner åter sade: »Innan de få veta eller se något, skola vi stå mitt ibland dem och dräpa dem; så skola vi göra slut på arbetet.»
När nu de judar som bodde i deras grannskap kommo och från alla håll uppmanade oss, väl tio gånger, att vi skulle draga oss tillbaka till dem,
då ställde jag upp folket i de lägsta och mest öppna delarna av staden bakom muren; jag ställde upp dem efter släkter, med sina svärd, spjut och bågar.
Och sedan jag hade besett allt, stod jag upp och sade till ädlingarna och föreståndarna och det övriga folket: »Frukten icke för dem; tänken på Herren, den store och fruktansvärde, och striden för edra bröder, edra söner och döttrar, edra hustrur och edra hus.»
Sedan våra fiender sålunda hade fått förnimma att saken var oss bekant, och att Gud hade gjort deras råd om intet, kunde vi alla vända tillbaka till muren, var och en till sitt arbete.
Från den dagen var ena hälften av mina tjänare sysselsatt med arbetet, under det att andra hälften stod väpnad med sina spjut, sköldar, bågar och pansar, medan furstarna stodo bakom hela Juda hus.
De som byggde på muren och de som lassade på och buro bördor gjorde sitt arbete med den ena handen, och med den andra höllo de vapnet.
Och de som byggde hade var och en sitt svärd bundet vid sin länd, under det att de byggde; och bredvid mig stod en basunblåsare.
Jag hade nämligen sagt till ädlingarna och föreståndarna och det övriga folket: »Arbetet är stort och vidsträckt, och vi äro spridda över muren, långt ifrån varandra.
Där I nu hören basunen ljuda, dit skolen I församla eder till oss; vår Gud skall strida för oss.»
Så gjorde ock vi vårt arbete, under det att hälften av folket stod väpnad med sina spjut från morgonrodnadens uppgång, till dess att stjärnorna kommo fram.
Vid samma tid sade jag ock till folket att var och en med sin tjänare skulle stanna över natten inne i Jerusalem, så att vi om natten kunna hava dem till vakt och om dagen till arbete.
Och varken jag eller mina bröder eller mina tjänare eller de som gjorde vakt hos mig lade av kläderna; vapnen höllos av var och en för lika nödvändiga som vatten.
Och männen av folket med sina hustrur hovo upp ett stort rop mot sina judiska bröder.
Några sade: »Vi med våra söner och döttrar äro många; låt oss få säd, så att vi hava att äta och kunna bliva vid liv.»
Och några sade: »Våra åkrar, vingårdar och hus måste vi pantsätta; låt oss få säd till att stilla vår hunger.»
Och andra sade: »Vi hava måst låna penningar på våra åkrar och vingårdar till skatten åt konungen.
Nu äro ju våra kroppar lika goda som våra bröders kroppar, och våra barn lika goda som deras barn; men ändå måste vi giva våra söner och döttrar i träldom, ja, några av våra döttrar hava redan blivit givna i träldom, utan att vi förmå göra något därvid, eftersom våra åkrar och vingårdar äro i andras händer.»
När jag nu hörde deras rop och hörde dessa ord, blev jag mycket vred.
Och sedan jag hade gått till råds med mig själv, förebrådde jag ädlingarna och föreståndarna och sade till dem: »Det är ocker I bedriven mot varandra.»
Därefter sammankallade jag en stor folkförsamling emot dem.
Och jag sade till dem: »Vi hava efter förmåga friköpt våra judiska bröder som voro sålda åt hedningarna.
Skolen nu I sälja edra bröder?
Skola de behöva sälja sig åt oss?»
Då tego de och hade intet att svara.
Och jag sade: »Vad I gören är icke rätt.
I borden ju vandra i vår Guds fruktan, så att våra fiender, hedningarna, ej finge orsak att smäda oss.
Också jag och mina bröder och mina tjänare hava penningar och säd att fordra av dem; låt oss nu avstå från vår fordran.
Given dem redan i dag tillbaka deras åkrar, vingårdar, olivplanteringar och hus, och skänken efter den ränta på penningarna, på säden, på vinet och oljan, som I haven att fordra av dem.»
De svarade: »Vi vilja giva det tillbaka och icke utkräva något av dem; vi vilja göra såsom du har sagt.»
Och jag tog en ed av dem, sedan jag hade tillkallat prästerna, att de skulle göra så.
Därjämte skakade jag fånget på min mantel och sade: »Var och en som icke håller detta sitt ord, honom må Gud så skaka bort ifrån hans hus och hans gods; ja, varde han så utskakad och tom på allt.»
Och hela församlingen sade: »Amen», och lovade HERREN.
Därefter gjorde folket såsom det var sagt.
Ytterligare är att nämna att från den dag då jag förordnades att vara ståthållare över dem i Juda land, alltså från Artasastas tjugonde regeringsår ända till hans trettioandra, tolv hela år, varken jag eller mina bröder åto av ståthållarkosten.
De förra ståthållarna, de som hade varit före mig, hade betungat folket och tagit av dem mat och vin till ett värde av mer än fyrtio siklar silver, och jämväl deras tjänare hade förfarit hårt mot folket.
Men så gjorde icke jag, ty jag fruktade Gud.
Dessutom höll jag i att arbeta på muren, och ingen åker köpte vi oss; och alla mina tjänare voro församlade vid arbetet där.
Och av judarna och deras föreståndare åto ett hundra femtio man vid mitt bord, förutom dem som kommo till oss ifrån folken runt omkring oss.
Och vad som tillreddes för var dag, nämligen en oxe och sex utsökta får, förutom fåglar, det tillreddes på min bekostnad; och var tionde dag anskaffades mycket vin av alla slag.
Men likväl krävde jag icke ut ståthållarkosten, eftersom arbetet tyngde så svårt på folket.
Tänk, min Gud, på allt vad jag har gjort för detta folk, och räkna mig det till godo!
När nu Sanballat och Tobia och araben Gesem och våra övriga fiender hörde att jag hade byggt upp muren, och att det icke mer fanns någon rämna i den -- om jag ock vid den tiden ännu icke hade satt in dörrar i portarna --
då sände Sanballat och Gesem bud till mig och läto säga: »Kom, låt oss träda tillsammans i Kefirim i Onos dal.»
De tänkte nämligen göra mig något ont.
Men jag skickade bud till dem och lät säga: »Jag har ett stort arbete för händer och kan icke komma ned.
Arbetet kan ju icke vila, såsom dock måste ske, om jag lämnade det och komme ned till eder.»
Och de sände samma bud till mig fyra gånger; men var gång gav jag dem samma svar som förut.
Då sände Sanballat för femte gången till mig sin tjänare med samma bud, och denne hade nu med sig ett öppet brev.
Däri var skrivet: »Det förljudes bland folken, och påstås jämväl av Gasmu, att du och judarna haven i sinnet att avfalla, och att det är därför du bygger upp muren, ja, att du vill bliva deras konung -- sådant säger man.
Du lär ock hava beställt profeter som i Jerusalem skola utropa och förkunna att du är konung i Juda.
Eftersom nu konungen nog får höra talas härom, därför må du nu komma, så att vi få rådslå med varandra.»
Då sände jag bud till honom och lät svara: »Intet av det du säger har någon grund, utan det är dina egna påfund.»
De ville nämligen alla skrämma oss, i tanke att vi då skulle förlora allt mod till arbetet, och att detta så skulle bliva ogjort.
Styrk du nu i stället mitt mod!
Men jag gick hem till Semaja, son till Delaja, son till Mehetabel; han höll sig då inne.
Och han sade: »Låt oss tillsammans gå till Guds hus, in i templet, och sedan stänga igen templets dörrar.
Ty de skola komma för att dräpa dig; om natten skola de komma för att dräpa dig.»
Men jag svarade: »Skulle en man sådan som jag vilja fly?
Eller kan väl en man av mitt slag gå in i templet och dock bliva vid liv?
Nej, jag vill icke gå dit.»
Jag förstod nämligen att Gud icke hade sänt honom, utan att han förebådade mig sådant, blott därför att Tobia och Sanballat hade lejt honom.
Han var lejd, för att jag skulle låta skrämma mig till att göra såsom han sade och därmed försynda mig; på detta sätt ville de framkalla ont rykte om mig, för att sedan kunna smäda mig.
Tänk, min Gud på Tobia, ävensom Sanballat, efter dessa hans gärningar, så ock på profetissan Noadja och de andra profeterna som ville skrämma mig!
Och muren blev färdig på tjugufemte dagen i månaden Elul, efter femtiotvå dagar.
När nu alla våra fiender hörde detta, betogos de, alla de kringboende folken, av fruktan, och sågo att de hade kommit illa till korta; ty de förstodo nu att detta arbete var vår Guds verk.
Vid denna tid sände ock Juda ädlingar många brev till Tobia, och brev från Tobia ankommo ock till dem.
Ty många i Juda voro genom ed förbundna med honom; han var nämligen måg till Sekanja, Aras son, och hans son Johanan hade tagit till hustru en dotter till Mesullam, Berekjas son.
Dessa plägade också inför mig tala gott om honom, och vad jag sade buro de fram till honom.
Tobia sände ock brev för att skrämma mig.
När nu muren var uppbyggd, satte jag in dörrarna; och dörrvaktare, sångare och leviter blevo anställda.
Och till befälhavare över Jerusalem satte jag min broder Hanani jämte Hananja, hövitsman i borgen, ty denne hölls för en pålitlig man och var gudfruktig mer än många andra.
Och jag sade till dem: »Jerusalems portar må icke öppnas, förrän solen är högt uppe; och medan vakten ännu står kvar, skall man stänga dörrarna och sätta bommarna för.
Och I skolen ställa ut vakter av Jerusalems invånare, var och en på hans post, så att envar får stå framför sitt eget hus.»
Och staden var vidsträckt och stor, men där fanns icke mycket folk, och husen voro icke uppbyggda.
Och min Gud ingav mig i hjärtat att jag skulle församla ädlingarna, föreståndarna och folket för att upptecknas i släktregister.
Då fann jag släktförteckningen över dem som först hade dragit upp, och jag fann däri så skrivet:
»Dessa voro de män från hövdingdömet, som drogo upp ur den landsflykt och fångenskap till vilken de hade blivit bortförda av Nebukadnessar, konungen i Babel, och som vände tillbaka till Jerusalem och till Juda, var och en till sin stad,
i det att de följde med Serubbabel, Jesua, Nehemja, Asarja, Raamja, Nahamani, Mordokai, Bilsan, Misperet, Bigvai, Nehum och Baana.
Detta var antalet män av Israels meniga folk:
Pareos' barn: två tusen ett hundra sjuttiotvå;
Sefatjas barn: tre hundra sjuttiotvå;
Aras barn: sex hundra femtiotvå;
Pahat-Moabs barn, av Jesuas och Joabs barn: två tusen åtta hundra aderton;
Elams barn: ett tusen två hundra femtiofyra;
Sattus barn: åtta hundra fyrtiofem;
Sackais barn: sju hundra sextio;
Binnuis barn: sex hundra fyrtioåtta;
Bebais barn: sex hundra tjuguåtta;
Asgads barn: två tusen tre hundra tjugutvå;
Adonikams barn: sex hundra sextiosju;
Bigvais barn: två tusen sextiosju;
Adins barn: sex hundra femtiofem;
Aters barn av Hiskia: nittioåtta;
Hasums barn: tre hundra tjuguåtta;
Besais barn: tre hundra tjugufyra;
Harifs barn: ett hundra tolv;
Gibeons barn: nittiofem;
männen från Bet-Lehem och Netofa: ett hundra åttioåtta;
männen från Anatot: ett hundra tjuguåtta;
männen från Bet-Asmavet: fyrtiotvå;
männen från Kirjat-Jearim, Kefira och Beerot: sju hundra fyrtiotre;
männen från Rama och Geba: sex hundra tjuguen;
männen från Mikmas: ett hundra tjugutvå;
männen från Betel och Ai: ett hundra tjugutre;
männen från det andra Nebo: femtiotvå;
den andre Elams barn: ett tusen två hundra femtiofyra;
Harims barn: tre hundra tjugu;
Jerikos barn: tre hundra fyrtiofem;
Lods, Hadids och Onos barn: sju hundra tjuguen;
Senaas barn: tre tusen nio hundra trettio.
Av prästerna: Jedajas barn av Jesuas hus: nio hundra sjuttiotre;
Immers barn: ett tusen femtiotvå;
Pashurs barn: ett tusen två hundra fyrtiosju;
Harims barn: ett tusen sjutton.
Av leviterna: Jesuas barn av Kadmiel, av Hodevas barn: sjuttiofyra;
av sångarna: Asafs barn: ett hundra fyrtioåtta;
av dörrvaktarna: Sallums barn, Aters barn, Talmons barn, Ackubs barn, Hatitas barn, Sobais barn: ett hundra trettioåtta.
Av tempelträlarna: Sihas barn, Hasufas barn, Tabbaots barn,
Keros' barn, Sias barn, Padons barn,
Lebanas barn, Hagabas barn, Salmais barn,
Hanans barn, Giddels barn, Gahars barn,
Reajas barn, Resins barn, Nekodas barn,
Gassams barn, Ussas barn, Paseas barn,
Besais barn, Meunims barn, Nefusesims barn,
Bakbuks barn, Hakufas barn, Harhurs barn,
Basluts barn, Mehidas barn, Harsas barn,
Barkos' barn, Siseras barn, Temas barn,
Nesias barn, Hatifas barn.
Av Salomos tjänares barn: Sotais barn, Soferets barn, Peridas barn,
Jaalas barn, Darkons barn, Giddels barn,
Sefatjas barn, Hattils barn, Pokeret-Hassebaims barn, Amons barn.
Tempelträlarna och Salomos tjänares barn utgjorde tillsammans tre hundra nittiotvå.
Och dessa voro de som drogo åstad från Tel-Mela, Tel-Harsa, Kerub, Addon och Immer, men som icke kunde uppgiva sina familjer och sin släkt, och huruvida de voro av Israel:
Delajas barn, Tobias barn, Nekodas barn, sex hundra fyrtiotvå.
Och av prästerna: Habajas barn, Hackos' barn, Barsillais barn, hans som tog en av gileaditen Barsillais döttrar till hustru och blev uppkallad efter deras namn.
Dessa sökte efter sina släktregister, men man kunde icke finna dem; därför blevo de såsom ovärdiga uteslutna från prästadömet.
Och ståthållaren tillsade dem att de icke skulle få äta av det högheliga, förrän en präst uppstode med urim och tummim.
Hela församlingen utgjorde sammanräknad fyrtiotvå tusen tre hundra sextio,
förutom deras tjänare och tjänarinnor, som voro sju tusen tre hundra trettiosju.
Och till dem hörde två hundra fyrtiofem sångare och sångerskor.
124920
Och de hade fyra hundra trettiofem kameler och sex tusen sju hundra tjugu åsnor.
Och somliga bland huvudmännen för familjerna gåvo skänker till arbetet.
Ståthållaren gav till kassan i guld ett tusen dariker, därtill femtio skålar och fem hundra trettio prästerliga livklädnader.
Och somliga bland huvudmännen för familjerna gåvo till arbetskassan i guld tjugu tusen dariker och i silver två tusen två hundra minor.
Och det övriga folkets gåvor utgjorde i guld tjugu tusen dariker och i silver två tusen minor, så ock sextiosju prästerliga livklädnader.
Och prästerna, leviterna, dörrvaktarna, sångarna, en del av meniga folket samt tempelträlarna, korteligen hela Israel, bosatte sig i sina städer.»
När sjunde månaden nalkades och Israels barn voro bosatta i sina städer, församlade sig folket, alla såsom en man, på den öppna platsen framför Vattenporten; och de bådo Esra, den skriftlärde, att hämta fram Moses lagbok, den som HERREN hade givit åt Israel.
Då framlade prästen Esra lagen för församlingen, för både män och kvinnor, alla som kunde förstå vad de hörde; detta var på första dagen i sjunde månaden.
Och han föreläste därur vid den öppna platsen framför Vattenporten, från dagningen till middagen, för män och kvinnor, dem som kunde förstå det; och allt folket lyssnade till lagboken.
Och Esra, den skriftlärde, stod på en hög träställning som man hade gjort för det ändamålet; och bredvid honom stodo Mattitja, Sema, Anaja, Uria, Hilkia och Maaseja på hans högra sida, och till vänster om honom Pedaja, Misael, Malkia, Hasum, Hasbaddana, Sakarja och Mesullam.
Och Esra öppnade boken, så att allt folket såg det, ty han stod högre än allt folket; och när han öppnade den, stod allt folket upp.
Och Esra lovade den store HERREN Gud, och allt folket svarade: »Amen, Amen», med uppräckta händer; och de böjde sig ned och tillbådo HERREN med ansiktet mot jorden.
Och Jesua, Bani, Serebja, Jamin, Ackub, Sabbetai, Hodia, Maaseja, Kelita, Asarja, Josabad, Hanan, Pelaja och de andra leviterna undervisade folket i lagen, medan folket stod där, var och en på sin plats.
Och de föreläste tydligt ur boken, ur Guds lag; och de utlade meningen, så att man förstod det som lästes.
Och Nehemja, han som var ståthållare, och prästen Esra, den skriftlärde, och leviterna, som undervisade folket, sade till allt folket: »Denna dag är helgad åt HERREN, eder Gud; sörjen icke och gråten icke.»
Ty allt folket grät, när de hörde lagens ord.
Och han sade ytterligare till dem: »Gån bort och äten eder bästa mat och dricken edert sötaste vin, och sänden omkring gåvor därav till dem som icke hava något tillrett åt sig, ty denna dag är helgad åt vår Herre.
Och varen icke bedrövade, ty fröjd i HERREN är eder starkhet.»
Också leviterna lugnade allt folket och sade: »Varen stilla, ty dagen är helig; varen icke bedrövade.»
Och allt folket gick bort och åt och drack; de sände ock omkring gåvor av den mat de hade tillagat och gjorde sig mycket glada; ty de hade aktat på det som man hade kungjort för dem.
Dagen därefter församlade sig huvudmännen för hela folkets familjer, så ock prästerna och leviterna, till Esra, den skriftlärde, för att giva närmare akt på lagens ord.
Och de funno skrivet i lagen att HERREN genom Mose hade bjudit att Israels barn skulle bo i lövhyddor under högtiden i sjunde månaden,
och att man skulle kungöra och låta utropa i alla deras städer och i Jerusalem och säga: »Gån ut på bergen och hämten löv av olivträd, planterade eller vilda, och löv av myrten, palmträd och andra lummiga träd, och gören lövhyddor, såsom det är föreskrivet.»
Då gick folket ut och hämtade sådant och gjorde sig hyddor på tak och på gårdar, var och en åt sig, så ock på gårdarna till Guds hus och på den öppna platsen vid Vattenporten och på den öppna platsen vid Efraimsporten.
Och hela församlingen, så många som hade kommit tillbaka ifrån fångenskapen, gjorde sig lövhyddor och bodde i dessa hyddor.
Ty från Jesuas, Nuns sons, dagar ända till den dagen hade Israels barn icke gjort så.
Och där rådde mycket stor glädje.
Och man föreläste ur Guds lagbok var dag, från den första dagen till den sista.
Och de höllo högtid i sju dagar, och på åttonde dagen hölls en högtidsförsamling på föreskrivet sätt.
Men på tjugufjärde dagen i samma månad församlade sig Israels barn och höllo fasta och klädde sig i sorgdräkt och strödde jord på sina huvuden.
Och de som voro av Israels släkt avskilde sig från alla främlingar och trädde så fram och bekände sina synder och sina fäders missgärningar.
Och de stodo upp, var och en på sin plats, och man föreläste ur HERRENS, deras Guds, lagbok under en fjärdedel av dagen; och under en annan fjärdedel bekände de sina synder och tillbådo HERREN, sin Gud.
Och Jesua och Bani, Kadmiel, Sebanja, Bunni, Serebja, Bani och Kenani trädde upp på leviternas upphöjning och ropade med hög röst till HERREN, sin Gud.
Och leviterna Jesua och Kadmiel, Bani, Hasabneja, Serebja, Hodia, Sebanja och Petaja sade: »Stån upp och loven HERREN, eder Gud, från evighet till evighet.
Ja, lovat vare ditt härliga namn, som är upphöjt över allt lov och pris.
Du allena är HERREN.
Du har gjort himlarna och himlarnas himmel och hela deras härskara, jorden och allt vad därpå är, haven och allt vad som är i dem, och det är du som behåller det allt vid liv; och himmelens härskara tillbeder dig.
Du är HERREN Gud, som utvalde Abram och förde honom ut från det kaldeiska Ur och gav honom namnet Abraham.
Och du fann hans hjärta fast i tron inför dig, och du slöt med honom det förbundet att du skulle giva åt hans säd kananéernas, hetiternas, amoréernas, perisséernas, jebuséernas och girgaséernas land, ja, giva det åt dem; och du uppfyllde dina ord, ty du är rättfärdig.
Och du såg till våra fäders betryck i Egypten och hörde deras rop vid Röda havet.
Du gjorde tecken och under på Farao och på alla hans tjänare och på allt folket i hans land; ty du förnam att dessa handlade övermodigt mot dem, och du gjorde dig ett namn, som är detsamma än i dag.
Havet klöv du itu för dem, så att de gingo mitt igenom havet på torr mark; men deras förföljare lät du sjunka i djupet såsom stenar, i väldiga vatten.
Du ledde dem om dagen med en molnstod, och om natten med en eldstod, för att lysa dem på den väg de skulle gå.
Och du steg ned på berget Sinai och talade till dem från himmelen och gav dem rättfärdiga rätter och riktiga lagar, goda stadgar och bud.
Du gav dem kunskap om din heliga sabbat och gav dem bud och stadgar och lag genom din tjänare Mose.
Och du gav dem bröd från himmelen, när de hungrade, och lät vatten komma ut ur klippan, när de törstade; och du tillsade dem att gå och taga i besittning det land som du med upplyft hand hade lovat giva åt dem.
Men våra fäder, de voro övermodiga; de voro hårdnackade, så att de icke hörde på dina bud.
De ville icke höra och tänkte icke på de under som du hade gjort med dem, utan voro hårdnackade och valde i sin gensträvighet en anförare, för att vända tillbaka till sin träldom.
Men du är en förlåtande Gud, nådig och barmhärtig, långmodig och stor i mildhet; och du övergav dem icke.
Nej, fastän de gjorde åt sig en gjuten kalv och sade: 'Detta är din Gud, han som har fört dig upp ur Egypten', och fastän de gjorde sig skyldiga till stora hädelser,
så övergav du dem likväl icke i öknen, efter din stora barmhärtighet.
Molnstoden vek om dagen icke ifrån dem, utan ledde dem på vägen, ej heller eldstoden om natten, utan lyste dem på den väg de skulle gå.
Din gode Ande sände du att undervisa dem, och ditt manna förvägrade du icke deras mun, och vatten gav du dem, när de törstade.
I fyrtio år försörjde du dem i öknen, så att intet fattades dem; deras kläder blevo icke utslitna, och deras fötter svullnade icke.
Och du gav dem riken och folk och utskiftade lotter åt dem på skilda håll; och de intogo Sihons land, det land som tillhörde konungen i Hesbon, och det land som tillhörde Og, konungen i Basan
Och du lät deras barn bliva talrika såsom stjärnorna på himmelen, och förde dem in i det land varom du hade sagt till deras fäder att de skulle komma dit och taga det i besittning.
Så kommo då barnen och togo landet i besittning, och du kuvade för dem landets inbyggare, kananéerna, och gav dessa i deras hand, både konungarna och folken där i landet, så att de gjorde med dem vad de ville.
Och de intogo befästa städer och ett bördigt land och kommo i besittning av hus, fulla med allt gott, och av uthuggna brunnar, vingårdar, olivplanteringar och fruktträd i myckenhet; och de åto och blevo mätta och feta och gjorde sig glada dagar av ditt myckna goda.
Men de blevo gensträviga och satte sig upp mot dig och kastade din lag bakom sin rygg och dräpte dina profeter, som varnade dem och ville omvända dem till dig; och de gjorde sig skyldiga till stora hädelser.
Då gav du dem i deras ovänners hand, så att dessa förtryckte dem; men när de i sin nöds tid ropade till dig, hörde du det från himmelen, och efter din stora barmhärtighet gav du dem frälsare, som frälste dem ur deras ovänners hand.
När de så kommo till ro, gjorde de åter vad ont var inför dig.
Då överlämnade du dem i deras fienders hand, så att dessa fingo råda över dem; men när de åter ropade till dig, då hörde du det från himmelen och räddade dem efter din barmhärtighet, många gånger.
Och du varnade dem och ville omvända dem till din lag; men de voro övermodiga och hörde icke på dina bud, utan syndade mot dina rätter, om vilka det gäller att den människa som gör efter dem får leva genom dem; de spjärnade emot i gensträvighet och voro hårdnackade och ville icke höra.
Du hade fördrag med dem i många år och varnade dem med din Ande genom dina profeter, men de lyssnade icke därtill; då gav du dem i de främmande folkens hand.
Men i din stora barmhärtighet gjorde du icke alldeles ände på dem och övergav dem icke; ty du är en nådig och barmhärtig Gud.
Och nu, vår Gud, du store, väldige och fruktansvärde Gud, du som håller förbund och bevarar nåd, nu må du icke akta för ringa all den vedermöda som har träffat oss, våra konungar, våra furstar, våra präster, våra fäder och hela ditt folk, ifrån de assyriska konungarnas dagar ända till denna dag.
Nej, du är rättfärdig vid allt det som har kommit över oss; ty du har visat dig trofast, men vi hava varit ogudaktiga.
Och våra konungar, våra furstar, våra präster och våra fäder hava icke gjort efter din lag och icke aktat på dina bud och på de varningar som du har låtit komma till dem.
Och fastän de sutto i sitt eget rike i det myckna goda som du hade givit dem, och i det rymliga och bördiga land som du hade upplåtit för dem, hava de ändå icke tjänat dig och icke omvänt sig från sina onda gärningar.
Se, vi äro nu andras tjänare; i det land som du gav åt våra fäder, för att de skulle äta dess frukt och dess goda, just där äro vi andras tjänare,
och sin rika avkastning giver det åt de konungar som du för våra synders skull har satt över oss.
Och de råda över våra kroppar och vår boskap såsom de vilja, och vi äro i stor nöd.»
På grund av allt detta slöto vi ett fast förbund och uppsatte det skriftligen; och på skrivelsen, som försågs med sigill, stodo våra furstars, våra leviters och våra prästers namn.
Följande namn stodo på skrivelserna som buro sigillen: Nehemja, ståthållaren, Hakaljas son, och Sidkia,
Seraja, Asarja, Jeremia,
Pashur, Amarja, Malkia,
Hattus, Sebanja, Malluk,
Harim, Meremot, Obadja,
Daniel, Ginneton, Baruk,
Mesullam, Abia, Mijamin,
Maasja, Bilgai, Semaja; dessa voro prästerna.
Och leviterna voro: Jesua, Asanjas son, Binnui, av Henadads barn, Kadmiel,
så ock deras bröder: Sebanja, Hodia, Kelita, Pelaja, Hanan,
Mika, Rehob, Hasabja,
Sackur, Serebja, Sebanja,
Hodia, Bani och Beninu.
Folkets huvudmän voro: Pareos, Pahat-Moab, Elam, Sattu, Bani,
Bunni, Asgad, Bebai,
Adonia, Bigvai, Adin,
Ater, Hiskia, Assur,
Hodia, Hasum, Besai,
Harif, Anatot, Nobai,
Magpias, Mesullam, Hesir,
Mesesabel, Sadok, Jaddua,
Pelatja, Hanan, Anaja,
Hosea, Hananja, Hassub,
Hallohes, Pilha, Sobek,
Rehum, Hasabna, Maaseja,
Ahia, Hanan, Anan,
Malluk, Harim och Baana.
Och det övriga folket, prästerna, leviterna, dörrvaktarna, sångarna, tempelträlarna och alla de som hade avskilt sig från de främmande folken och vänt sig till Guds lag, så ock deras hustrur, söner och döttrar, alla som hade kommit till moget förstånd,
dessa slöto sig till sina förnämligare bröder och gingo ed och svuro att de skulle vandra efter Guds lag, den som hade blivit given genom Guds tjänare Mose, och att de skulle hålla och göra efter alla HERRENS, vår HERRES, bud och rätter och stadgar,
att vi icke skulle giva våra döttrar åt de främmande folken, ej heller taga deras döttrar till hustrur åt våra söner.
Och när de främmande folken förde in handelsvaror eller något slags säd till salu på sabbatsdagen, skulle vi icke köpa det av dem på sabbat eller helgdag; och vi skulle låta vart sjunde år vara friår och då avstå från alla slags krav.
Och vi fastställde för oss den förpliktelsen att såsom vår gärd årligen erlägga en tredjedels sikel till tjänsten i vår Guds hus,
nämligen till skådebröden, och till det dagliga brännoffret, och till offren på sabbaterna, vid nymånaderna och högtiderna, och till tackoffren, och till syndoffren för Israels försoning, och till allt arbete i vår Guds hus.
Och vi, prästerna, leviterna och folket, kastade lott angående vedoffret, huru man årligen skulle föra det till vår Guds hus på bestämda tider, efter våra familjer, för att antändas på HERRENS, vår Guds, altare, såsom det är föreskrivet i lagen.
Och vi skulle årligen föra till HERRENS hus förstlingen av vår mark, och förstlingen av all frukt på alla slags träd,
och de förstfödda av våra söner och av vår boskap, såsom det är föreskrivet i lagen; vi skulle föra till vår Guds hus de förstfödda både av våra fäkreatur och av vår småboskap, till prästerna som gjorde tjänst i vår Guds hus.
Och förstlingen av vårt mjöl och våra offergärder, så ock av allt slags trädfrukt, av vin och olja skulle vi föra till prästerna, in i kamrarna i vår Guds hus, och tionden av vår jord till leviterna; ty det var leviterna som skulle uppbära tionden i alla de städer vid vilka vi brukade jorden.
Och en präst, en av Arons söner, skulle vara med leviterna, när leviterna uppburo tionden; och själva skulle leviterna föra tionden av sin tionde upp till vår Guds hus, in i förrådshusets kamrar.
Ty såväl de övriga israeliterna som Levi barn skulle föra sin offergärd av säd, vin och olja in i dessa kamrar, där helgedomens kärl och de tjänstgörande prästerna, ävensom dörrvaktarna och sångarna voro.
Alltså skulle vi icke försumma vår Guds hus.
Och folkets furstar bodde i Jerusalem; men det övriga folket kastade lott, för att så var tionde man skulle utses att bo i Jerusalem, den heliga staden, medan nio tiondedelar skulle bo i de andra städerna.
Och folket välsignade alla de män som frivilligt bosatte sig i Jerusalem.
Och de huvudmän i hövdingdömet, som bodde i Jerusalem, bodde var och en där han hade sin arvsbesittning, i sin stad; vanliga israeliter, präster, leviter och tempelträlar, så ock Salomos tjänares barn.
I Jerusalem bodde en del av Juda barn och en del av Benjamins barn, nämligen: Av Juda barn: Ataja, son till Ussia, son till Sakarja, son till Amarja, son till Sefatja, son till Mahalalel, av Peres' barn,
så ock Maaseja, son till Baruk, son till Kol-Hose, son till Hasaja, son till Adaja, son till Jojarib, son till Sakarja, silonitens son.
Peres' barn som bodde i Jerusalem utgjorde tillsammans fyra hundra sextioåtta stridbara män.
Och Benjamins barn voro dessa: Sallu, son till Mesullam, son till Joed, son till Pedaja, son till Kolaja, son till Maaseja, son till Itiel, son till Jesaja,
och näst honom Gabbai och Sallai, nio hundra tjuguåtta.
Joel, Sikris son, var tillsyningsman över dem, och Juda, Hassenuas son, var den andre i befälet över staden.
Av prästerna: Jedaja, Jojaribs son, Jakin
samt Seraja, son till Hilkia, son till Mesullam, son till Sadok, son till Merajot, son till Ahitub, fursten i Guds hus,
så ock deras bröder, som förrättade sysslorna i huset, åtta hundra tjugutvå; vidare Adaja, son till Jeroham, son till Pelalja, son till Amsi, son till Sakarja, son till Pashur, son till Malkia,
så ock hans bröder, huvudmän för familjer, två hundra fyrtiotvå; vidare Amassai, son till Asarel, son till Asai, son till Mesillemot, son till Immer,
så ock deras bröder, dugande män, ett hundra tjuguåtta; och tillsyningsman över dem var Sabdiel, Haggedolims son.
Och av leviterna: Semaja, son till Hassub, son till Asrikam, son till Hasabja, son till Bunni,
så ock Sabbetai och Josabad, som hade uppsikten över de yttre sysslorna vid Guds hus och hörde till leviternas huvudmän,
vidare Mattanja, son till Mika, son till Sabdi, son till Asaf, sånganföraren, som vid bönen tog upp lovsången, och Bakbukja, den av hans bröder, som var närmast efter honom, och Abda, son till Sammua, son till Galal, son till Jeditun.
Leviterna i den heliga staden utgjorde tillsammans två hundra åttiofyra.
Och dörrvaktarna, Ackub, Talmon och deras bröder, som höllo vakt vid portarna, voro ett hundra sjuttiotvå.
Och de övriga israeliterna, prästerna och leviterna bodde i alla de andra städerna i Juda, var och en i sin arvedel.
Men tempelträlarna bodde på Ofel, och Siha och Gispa hade uppsikten över tempelträlarna.
Och tillsyningsman bland leviterna i Jerusalem vid sysslorna i Guds hus var Ussi, son till Bani, son till Hasabja, son till Mattanja, son till Mika, av Asafs barn, sångarna.
Ty ett kungligt påbud var utfärdat angående dem, och en bestämd utanordning var för var dag fastställd för sångarna.
Och Petaja, Mesesabels son, av Seras, Judas sons, barn, gick konungen till handa i var sak som rörde folket.
Och i byarna med tillhörande utmarker bodde ock en del av Juda barn: i Kirjat-Arba och underlydande orter, I Dibon och underlydande orter, i Jekabseel och dess byar,
vidare i Jesua, Molada, Bet-Pelet
och Hasar-Sual, så ock i Beer-Seba och underlydande orter,
i Siklag, ävensom i Mekona och underlydande orter,
i En-Rimmon, Sorga, Jarmut,
Sanoa, Adullam och deras byar, i Lakis med dess utmarker, i Aseka och underlydande orter; och de hade sina boningsorter från Beer- Seba ända till Hinnoms dal.
Och Benjamins barn hade sina boningsorter från Geba: i Mikmas och Aja, så ock i Betel och underlydande orter,
i Anatot, Nob, Ananja,
Hasor, Rama, Gittaim,
Hadid, Seboim, Neballat,
Lod, Ono, och Timmermansdalen.
Och av leviterna blevo några avdelningar från Juda räknade till Benjamin.
Och dessa voro de präster och leviter som drogo upp med Serubbabel, Sealtiels son, och Jesua: Seraja, Jeremia, Esra,
Amarja, Malluk, Hattus,
Sekanja, Rehum, Meremot,
Iddo, Ginnetoi, Abia,
Mijamin, Maadja, Bilga,
Semaja, Jojarib, Jedaja,
Sallu, Amok, Hilkia och Jedaja.
Dessa voro huvudmän för prästerna och för sina bröder i Jesuas tid.
Och leviterna voro: Jesua, Binnui, Kadmiel, Serebja, Juda och Mattanja, som jämte sina bröder förestod lovsången;
vidare Bakbukja och Unno, deras bröder, som hade sina platser mitt emot dem, så att var avdelning hade sin tjänstgöring.
Och Jesua födde Jojakim, och Jojakim födde Eljasib, och Eljasib Jojada,
och Jojada födde Jonatan, och Jonatan födde Jaddua.
Och i Jojakims tid voro huvudmännen för prästernas familjer följande: för Seraja Meraja, för Jeremia Hananja,
för Esra Mesullam, för Amarja Johanan,
för Malluki Jonatan, för Sebanja Josef,
för Harim Adna, för Merajot Helkai,
för Iddo Sakarja, för Ginneton Mesullam,
för Abia Sikri, för Minjamin, för Moadja Piltai,
för Bilga Sammua, för Semaja Jonatan,
för Jojarib Mattenai, för Jedaja Ussi,
för Sallai Kallai, för Amok Eber,
för Hilkia Hasabja, för Jedaja Netanel.
I Eljasibs, Jojadas, Johanans och Jadduas tid blevo huvudmännen för leviternas familjer upptecknade, ävenså prästerna under persern Darejaves' regering.
Huvudmännen för Levi barns familjer äro upptecknade i krönikeboken, ända till Johanans, Eljasibs sons, tid.
Och leviternas huvudmän voro Hasabja, Serebja och Jesua, Kadmiels son, samt deras bröder, som stodo mitt emot dem för att lova och tacka, såsom gudsmannen David hade bjudit, den ena tjänstgörande avdelningen jämte den andra.
Mattanja, Bakbukja, Obadja, Mesullam, Talmon och Ackub höllo såsom dörrvaktare vakt över förrådshusen vid portarna.
Dessa levde i Jojakims, Jesuas sons, Josadaks sons, tid, och i Nehemjas, ståthållarens, och i prästen Esras, den skriftlärdes, tid.
Och när Jerusalems mur skulle invigas, uppsökte man leviterna på alla deras orter och förde dem till Jerusalem för att hålla invignings- och glädjehögtid under tacksägelse och sång, med cymbaler, psaltare och harpor.
Då församlade sig sångarnas barn såväl från nejden runt omkring Jerusalem som från netofatiternas byar,
ävensom från Bet-Haggilgal och från Gebas och Asmavets utmarker; ty sångarna hade byggt sig byar runt omkring Jerusalem.
Och prästerna och leviterna renade sig och renade sedan folket, portarna och muren.
Och jag lät Juda furstar stiga upp på muren.
Därefter anordnade jag två stora lovsångskörer och högtidståg; den ena kören gick till höger ovanpå muren, fram till Dyngporten.
Och dem följde Hosaja och ena hälften av Juda furstar
samt Asarja, Esra och Mesullam,
Juda, Benjamin, Semaja och Jeremia,
ävensom några av prästerna söner med trumpeter, vidare Sakarja, son till Jonatan, son till Semaja, son till Mattanja, son till Mikaja, son till Sackur, son till Asaf,
så ock hans bröder Semaja, Asarel, Milalai, Gilalai, Maai, Netanel och Juda samt Hanani, med gudsmannen Davids musikinstrumenter; och Esra, den skriftlärde, gick i spetsen för dem.
Och de gingo över Källporten och rakt fram uppför trapporna till Davids stad, på trappan i muren ovanför Davids hus, ända fram till Vattenporten mot öster.
Och efter den andra lovsångskören, som gick åt motsatt håll, följde jag med andra hälften av folket, ovanpå muren, upp genom Ugnstornet ända till Breda muren,
vidare över Efraimsporten, Gamla porten och Fiskporten och genom Hananeltornet, ända fram till Fårporten; och de stannade vid Fängelseporten.
Sedan trädde de båda lovsångskörerna upp i Guds hus, och likaså jag och ena hälften av föreståndarna jämte mig,
så ock prästerna Eljakim, Maaseja, Minjamin, Mikaja, Eljoenai, Sakarja och Hananja, med trumpeterna,
och Maaseja, Semaja, Eleasar, Ussi, Johanan, Malkia, Elam och Eser.
Och sångarna läto sången ljuda under Jisrajas anförarskap.
Och de offrade på den dagen stora offer och voro glada, ty Gud hade berett dem stor glädje; också kvinnor och barn voro glada.
Och glädjen från Jerusalem hördes vida omkring.
Vid samma tid tillsattes män som skulle förestå förrådskamrarna där offergärder, förstling och tionde nedlades; de skulle i dem hopsamla från stadsåkrarna det som efter lagen tillkom prästerna och leviterna.
Ty glädje rådde i Juda över att prästerna och leviterna nu gjorde sin tjänst.
Dessa iakttogo nu vad som var att iakttaga vid gudstjänsten och vid reningarna, och likaså gjorde sångarna och dörrvaktarna sin tjänst, såsom David och hans son Salomo hade bjudit.
Ty redan i fordom tid, på Davids och Asafs tid, hans som var anförare för sångarna, sjöngos lov- och tacksägelsesånger till Gud.
Och nu under Serubbabels och Nehemjas tid gav hela Israel åt sångarna och dörrvaktarna vad som tillkom dem för var dag; och man gav åt leviterna deras helgade andel, och leviterna gåvo åt Arons söner deras helgade andel.
Vid samma tid föreläste man ur Moses bok för folket, och man fann däri skrivet att ingen ammonit eller moabit någonsin skulle få komma in i Guds församling,
därför att de icke hade kommit Israels barn till mötes med mat och dryck, utan hade lejt Bileam emot dem till att förbanna dem; fastän vår Gud förvandlade förbannelsen till välsignelse.
Och när de hade hört lagen, avskilde de allt slags främmande folk från Israel.
Men en tid förut hade prästen Eljasib, som var satt att förestå kammaren i vår Guds hus, och som var en frände till Tobia,
åt denne inrett en stor kammare, där man förut plägade lägga in spisoffret, rökelsen och kärlen och den tionde av säd, vin och olja, som var bestämd åt leviterna, sångarna och dörrvaktarna, så ock offergärden åt prästerna.
Men under allt detta var jag icke i Jerusalem; ty i den babyloniske konungen Artasastas trettioandra regeringsår hade jag återkommit till konungen.
Men sedan jag efter någon tid hade utbett mig tillstånd av konungen,
begav jag mig till Jerusalem.
Och när jag där förnam det onda som Eljasib hade gjort till förmån för Tobia, då han hade inrett åt honom en kammare i förgårdarna till Guds hus,
misshagade detta mig högeligen; och jag lät kasta allt Tobias bohag ut ur kammaren.
Därefter tillsade jag att man skulle rena kamrarna, och jag lät åter ställa in i dem Guds hus' kärl, så ock spisoffret och rökelsen.
Och när jag vidare fick veta att man icke hade givit åt leviterna vad dem tillkom, varför ock leviterna och sångarna, i stället för att förrätta sina sysslor, hade avvikit var och en till sitt jordagods,
då förebrådde jag föreståndarna detta och sade: »Varför har Guds hus blivit så försummat?»
Och jag hämtade dem tillhopa och lät dem inställa sig på sina platser.
Och hela Juda förde fram till förrådshusen sin tionde av säd, vin och olja;
och jag satte prästen Selemja och Sadok, den skriftlärde, och Pedaja, en av leviterna, till förvaltare över förrådshusen och gav dem till biträde Hanan, son till Sackur, son till Mattanja; ty dessa voro ansedda såsom pålitliga män, och de skulle nu ombesörja utdelningen åt sina bröder.
Tänk fördenskull på mig, min Gud, och låt icke de fromma gärningar bliva utplånade, som jag har gjort för min Guds hus och för tjänstgöringen där!
Vid samma tid såg jag i Juda huru man trampade vinpressarna på sabbaten och förde hem säd, som man lastade på åsnor, så ock vin, druvor och fikon och annat lastgods av olika slag, och huru man förde sådant till Jerusalem på sabbatsdagen; och jag varnade dem, när de sålde dessa livsförnödenheter.
Och tyrierna, som vistades där, förde in fisk och alla slags varor och sålde dem på sabbaten till judarna, och detta i Jerusalem.
Då förebrådde jag Juda ädlingar detta och sade till dem: »Huru kunnen I handla så illa och därmed ohelga sabbatsdagen?
Var det icke därför att edra fäder gjorde sådant som vår Gud lät all denna olycka komma över oss och över denna stad?
Och nu dragen I ännu större vrede över Israel genom att så ohelga sabbaten.»
Och så snart det begynte bliva mörkt i Jerusalems portar före sabbaten, tillsade jag att man skulle stänga dörrarna; jag tillsade ock att man icke skulle öppna dem förrän efter sabbaten.
Och jag ställde några av mina tjänare på vakt vid portarna, för att intet lastgods skulle kunna föras in på sabbatsdagen.
Då stannade köpmän och försäljare av alla slags varor utanför Jerusalem över natten, och det både en och två gånger.
Men jag varnade dem och sade till dem: »Varför stannen I över natten framför muren?
Om I ännu en gång gören så, skall jag låta min hand drabba eder.»
Och jag tillsade leviterna att de skulle rena sig och komma och hålla vakt vid portarna, för att sabbatsdagen måtte hållas helig.
Tänk ock därför på mig, min Gud, och hav misskund med mig efter din stora nåd!
På den tiden såg jag också judiska män som hade tagit till sig asdoditiska, ammonitiska och moabitiska kvinnor.
Och deras barn talade till hälften asdoditiska -- ty judiska kunde de icke tala riktigt -- eller ock något av de andra folkens tungomål.
Då förebrådde jag dem detta och uttalade förbannelser över dem, ja, några av dem slog jag och ryckte jag i skägget.
Och jag besvor dem vid Gud och sade: »I skolen icke giva edra döttrar åt deras söner, ej heller skolen I av deras döttrar taga hustrur åt edra söner eller åt eder själva.
Var det icke med sådant som Salomo, Israels konung, försyndade sig?
Det fanns bland de många folken ingen konung som var hans like, ty han var älskad av sin Gud, och Gud satte honom till konung över hela Israel.
Likväl kommo de främmande kvinnorna också honom att synda.
Och nu skulle vi om eder få höra att I haven gjort allt detta stora onda och varit otrogna mot vår Gud, i det att I haven tagit till eder främmande kvinnor!»
Och en son till Jojada, översteprästen Eljasibs son, var måg till horoniten Sanballat; honom drev jag bort ifrån mig.
Tänk på dem, min Gud, därför att de hava befläckat prästadömet och prästadömets och leviternas förbund!
Så renade jag folket ifrån allt främmande väsen; och jag fastställde vad prästerna och leviterna skulle iakttaga, var och en i sin syssla,
och huru vedoffret på bestämda tider skulle avlämnas, och huru med förstlingsgåvorna skulle förfaras.
Tänk härpå, min Gud, och räkna mig det till godo!
I Ahasveros' tid -- den Ahasveros' som regerade från Indien ända till Etiopien, över ett hundra tjugusju hövdingdömen --
under den tiden, medan konung Ahasveros satt på konungatronen i Susans borg, tilldrog sig följande.
I sitt tredje regeringsår gjorde han ett gästabud för alla sina furstar och tjänare, varvid Persiens och Mediens härförare och hans förnämsta män och furstarna i hövdingdömena voro samlade inför honom.
Och han lät dem under många dagar se sin konungsliga härlighet och rikedom och sin storhets glans och prakt -- under ett hundra åttio dagar.
Och när dessa dagar hade gått till ända, gjorde konungen ett sju dagars gästabud för allt det folk som fanns i Susans borg, både stora och små, i den inhägnade trädgård som hörde till konungapalatset.
Där hängde tapeter av linne, bomull och mörkblått tyg, uppsatta med vita och purpurröda snören i ringar av silver och på pelare av vit marmor.
Soffor av guld och silver stodo på ett golv som var inlagt med grön och vit marmor och med pärlglänsande och svart sten.
Och dryckerna sattes fram i gyllene kärl, det ena icke likt det andra, och konungsligt vin fanns i myckenhet, såsom det hövdes hos en konung.
Och när man drack, gällde den lagen att intet tvång skulle råda; ty konungen hade befallt alla sina hovmästare att de skulle rätta sig efter vars och ens önskan.
Samtidigt gjorde ock Vasti, drottningen, ett gästabud för kvinnorna i konung Ahasveros' kungliga palats.
När då på sjunde dagen konungens hjärta var glatt av vinet, befallde han Mehuman, Bisseta, Harebona, Bigeta, Abageta, Setar och Karkas, de sju hovmän som gjorde tjänst hos konung Ahasveros,
att de skulle föra drottning Vasti, prydd med kunglig krona, inför konungen, för att han skulle låta folken och furstarna se hennes skönhet, ty hon var fager att skåda.
Men drottning Vasti ville icke komma, fastän konungen befallde henne det genom hovmännen.
Då blev konungen mycket förtörnad. och hans vrede upptändes.
Och konungen frågade de vise som voro kunniga i tidstecknens tydning (ty konungens ärenden plägade så läggas fram för alla i lag och rätt kunniga;
och han hade vid sin sida Karsena, Setar, Admata, Tarsis, Meres, Marsena och Memukan, de sju furstar i Persien och Medien, som voro konungens närmaste män och innehade främsta platsen i riket); han frågade:
»Vad skall man efter lag göra med drottning Vasti, då hon nu icke har gjort vad konung Ahasveros befallde genom hovmännen?»
Memukan svarade inför konungen och furstarna: »Icke mot konungen allena har drottning Vasti gjort illa, utan mot alla furstar och alla folk i alla konung Ahasveros' hövdingdömen.
Ty vad drottningen har gjort skall komma ut bland alla kvinnor, och skall leda till att de förakta sina män, då de ju kunna säga: 'Konung Ahasveros befallde att man skulle föra drottning Vasti inför honom, men hon kom icke.'
Ja, redan i dag skola furstinnorna i Persien och Medien, när de få höra vad drottningen har gjort, åberopa detta inför alla konungens furstar, och därav skall komma förakt och förtret mer än nog.
Om det så täckes konungen, må han därför låta en kunglig befallning utgå -- och må denna upptecknas i Persiens och Mediens lagar, så att den bliver orygglig -- att Vasti icke mer skall få komma inför konung Ahasveros' ansikte; och hennes konungsliga värdighet give konungen åt en annan, som är bättre än hon.
När så den förordning som konungen utfärdar bliver kunnig i hela hans rike, så stort det är, då skola alla kvinnor giva sina män tillbörlig ära, både stora och små.»
Detta tal behagade konungen och furstarna, och konungen gjorde såsom Memukan hade sagt.
Skrivelser blevo sända till alla konungens hövdingdömen, till vart hövdingdöme med dess skrift och till vart folk på dess tungomål, att envar man skulle vara herre i sitt hus och tala sitt folks tungomål.
Efter en tids förlopp, sedan konung Ahasveros' vrede hade lagt sig, tänkte han åter på Vasti och vad hon hade gjort, och vad som var beslutet om henne.
Då sade konungens män som betjänade honom: »Må man för konungens räkning söka upp unga och fagra jungfrur,
och må konungen i sitt rikes alla hövdingdömen förordna vissa män som samla tillhopa alla dessa unga och fagra jungfrur till fruhuset i Susans borg och överlämna dem åt konungens hovman Hege, kvinnovaktaren, och man give dem vad nödigt är till deras beredelse.
Och den kvinna som konungen finner behag i blive drottning i Vastis ställe.»
Detta tal behagade konungen, och han gjorde så.
I Susans borg fanns då en judisk man som hette Mordokai, son till Jair, son till Simei, son till Kis, en benjaminit;
denne hade blivit bortförd från Jerusalem med de fångar som fördes bort tillsammans med Jekonja, Juda konung, när denne fördes bort av Nebukadnessar, konungen i Babel.
Han var fosterfader åt Hadassa, som ock kallades Ester, hans farbroders dotter; ty hon hade varken fader eller moder.
Hon var en flicka med skön gestalt, fager att skåda; och efter hennes faders och moders död hade Mordokai upptagit henne såsom sin egen dotter.
Då nu konungens befallning och påbud blev kunnigt, och många unga kvinnor samlades tillhopa till Susans borg och överlämnades åt Hegai, blev ock Ester hämtad till konungshuset och överlämnad åt kvinnovaktaren Hegai.
Och flickan behagade honom och fann nåd inför honom; därför skyndade han att giva henne vad nödigt var till hennes beredelse, så ock den kost hon skulle hava, ävensom att giva henne från konungshuset de sju tärnor som utsågos åt henne.
Och han lät henne med sina tärnor flytta in i den bästa delen av fruhuset.
Men om sitt folk och sin släkt hade Ester icke yppat något, ty Mordokai hade förbjudit henne att yppa något därom.
Och Mordokai gick var dag fram och åter utanför gården till fruhuset, för att få veta huru det stod till med Ester, och vad som vederfors henne.
Nu var det så, att när ordningen kom till den ena eller andra av de unga kvinnorna att gå in till konung Ahasveros, sedan med henne hade förfarits i tolv månader såsom det var påbjudet om kvinnorna (så lång tid åtgick nämligen till att bereda dem: sex månader med myrraolja och sex månader med välluktande kryddor och annat som var nödigt till kvinnornas beredelse),
när alltså en kvinna gick in till konungen, då fick hon taga med sig ifrån fruhuset till konungshuset allt vad hon begärde.
Och sedan hon om aftonen hade gått ditin, skulle hon om morgonen, när hon gick tillbaka, gå in i det andra fruhuset och överlämnas åt konungens hovman Saasgas, som hade vakten över bihustrurna.
Hon fick sedan icke mer komma in till konungen, om icke konungen hade funnit sådant behag i henne, att hon uttryckligen blev kallad till honom.
Då nu ordningen att gå in till konungen kom till Ester, dotter till Abihail, farbroder till Mordokai, som hade upptagit henne till sin dotter, begärde hon intet annat än det som konungens hovman Hegai, kvinnovaktaren, rådde henne till.
Och Ester fann nåd för allas ögon, som sågo henne.
Ester blev hämtad till konung Ahasveros i hans kungliga palats i tionde månaden, det är månaden Tebet, i hans sjunde regeringsår.
Och Ester blev konungen kärare än alla de andra kvinnorna, och hon fann nåd och ynnest inför honom mer än alla de andra jungfrurna, så att han satte en kunglig krona på hennes huvud och gjorde henne till drottning i Vastis ställe.
Och konungen gjorde ett stort gästabud för alla sina furstar och tjänare, ett gästabud till Esters ära; och han beviljade skattelindring åt sina hövdingdömen och delade ut skänker, såsom det hövdes en konung.
När sedermera jungfrur för andra gången samlades tillhopa och Mordokai satt i konungens port
(men Ester hade, såsom Mordokai bjöd henne, icke yppat något om sin släkt och sitt folk, ty Ester gjorde efter Mordokais befallning, likasom när hon var under hans vård),
vid den tiden, under det att Mordokai satt i konungens port, blevo Bigetan och Teres, två av de hovmän hos konungen, som höllo vakt vid tröskeln, förbittrade på konung Ahasveros och sökte tillfälle att bära hand på honom.
Härom fick Mordokai kunskap, och han berättade det för drottning Ester; därefter omtalade Ester det för konungen på Mordokais vägnar.
Saken blev nu undersökt och så befunnen; och de blevo båda upphängda på trä.
Och detta upptecknades i krönikan, för konungen.
En tid härefter upphöjde konung Ahasveros agagiten Haman, Hammedatas son, till hög värdighet och gav honom främsta platsen bland alla de furstar som voro hos honom.
Och alla konungens tjänare som voro i konungens port böjde knä och föllo ned för Haman, ty så hade konungen bjudit om honom.
Men Mordokai böjde icke knä och föll icke ned för honom.
Då sade konungens tjänare som voro i konungens port till Mordokai: »Varför överträder du konungens bud?»
Och när de dag efter dag hade sagt så till honom, utan att han lyssnade till dem, berättade de det för Haman, för att se om Mordokais förklaring skulle få gälla: ty han hade berättat för dem att han var en jude.
När nu Haman såg att Mordokai icke böjde knä eller föll ned för honom, uppfylldes han med vrede.
Men det syntes honom för ringa att bära hand allenast på Mordokai, sedan man berättat för honom av vilket folk Mordokai var, utan Haman sökte tillfälle att utrota alla judar som funnos i Ahasveros' hela rike, därför att de voro Mordokais landsmän.
I första månaden, det är månaden Nisan, i Ahasveros' tolfte regeringsår, kastades pur , det är lott , inför Haman om var särskild dag och var särskild månad intill tolfte månaden, det är månaden Adar.
Och Haman sade till konung Ahasveros: »Här finnes ett folk som bor kringspritt och förstrött bland de andra folken i ditt rikes alla hövdingdömen.
Deras lagar äro olika alla andra folks, och de göra icke efter konungens lagar; därför är det icke konungen värdigt att låta dem vara.
Om det så täckes konungen, må fördenskull en skrivelse utfärdas, att man skall förgöra dem.
Tio tusen talenter silver skall jag då kunna väga upp åt tjänstemännen till att läggas in i konungens skattkamrar.»
Då tog konungen ringen av sin hand och gav den åt agagiten Haman, Hammedatas son, judarnas ovän.
Därefter sade konungen till Haman: »Silvret vare dig skänkt, och med folket må du göra såsom du finner för gott.»
Så blevo då konungens sekreterare tillkallade på trettonde dagen i första månaden, och en skrivelse, alldeles sådan som Haman ville, utfärdades till konungens satraper och till ståthållarna över de särskilda hövdingdömena och till furstarna över de särskilda folken, till vart hövdingdöme med dess skrift och till vart folk på dess tungomål.
I konung Ahasveros' namn utfärdades skrivelsen, och den beseglades med konungens ring.
Sedan kringsändes med ilbud brev till alla konungens hövdingdömen, att man skulle utrota, dräpa och förgöra judarna, både unga och gamla, både barn och kvinnor, alla på en och samma dag, nämligen på trettonde dagen i tolfte månaden, det är månaden Adar, varvid ock deras ägodelar såsom byte skulle givas till plundring.
I skrivelsen stod att i vart särskilt hövdingdöme ett påbud, öppet för alla folk, skulle utfärdas, som innehöll att de skulle vara redo den dagen.
Och på grund av konungens befallning drogo ilbuden med hast åstad, så snart påbudet hade blivit utfärdat i Susans borg.
Men konungen och Haman satte sig ned till att dricka, under det att bestörtning rådde i staden Susan.
När Mordokai fick veta allt vad som hade skett, rev han sönder sina kläder och klädde sig i säck och aska, och gick så ut i staden och uppgav högljudda och bittra klagorop.
Och han begav sig till konungens port och stannade framför den, ty in i konungens port fick ingen komma, som var klädd i sorgdräkt.
Och i vart hövdingdöme dit konungens befallning och påbud kom blev stor sorg bland judarna, och de fastade, gräto och klagade, ja, de flesta satte sig i säck och aska.
När nu Esters tjänarinnor och hovmän kommo och berättade detta för henne, blev drottningen högeligen förskräckt; och hon skickade ut kläder till Mordokai, för att man skulle kläda honom i dem och taga av honom sorgdräkten; men han tog icke emot dem.
Då kallade Ester till sig Hatak, en av de hovmän som konungen hade anställt i hennes tjänst, och bjöd honom att gå till Mordokai, för att få veta vad som var på färde, och varför han gjorde så.
När då Hatak kom ut till Mordokai på den öppna platsen i staden framför konungens port,
berättade Mordokai för honom allt vad som hade hänt honom, och uppgav beloppet av den penningsumma som Haman hade lovat väga upp till konungens skattkamrar, för att han skulle få förgöra judarna.
Och en avskrift av det skrivna påbud som hade blivit utfärdat i Susan om att de skulle utrotas lämnade han honom ock, för att han skulle visa Ester den och berätta allt för henne, och ålägga henne att gå in till konungen och bedja honom om misskund och söka nåd hos honom för sitt folk.
Och Hatak kom och berättade för Ester vad Mordokai hade sagt.
Då bjöd Ester Hatak att gå till Mordokai och säga:
»Alla konungens tjänare och folket i konungens hövdingdömen veta, att om någon, vare sig man eller kvinna, går in till konungen på den inre gården utan att vara kallad, så gäller för var och en samma lag: att han skall dödas, såframt icke konungen räcker ut mot honom den gyllene spiran, till tecken på att han får leva.
Men jag har icke på trettio dagar varit kallad att komma till konungen.»
När man nu berättade för Mordokai vad Ester hade sagt,
sade Mordokai att man skulle giva Ester detta svar: »Tänk icke att du ensam bland alla judar skall slippa undan, därför att du är i konungens hus.
Nej, om du tiger stilla vid detta tillfälle, så skall nog hjälp och räddning beredas judarna från något annat håll, men du och din faders hus, I skolen förgöras.
Vem vet om du icke just för en sådan tid som denna har kommit till konungslig värdighet?»
Då lät Ester giva Mordokai detta svar:
»Gå åstad och församla alla judar som finnas i Susan, och hållen fasta för mig; I skolen icke äta eller dricka något under tre dygn, vare sig dag eller natt.
Jag med mina tärnor vill ock sammalunda fasta; därefter vill jag gå in till konungen, fastän det är emot lagen.
Och skall jag gå förlorad, så må det då ske.»
Och Mordokai gick bort och gjorde alldeles såsom Ester hade bjudit honom.
På tredje dagen klädde Ester sig i konungslig skrud och trädde in på den inre gården till konungshuset, mitt emot själva konungshuset; konungen satt då på sin konungatron i det kungliga palatset, mitt emot palatsets dörr.
När nu konungen såg drottning Ester stå på gården, fann hon nåd för hans ögon, så att konungen räckte ut mot Ester den gyllene spira, som han hade i sin hand; då gick Ester fram och rörde vid ändan av spiran.
Och konungen sade till henne: »Vad önskar du, drottning Ester, och vad är din begäran?
Gällde den ock hälften av riket, så skall den beviljas dig.»
Ester svarade: »Om det så täckes konungen, må konungen jämte Haman i dag komma till ett gästabud, som jag har tillrett för honom.»
Då sade konungen: »Skynden att hämta hit Haman, för att så må ske, som Ester har begärt.»
Så kommo då konungen och Haman till gästabudet, som Ester hade tillrett.
Och när vinet dracks, sade konungen till Ester: »Vad är din bön?
Den vare dig beviljad.
Och vad är din begäran?
Gällde den ock hälften av riket, så skall den uppfyllas.»
Ester svarade och sade: »Min bön och min begäran är:
om jag har funnit nåd för konungens ögon, och det täckes konungen att bevilja min bön och uppfylla min begäran, så må konungen och Haman komma till ännu ett gästabud, som jag vill tillreda för dem; då skall jag i morgon göra såsom konungen har befallt.»
Och Haman gick därifrån den dagen, glad och väl till mods.
Men när han fick se Mordokai i konungens port och denne varken stod upp eller ens rörde sig för honom, då uppfylldes Haman med vrede mot Mordokai.
Men Haman betvang sig och gick hem; därefter sände han och lät hämta sina vänner och sin hustru Seres.
Och Haman talade för dem om sin rikedom och härlighet och om sina många barn och om all den storhet, som konungen hade givit honom, och om huru konungen i allt hade upphöjt honom över de andra furstarna och konungens övriga tjänare.
Och Haman sade ytterligare: »Icke heller har drottning Ester låtit någon annan än mig komma med konungen till det gästabud, som hon hade tillrett; och jämväl i morgon är jag bjuden till henne, jämte konungen.
Men vid allt detta kan jag dock icke vara till freds, så länge jag ser juden Mordokai sitta i konungens port.»
Då sade hans hustru Seres och alla hans vänner till honom: »Låt resa upp en påle, femtio alnar hög, och bed i morgon konungen, att Mordokai må bliva upphängd därpå; då kan du glad komma med konungen till gästabudet.»
Detta behagade Haman, och han lät resa upp pålen.
Den natten kunde konungen icke sova; därför lät han hämta krönikan, där minnesvärda händelser voro upptecknade, och man föreläste ur den för konungen.
Då fann man där skrivet, att Mordokai hade berättat, hurusom Bigetana och Teres, två av de hovmän, som höllo vakt vid tröskeln, hade sökt tillfälle att bära hand på konung Ahasveros.
Konungen frågade: »Vilken ära och upphöjelse har vederfarits Mordokai för detta?»
Konungens män, som betjänade honom, svarade: »Intet sådant har vederfarits honom.»
Då sade konungen: »Är någon nu tillstädes på gården?»
Och Haman hade just kommit in på den yttre gården till konungshuset för att bedja konungen, att Mordokai måtte bliva upphängd på den påle, som han hade låtit sätta upp för hans räkning.
Så svarade honom då konungens tjänare: »Ja, Haman står därute på gården.»
Konungen sade: »Låt honom komma in.»
När då Haman kom in, sade konungen till honom: »Huru skall man göra med den man, som konungen vill ära?»
Men Haman tänkte i sitt hjärta: »Vem skulle konungen vilja bevisa ära mer än mig?»
Därför sade Haman till konungen: »Om konungen vill ära någon,
så skall man hämta en konungslig klädnad, som konungen själv har burit, och en häst, som konungen själv har ridit på, och på vilkens huvud en kunglig krona är fäst;
och man skall överlämna klädnaden och hästen åt en av konungens förnämsta furstar, och klädnaden skall sättas på den man, som konungen vill ära, och man skall föra honom ridande på hästen fram på den öppna platsen i staden och utropa framför honom: 'Så gör man med den man, som konungen vill ära.'»
Då sade konungen till Haman: »Skynda dig att taga klädnaden och hästen, såsom du har sagt, och gör så med juden Mordokai, som sitter i konungens port.
Underlåt intet av allt vad du har sagt.»
Så tog då Haman klädnaden och hästen och satte klädnaden på Mordokai och förde honom ridande fram på den öppna platsen i staden och utropade framför honom: »Så gör man med den man, som konungen vill ära.»
Och Mordokai vände tillbaka till konungens port; men Haman skyndade hem, sörjande och med överhöljt huvud.
Och när Haman förtäljde för sin hustru Seres och alla sina vänner vad som hade hänt honom, sade hans vise män och hans hustru Seres till honom: »Om Mordokai, som du har begynt att stå tillbaka för, är av judisk börd, så förmår du intet mot honom, utan skall komma alldeles till korta för honom.»
Medan de ännu så talade med honom, kommo konungens hovmän för att skyndsamt hämta Haman till gästabudet, som Ester hade tillrett.
Så kommo då konungen och Haman till gästabudet hos drottning Ester.
Och när vinet dracks, sade konungen till Ester, också nu på andra dagen: »Vad är din bön, drottning Ester?
Den vare dig beviljad.
Och vad är din begäran?
Gällde den ock hälften av riket, så skall den uppfyllas.»
Drottning Ester svarade och sade: »Om jag har funnit nåd för dina ögon, o konung, och det så täckes konungen, så blive mitt liv mig skänkt på min bön, och mitt folks på min begäran.
Ty vi äro sålda, jag och mitt folk, till att utrotas, dräpas och förgöras.
Om vi allenast hade blivit sålda till trälar och trälinnor, så skulle jag hava tegat; ty den olyckan vore icke sådan, att vi borde besvära konungen därmed.»
Då svarade konung Ahasveros och sade till drottning Ester: »Vem är den, och var är den, som har fördristat sig att så göra?»
Ester sade: »En hätsk och illvillig man är det: den onde Haman där.»
Då blev Haman förskräckt för konungen och drottningen.
Och konungen stod upp i vrede och lämnade gästabudet och gick ut i palatsets trädgård; men Haman trädde fram för att bedja drottning Ester om sitt liv, ty han såg, att konungen hade beslutit hans ofärd.
När konungen därefter kom tillbaka till gästabudssalen från palatsets trädgård, hade Haman sjunkit ned mot den soffa, där Ester satt; då sade konungen: »Vill han ock öva våld mot drottningen, härinne i min närvaro?»
Knappt hade detta ord gått över konungens läppar, förrän man höljde över Hamans ansikte.
Och Harebona, en av hovmännen hos konungen, sade: »Vid Hamans hus står redan en påle, femtio alnar hög, som Haman låtit resa upp för Mordokai, vilkens ord en gång var konungen till sådant gagn.»
Då sade konungen: »Hängen upp honom på den.»
Så hängde de upp Haman på den påle, som han hade låtit sätta upp för Mordokai.
Sedan lade sig konungens vrede.
Samma dag gav konung Ahasveros åt drottning Ester Hamans, judarnas oväns, hus.
Och Mordokai fick tillträde till konungen, ty Ester hade nu omtalat, vad han var för henne.
Och konungen tog av sig ringen, som han hade låtit taga ifrån Haman, och gav den åt Mordokai.
Och Ester satte Mordokai över Hamans hus.
Och Ester talade ytterligare inför konungen, i det att hon föll ned för hans fötter; hon bönföll honom gråtande, att han skulle avvända agagiten Hamans onda råd och det anslag, som denne hade förehaft mot judarna.
Då räckte konungen ut den gyllene spiran mot Ester; och Ester stod upp och trädde fram inför konungen
och sade: »Om det så täckes konungen, och om jag har funnit nåd inför honom, och det synes konungen vara riktigt och jag är honom till behag, så må en skrivelse utfärdas för att återkalla de brev, som innehöllo agagiten Hamans, Hammedatas sons, anslag, och som han skrev för att förgöra judarna i alla konungens hövdingdömen.
Ty huru skulle jag kunna uthärda att se den olycka, som eljest träffade mitt folk?
Ja, huru skulle jag kunna uthärda att se mina landsmän förgöras?»
Då sade konung Ahasveros till drottning Ester och till juden Mordokai: »Se, Hamans hus har jag givit åt Ester, och han själv har blivit upphängd på en påle, därför att han ville bära hand på judarna.
Men utfärden nu ock I en skrivelse angående judarna i konungen namn, såsom I finnen för gott, och beseglen den med konungens ring.
Ty en skrivelse, som är utfärdad i konungens namn och beseglad med konungens ring, kan icke återkallas.»
Så blevo nu strax konungens sekreterare tillkallade, på tjugutredje dagen i tredje månaden, det är månaden Sivan, och en skrivelse, alldeles sådan som Mordokai ville, utfärdades till judarna och till satraperna, ståthållarna och furstarna i hövdingdömena, från Indien ända till Etiopien, ett hundra tjugusju hövdingdömen, till vart hövdingdöme med dess skrift och till vart folk på dess tungomål, jämväl till judarna med deras skrift och på deras tungomål.
Han utfärdade skrivelsen i konung Ahasveros' namn och beseglade den med konungens ring.
Därefter kringsände han brev med ilbud till häst, som redo på kungliga travare från stuterierna,
att konungen tillstadde judarna i var särskild stad att församla sig till försvar för sitt liv och att i vart folk och hövdingdöme utrota, dräpa och förgöra alla väpnade skaror, som angrepe dem, ävensom barn och kvinnor, varvid deras ägodelar såsom byte skulle givas till plundring,
detta på en och samma dag i alla konung Ahasveros' hövdingdömen, nämligen på trettonde dagen i tolfte månaden, det är månaden Adar.
I skrivelsen stod, att i vart särskilt hövdingdöme ett påbud, öppet för alla folk, skulle utfärdas, som innehöll, att judarna skulle vara redo till den dagen att hämnas på sina fiender.
Och på grund av konungens befallning drogo ilbuden på de kungliga travarna skyndsamt och med hast åstad, så snart påbudet hade blivit utfärdat i Susans borg.
Men Mordokai gick ut från konungen i konungslig klädnad av mörkblått och vitt tyg och med en stor gyllene krona och en mantel av vitt och purpurrött tyg, under det att staden Susan jublade och var glad.
För judarna hade nu uppgått ljus och glädje, fröjd och ära.
Och i vart hövdingdöme och i var stad, dit konungens befallning och påbud kom, blev glädje och fröjd bland judarna, och de höllo gästabud och högtid.
Och många ur de främmande folken blevo judar, ty förskräckelse för judarna hade fallit över dem.
På trettonde dagen i tolfte månaden, det är månaden Adar, den dag då konungens befallning och påbud skulle verkställas, och då judarnas fiender hade hoppats att bliva dem övermäktiga -- fastän det vände sig så, att judarna i stället skulle bliva sina motståndare övermäktiga --
på den dagen församlade sig judarna i sina städer, i alla konung Ahasveros' hövdingdömen, för att kasta sig över dem, som sökte deras ofärd; och ingen kunde stå dem emot, ty förskräckelse för dem hade fallit över alla folk.
Och alla furstarna i hövdingdömena och satraperna och ståthållarna och konungens tjänstemän understödde judarna, ty förskräckelse för Mordokai hade fallit över dem.
Ty Mordokai var nu stor i konungens hus, och hans rykte gick ut i alla hövdingdömen, eftersom denne Mordokai lev allt större och större.
Och judarna anställde med sina svärd ett nederlag överallt bland sina fiender och dräpte och förgjorde dem och förforo såsom de ville med sina motståndare.
I Susans borg dräpte och förgjorde judarna fem hundra män.
Och Parsandata, Dalefon, Aspata,
Porata, Adalja, Aridata,
Parmasta, Arisai, Aridai och Vajsata,
judarnas ovän Hamans, Hammedatas sons, tio söner dräpte de; men till plundring räckte de icke ut sin hand.
Samma dag fick konungen veta huru många som hade blivit dräpta i Susans borg.
Då sade konungen till drottning Ester: »I Susans borg hava judarna dräpt och förgjort fem hundra män utom Hamans tio söner; vad skola de då icke hava gjort i konungens övriga hövdingdömen?
Vad är nu din bön?
Den vare dig beviljad.
Och vad är ytterligare din begäran?
Den skall uppfyllas.»
Ester svarade: »Om det så täckes konungen, så må det också i morgon tillstädjas de judar, som äro i Susan, att göra efter påbudet för i dag; och må Hamans tio söner bliva upphängda på pålen.»
Då befallde konungen, att så skulle ske, och påbudet blev utfärdat i Susan; därefter blevo Hamans tio söner upphängda.
och de judar, som voro i Susan, församlade sig också på fjortonde dagen i månaden Adar och dräpte i Susan tre hundra män; men till plundring räckte de icke ut sin hand.
Och de övriga judarna, de som voro i konungen hövdingdömen, församlade sig till försvar för sitt liv och skaffade sig ro för sina fiender, i det att dräpte sjuttiofem tusen av dessa sina motståndare; men till plundring räckte de icke ut sin hand.
Detta skedde på trettonde dagen i månaden Adar; men på fjortonde dagen vilade de och firade den såsom en gästabuds- och glädjedag.
De judar åter, som voro i Susan, hade församlat sig både den trettonde dagen och på den fjortonde; men de vilade på den femtonde dagen och firade den såsom en gästabuds- och glädjedag.
Därför fira judarna på landsbygden, de som bo i landsortsstäderna, den fjortonde dagen i månaden Adar såsom en glädje-, gästabuds- och högtidsdag, på vilken de sända gåvor till varandra av den mat de hava tillagat.
Och Mordokai tecknade upp dessa händelser och sände skrivelser till alla judar i konung Ahasveros' hövdingdömen, både nära och fjärran,
och stadgade såsom lag för dem, att de alltid, år efter år, skulle fira den fjortonde och den femtonde dagen i månaden Adar,
eftersom det var på dessa dagar som judarna hade fått ro för sina fiender, och eftersom i denna månad deras bedrövelse hade blivit förvandlad till glädje och deras sorg till högtid.
Därför skulle de fira dessa dagar såsom gästabuds- och glädjedagar, på vilka de skulle sända gåvor till varandra av den mat de hade tillagat, så ock skänker till de fattiga.
Och judarna antogo såsom sed, vad de nu hade begynt att göra, det varom Mordokai hade skrivit till dem --
detta eftersom agagiten Haman, Hammedatas son, alla judars ovän, hade förehaft sitt anslag mot judarna till att förgöra dem och hade kastat pur , det är lott , till att plötsligt överfalla och förgöra dem;
varemot konungen, när han hade fått veta detta, hade givit befallning och utfärdat en skrivelse om att det onda anslag, som denne hade förehaft mot judarna, skulle vända tillbaka på hans eget huvud, så att han själv och hans söner hade blivit upphängda på pålen.
Fördenskull blevo dessa dagar kallade purim efter ordet pur ; och fördenskull, i anledning av allt som stod i detta brev, och vad de själva härav hade sett, och vad som hade vederfarits dem,
stadgade judarna och antogo såsom orygglig sed för sig och sina efterkommande och för alla, som slöto sig till dem, att alltid, år efter år, fira dessa båda dagar, efter föreskriften om dem och på den för dem bestämda tiden,
och att dessa dagar skulle ihågkommas och firas i alla tider, i var släkt, i vart hövdingdöme och i var stad, så att dessa purimsdagar oryggligt skulle hållas bland judarna och deras åminnelse icke upphöra bland deras efterkommande.
Men drottning Ester, Abihails dotter, och juden Mordokai uppsatte ånyo en skrivelse, i eftertryckliga ordalag, för att stadga såsom en lag, vad som föreskrevs i detta nya brev om purim.
Och skrivelser, vänligt och välvilligt avfattade, utsändes till alla judar i de ett hundra tjugusju hövdingdömena i Ahasveros' rike,
för att stadga såsom lag, att de skulle fira dessa purimsdagar på deras bestämda tider så, som juden Mordokai och drottning Ester stadgade för dem, och så, som de stadgade för sig själva och sina efterkommande, nämligen med föreskrivna fastor och övliga klagorop.
Alltså blevo genom Esters befallning dessa föreskrifter om purim stadgade såsom lag; och den tecknades upp i en bok.
Och konung Ahasveros tog skatt både av fastlandet och av öarna i havet.
Och allt vad han i sin makt och sin väldighet gjorde, ävensom berättelsen om den storhet, till vilken konungen upphöjde Mordokai, det finnes upptecknat i de mediska och persiska konungarnas krönika.
Ty juden Mordokai var konung Ahasveros' närmaste man, och han var stor bland judarna och älskad av alla sina bröder, eftersom han sökte sitt folks bästa och lade sig ut för alla sina landsmän till deras välfärd.
I Us' land levde en man som hette Job; han var en ostrafflig och redlig man, som fruktade Gud och flydde det onda.
Åt honom föddes sju söner och tre döttrar;
och han ägde sju tusen får, tre tusen kameler, fem hundra par oxar och fem hundra åsninnor, därtill tjänare i stor mängd.
Så var denne man mäktigare än någon annan i Österlandet.
Och hans söner hade för sed att gå åstad och hålla gästabud, den ena dagen i den enes hus, den andra dagen i den andres; de sände då och inbjödo sina tre systrar att äta och dricka tillsammans med dem.
När så en omgång av gästabudsdagar var till ända, sände Job efter dem för att helga dem; bittida om morgonen offrade han då ett brännoffer för var och en av dem.
Ty Job tänkte »Kanhända hava mina barn syndat och i sina hjärtan talat förgripligt om Gud».
Så gjorde Job för var gång.
Men nu hände sig en dag att Guds söner kommo och trädde fram inför HERREN, och Åklagaren kom också med bland dem.
Då frågade HERREN Åklagaren: »Varifrån kommer du?»
Åklagaren svarade HERREN och sade: »Från en vandring utöver jorden och från en färd omkring på den.»
Då sade HERREN till Åklagaren: »Har du givit akt på min tjänare Job?
Ty på jorden finnes icke hans like i ostrafflighet och redlighet, ingen som så fruktar Gud och flyr det onda.»
Åklagaren svarade HERREN och sade: »Är det då för intet som Job fruktar Gud?
Du har ju på allt sätt beskärmat honom och hans hus och allt vad han äger; du har välsignat hans händers verk, och hans boskapshjordar hava utbrett sig i landet.
Man räck ut din hand och kom vid detta allt som han äger; förvisso skall han då mitt i ansiktet tala förgripliga ord mot dig.»
HERREN sade till Åklagaren: »Välan, allt vad han äger vare givet i din hand; allenast mot honom själv må du icke räcka ut din hand.»
Så gick Åklagaren bort ifrån HERRENS ansikte.
När nu en dag hans söner och döttrar höllo måltid och drucko vin i den äldste broderns hus,
Kom en budbärare till Job och sade: »Oxarna gingo för plogen, och åsninnorna betade därbredvid;
då föllo sabéerna in och rövade bort dem, och folket slogo de med svärdsegg.
Jag var den ende som kom undan, för att jag skulle underrätta dig därom.»
Medan denne ännu talade, kom åter en och sade: »Guds eld föll ifrån himmelen och slog ned bland småboskapen och folket och förtärde dem.
Jag var den ende som kom undan, för att jag skulle underrätta dig därom.»
Medan denne ännu talade, kom åter en och sade: Kaldéerna ställde upp sitt manskap i tre hopar och föllo så över kamelerna och rövade bort dem, och folket slogo de med svärdsegg.
Jag var den ende som kom undan, för att jag skulle underrätta dig därom.»
Under det att denne ännu talade, kom åter en annan och sade: Dina söner och döttrar höllo måltid och drucko vin i den äldste broderns hus;
då kom en stark storm fram över öknen och tog tag i husets fyra hörn, och det föll omkull över folket, så att de förgingos.
Jag var den ende som kom undan, för att jag skulle underrätta dig därom.»
Då stod Job upp och rev sönder sin mantel och skar av håret på sitt huvud.
Och han föll ned till jorden och tillbad
och sade: »Naken kom jag ur min moders liv, och naken skall jag vända åter dit; HERREN gav, och HERREN tog.
Lovat vare HERRENS namn!»
Vid allt detta syndade Job icke och talade intet lasteligt mot Gud.
Åter hände sig en dag att Guds söner kommo och trädde fram inför HERREN; och Åklagaren kom också med bland dem och trädde fram inför HERREN.
Då frågade HERREN Åklagaren: »Varifrån kommer du?»
Åklagaren svarade HERREN och sade: »Från en vandring utöver jorden och från en färd omkring på den.»
Då sade HERREN till Åklagaren: »Har du givit akt på min tjänare Job?
Ty på jorden finnes icke hans like i ostrafflighet och redlighet, ingen som så fruktar Gud och flyr det onda; och ännu håller han fast vid sin ostrafflighet.
Så har du då uppeggat mig mot honom till att utan sak fördärva honom.»
Åklagaren svarade HERREN och sade: »Hud för hud; allt vad man äger giver man ju för att själv slippa undan.
Men räck ut din hand och kom vid hans kött och ben; förvisso skall han då mitt i ansiktet tala förgripliga ord mot dig.»
HERREN sade till Åklagaren: »Välan, han vare given i din hand; allenast hans liv må du skona.»
Så gick Åklagaren bort ifrån HERRENS ansikte och slog Job med svåra bulnader, ifrån fotbladet ända till hjässan.
Och han tog sig en lerskärva att skrapa sig med, där han satt mitt i askan.
Då sade hans hustru till honom: »Håller du ännu fast vid din ostrafflighet?
Tala fritt ut om Gud, och dö.»
Man han svarade henne: »Du talar såsom en dåraktig kvinna skulle tala.
Om vi taga emot det goda av Gud, skola vi då icke också taga emot det onda?»
Vid allt detta syndade Job icke med sina läppar.
Men tre vänner till Job fingo höra om alla de olyckor som hade träffat honom, och de kommo så, var och en från sin ort; Elifas från Teman, Bildad från Sua och Sofar från Naama.
Och de avtalade med varandra att de skulle begiva sig åstad för att ömka honom och trösta honom.
Men när de, ännu på avstånd, lyfte upp sina ögon och sågo att de icke mer kunde känna igen honom, brusto de ut i gråt och revo sönder sina mantlar och kastade stoft mot himmelen, ned över sina huvuden.
Sedan sutto de med honom på jorden i sju dagar och sju nätter, utan att någon av dem talade ett ord till honom, eftersom de sågo att hans plåga var mycket stor.
Därefter upplät Job sin mun och förbannade sin födelsedag;
Job tog till orda och sade:
Må den dag utplånas, på vilken jag föddes, och den natt som sade: »Ett gossebarn är avlat.»
Må den dagen vändas i mörker, må Gud i höjden ej fråga efter den och intet dagsljus lysa däröver.
Mörkret och dödsskuggan börde den åter, molnen lägre sig över den; förskräcke den allt som kan förmörka en dag.
Den natten må gripas av tjockaste mörker; ej må den få fröjda sig bland årets dagar, intet rum må den finna inom månadernas krets.
Ja, ofruktsam blive den natten, aldrig höje sig jubel under den.
Må den förbannas av dem som besvärja dagar, av dem som förmå mana upp Leviatan.
Må dess grynings stjärnor förmörkas, efter ljus må den bida, utan att det kommer, morgonrodnadens ögonbryn må den aldrig få se;
eftersom den ej tillslöt dörrarna till min moders liv, ej lät olyckan förbliva dold för mina ögon.
Varför fick jag ej dö strax i modersskötet, förgås vid det jag kom ut ur min moders liv?
Varför funnos knän mig till mötes, och varför bröst, där jag fick di?
Hade så icke skett, låge jag nu i ro, jag finge då sova, jag njöte då min vila,
vid sidan av konungar och rådsherrar i landet, män som byggde sig palatslika gravar,
ja, vid sidan av furstar som voro rika på guld och hade sina hus uppfyllda av silver;
eller vore jag icke till, lik ett nedgrävt foster, lik ett barn som aldrig fick se ljuset.
Där hava ju de ogudaktiga upphört att rasa, där få de uttröttade komma till vila;
där hava alla fångar fått ro, de höra där ingen pådrivares röst.
Små och stora äro där varandra lika, trälen har där blivit fri ifrån sin herre.
Varför skulle den olycklige skåda ljuset?
Ja, varför gives liv åt dem som plågas så bittert,
åt dem som vänta efter döden, utan att den kommer, och spana därefter mer än efter någon skatt,
åt dem som skulle glädjas -- ja, intill jubel -- och fröjda sig, allenast de funne sin grav;
varför åt en man vilkens väg är höljd i mörker, åt en man så kringstängd av Gud?
Suckan har ju blivit mitt dagliga bröd, och såsom vatten strömma mina klagorop.
ty det som ingav mig förskräckelse, det drabbar mig nu, och vad jag fruktade för, det kommer över mig.
Jag får ingen rast, ingen ro, ingen vila; ångest kommer över mig.
Därefter tog Elifas från Teman till orda och sade:
Misstycker du, om man dristar tala till dig?
Vem kan hålla tillbaka sina ord?
Se, många har du visat till rätta, och maktlösa händer har du stärkt;
dina ord hava upprättat den som stapplade, och åt vacklande knän har du givit kraft.
Men nu, då det gäller dig själv, bliver du otålig, när det är dig det drabbar, förskräckes du.
Skulle då icke din gudsfruktan vara din tillförsikt och dina vägars ostrafflighet ditt hopp?
Tänk efter: när hände det att en oskyldig fick förgås? och var skedde det att de redliga måste gå under?
Nej, så har jag sett det gå, att de som plöja fördärv och de som utså olycka, de skörda och sådant;
för Guds andedräkt förgås de och för en fnysning av hans näsa försvinna de.
Ja, lejonets skri och rytarens röst måste tystna, och unglejonens tänder brytas ut;
Det gamla lejonet förgås, ty det finner intet rov, och lejoninnans ungar bliva förströdda.
Men till mig smög sakta ett ord, mitt öra förnam det likasom en viskning,
När tankarna svävade om vid nattens syner och sömnen föll tung på människorna,
då kom en förskräckelse och bävan över mig, med rysning fyllde den alla ben i min kropp.
En vindpust for fram över mitt ansikte, därvid reste sig håren på min kropp.
Och något trädde inför mina ögon, en skepnad vars form jag icke skönjde; och jag hörde en susning och en röst:
»Kan då en människa hava rätt mot Gud eller en man vara ren inför sin skapare?
Se, ej ens på sina tjänare kan han förlita sig, jämväl sina änglar måste han tillvita fel;
huru mycket mer då dem som bo i hyddor av ler, dem som hava sin grundval i stoftet!
De krossas sönder så lätt som mal;
när morgon har bytts till afton, ligga de slagna; innan man aktar därpå, hava de förgåtts för alltid.
Ja, deras hyddas fäste ryckes bort för dem, oförtänkt måste de dö.»
Ropa fritt; vem finnes, som svarar dig, och till vilken av de heliga kan du vända dig?
Se, dåren dräpes av sin grämelse, och den fåkunnige dödas av sin bitterhet.
Jag såg en dåre, fast var han rotad, men plötsligt måste jag ropa ve över hans boning.
Ty hans barn gå nu fjärran ifrån frälsning, de förtrampas i porten utan räddning.
Av hans skörd äter vem som är hungrig, den rövas bort, om och hägnad med törnen; efter hans rikedom gapar ett giller.
Ty icke upp ur stoftet kommer fördärvet, ej ur marken skjuter olyckan upp;
nej, människan varder född till olycka, såsom eldgnistor måste flyga mot höjden.
Men vore det nu jag, så sökte jag nåd hos Gud, åt Gud hemställde jag min sak,
åt honom som gör stora och outrannsakliga ting, under, flera än någon kan räkna,
åt honom som låter regnet falla på jorden och sänder vatten ned över markerna,
när han vill upphöja de ringa och förhjälpa de sörjande till frälsning.
Han är den som gör de klokas anslag om intet, så att deras händer intet uträtta med förnuft;
han fångar de visa i deras klokskap och låter de illfundiga förhasta sig i sina rådslag:
mitt på dagen råka de ut för mörker och famla mitt i ljuset, likasom vore det natt.
Så frälsar han från deras tungors svärd, han frälsar den fattige ur den övermäktiges hand.
Den arme kan så åter hava ett hopp, och orättfärdigheten måste tillsluta sin mun.
Ja, säll är den människa som Gud agar; den Allsmäktiges tuktan må du icke förkasta.
Ty om han och sargar, så förbinder han ock, om han slår, så hela ock hans händer.
Sex gånger räddar han dig ur nöden, ja, sju gånger avvändes olyckan från dig.
I hungerstid förlossar han dig från döden och i krig undan svärdets våld.
När tungor svänga gisslet, gömmes du undan; du har intet att frukta, när förhärjelse kommer.
Ja, åt förhärjelse och dyr tid kan du då le, för vilddjur behöver du ej heller känna fruktan;
ty med markens stenar står du i förbund, och med djuren på marken har du ingått fred.
Och du får se huru din hydda står trygg; när du synar din boning, saknas intet däri.
Du får ock se huru din ätt förökas, huru din avkomma bliver såsom markens örter.
I graven kommer du, när du har hunnit din mognad, såsom sädesskylen bärgas, då dess tid är inne.
Se, detta hava vi utrannsakat, och så är det; hör därpå och betänk det väl.
Då tog Job till orda och sade:
Ack att min grämelse bleve vägd och min olycka lagd jämte den på vågen!
Se, tyngre är den nu än havets sand, därför kan jag icke styra mina ord.
Ty den Allsmäktiges pilar hava träffat mig, och min ande indricker deras gift; ja, förskräckelser ifrån Gud ställa sig upp mot mig.
Icke skriar vildåsnan, när hon har friskt gräs, icke råmar oxen, då han står vid sitt foder?
Men vem vill äta den mat som ej har smak eller sälta, och vem finner behag i slemörtens saft?
Så vägrar nu min själ att komma vid detta, det är för mig en vämjelig spis.
Ack att min bön bleve hörd, och att Gud ville uppfylla mitt hopp!
O att det täcktes Gud att krossa mig, att räcka ut sin hand och avskära mitt liv!
Då funnes ännu för mig någon tröst, jag kunde då jubla, fastän plågad utan förskoning; jag har ju ej förnekat den Heliges ord.
Huru stor är då min kraft, eftersom jag alltjämt bör hoppas?
Och vad väntar mig för ände, eftersom jag skall vara tålig?
Min kraft är väl ej såsom stenens, min kropp är väl icke av koppar?
Nej, förvisso gives ingen hjälp för mig, var utväg har blivit mig stängd.
Den förtvivlade borde ju röna barmhärtighet av sin vän, men se, man övergiver den Allsmäktiges fruktan,
Mina bröder äro trolösa, de äro såsom regnbäckar, ja, lika bäckarnas rännilar, som snart sina ut,
som väl kunna gå mörka av vinterns flöden, när snön har fallit och gömt sig i dem,
men som åter försvinna, när de träffas av hettan, och torka bort ifrån sin plats, då värmen kommer.
Vägfarande där i trakten vika av till dem, men de finna allenast ödslighet och måste förgås.
Temas vägfarande skådade dithän, Sabas köpmanståg hoppades på dem;
men de kommo på skam i sin förtröstan, de sågo sig gäckade, när de hade hunnit ditfram.
Ja, likaså ären I nu ingenting värda, handfallna stån I av förfäran och förskräckelse.
Har jag då begärt att I skolen giva mig gåvor, taga av edert gods för att lösa mig ut,
att I skolen rädda mig undan min ovän, köpa mig fri ur våldsverkares hand?
Undervisen mig, så vill jag tiga, lären mig att förstå vari jag har farit vilse.
Gott är förvisso uppriktigt tal, men tillrättavisning av eder, vad båtar den?
Haven I då i sinnet att hålla räfst med ord, och skall den förtvivlade få tala för vinden?
Då kasten I väl också lott om den faderlöse, då lären I väl köpslå om eder vän!
Dock, må det nu täckas eder att akta på mig; icke vill jag ljuga eder mitt i ansiktet.
Vänden om!
Må sådan orätt icke ske; ja, vänden ännu om, ty min sak är rättfärdig!
Skulle väl orätt bo på min tunga, och min mun, skulle den ej förstå vad fördärvligt är?
En stridsmans liv lever ju människan på jorden, och hennes dagar äro såsom dagakarlens dagar.
Hon är lik en träl som flämtar efter skugga, lik en dagakarl som får bida efter sin lön.
Så har jag fått till arvedel månader av elände; nätter av vedermöda hava blivit min lott.
Så snart jag har lagt mig, är min fråga: »När skall jag då få stå upp?»
Ty aftonen synes mig så lång; jag är övermätt av oro, innan morgonen har kommit.
Med förruttnelsens maskar höljes min kropp, med en skorpa lik jord; min hud skrymper samman och faller sönder.
Mina dagar fly snabbare än vävarens spole; de försvinna utan något hopp.
Tänk därpå att mitt liv är en fläkt, att mitt öga icke mer skall få se någon lycka.
Den nu ser mig, hans öga skall ej vidare skåda mig; bäst din blick vilar på mig, är jag icke mer.
Såsom ett moln som har försvunnit och gått bort, så är den som har farit ned i dödsriket; han kommer ej åter upp därifrån.
Aldrig mer vänder han tillbaka till sitt hus, och hans plats vet icke av honom mer.
Därför vill jag nu icke lägga band på min mun, jag vill taga till orda i min andes ångest, jag vill klaga i min själs bedrövelse.
Icke är jag väl ett hav eller ett havsvidunder, så att du måste sätta ut vakt mot mig?
När jag hoppas att min bädd skall trösta mig, att mitt läger skall lindra mitt bekymmer,
då förfärar du mig genom drömmar, och med syner förskräcker du mig.
Nej, hellre vill jag nu bliva kvävd, hellre dö än vara blott knotor!
Jag är led vid detta; aldrig kommer jag åter till liv.
Låt mig vara; mina dagar äro ju fåfänglighet.
Vad är då en människa, att du gör så stor sak av henne, aktar på henne så noga,
synar henne var morgon, prövar henne vart ögonblick?
Huru länge skall det dröja, innan du vänder din blick ifrån mig, lämnar mig i fred ett litet andetag?
Om jag än har syndar, vad skadar jag därmed dig, du människornas bespejare?
Varför har du satt mig till ett mål för dina angrepp och låtit mig bliva en börda för mig själv?
Varför vill du icke förlåta mig min överträdelse, icke tillgiva mig min missgärning?
Nu måste jag ju snart gå till vila i stoftet; om du söker efter mig, så är jag icke mer.
Därefter tog Bildad från Sua till orda och sade:
Huru länge vill du hålla på med sådant tal och låta din muns ord komma såsom en väldig storm?
Skulle väl Gud kunna kränka rätten?
Kan den Allsmäktige kränka rättfärdigheten?
Om dina barn hava syndat mot honom och han gav dem i sina överträdelsers våld,
så vet, att om du själv söker Gud och beder till den Allsmäktige om misskund,
då, om du är ren och rättsinnig, ja, då skall han vakna upp till din räddning och upprätta din boning, så att du bor där i rättfärdighet;
och så skall din första tid synas ringa, då nu din sista tid har blivit så stor.
Ty fråga framfarna släkten, och akta på vad fäderna hava utrönt
-- vi själva äro ju från i går och veta intet, en skugga äro våra dagar på jorden;
men de skola undervisa dig och säga dig det, ur sina hjärtan skola de hämta fram svar:
»Icke kan röret växa högt, där marken ej är sank, eller vassen skjuta i höjden, där vatten ej finnes?
Nej, bäst den står grön, ej mogen för skörd, måste den då vissna, före allt annat gräs.
Så går det alla som förgäta Gud; den gudlöses hopp måste varda om intet.
Ty hans tillförsikt visar sig bräcklig och hans förtröstan lik spindelns väv.
Han förlitar sig på sitt hus, men det har intet bestånd; han tryggar sig därvid, men det äger ingen fasthet.
Lik en frodig planta växer han i solens sken, ut över lustgården sträcka sig hans skott;
kring stenröset slingra sig hans rötter, mellan stenarna bryter han sig fram.
Men när så Gud rycker bort honom från hans plats, då förnekar den honom: 'Aldrig har jag sett dig.'
Ja, så går det med hans levnads fröjd, och ur mullen få andra växa upp.»
Se, Gud föraktar icke den som är ostrafflig, han håller ej heller de onda vid handen.
Så bida då, till dess han fyller din mun med löje och dina läppar med jubel.
De som hata dig varda då höljda med skam, och de ogudaktigas hyddor skola ej mer vara till.
Därefter tog Job till orda och sade:
Ja, förvisso vet jag att så är; huru skulle en människa kunna hava rätt mot Gud?
Vill han gå till rätta med henne, så kan hon ej svara honom på en sak bland tusen.
Han som är så vis i förstånd och så väldig i kraft, vem kan trotsa honom och dock slippa undan;
honom som oförtänkt flyttar bort berg och omstörtar dem i sin vrede;
honom som kommer jorden att vackla från sin plats, och dess pelare bäva därvid;
honom som befaller solen, så går hon icke upp, och som sätter stjärnorna under försegling;
honom som helt allena spänner ut himmelen och skrider fram över havets toppar;
honom som har gjort Karlavagnen och Orion, Sjustjärnorna och söderns Stjärngemak;
honom som gör stora och outrannsakliga ting och under, flera än någon kan räkna?
Se, han far förbi mig, innan jag hinner att se det, han drager framom mig, förrän jag bliver honom varse.
Se, han griper sitt rov; vem kan hindra honom?
Vem kan säga till honom: »Vad gör du?»
Gud, han ryggar icke sin vrede; för honom har Rahabs följe måst böja sig;
huru skulle jag då våga svara honom, välja ut ord till att tala med honom?
Nej, om jag än hade rätt, tordes jag dock ej svara; jag finge anropa min motpart om misskund.
Och om han än svarade mig på mitt rop, så kunde jag ej tro att han lyssnade till min röst.
Ty med storm hemsöker han mig och slår mig med sår på sår, utan sak.
Han unnar mig icke att hämta andan; nej, med bedrövelser mättar han mig.
Gäller det försteg i kraft: »Välan, jag är redo!», gäller det rätt: »Vem ställer mig till ansvar?»
Ja, hade jag än rätt, så dömde min mun mig skyldig; vore jag än ostrafflig, så läte han mig synas vrång.
Men ostrafflig är jag!
Jag aktar ej mitt liv, jag frågar icke efter, om jag får leva.
Det må gå som det vill, nu vare det sagt: han förgör den ostrafflige jämte den ogudaktige.
Om en landsplåga kommer med plötslig död, så bespottar han de oskyldigas förtvivlan.
Jorden är given i de ogudaktigas hand, och täckelse sätter han för dess domares ögon.
Är det ej han som gör det, vem är det då?
Min dagar hasta undan snabbare än någon löpare, de fly bort utan att hava sett någon lycka;
de ila åstad såsom en farkost av rör, såsom en örn, när han störtar sig ned på sitt byte.
Om jag än besluter att förgäta mitt bekymmer, att låta min sorgsenhet fara och göra mig glad,
Så måste jag dock bäva för alla mina kval; jag vet ju att du icke skall döma mig fri.
Nej, såsom skyldig måste jag stå där; varför skulle jag då göra mig fåfäng möda?
Om jag än tvår mig i snö och renar mina händer i lutsalt,
så skall du dock sänka mig ned i pölen, så att mina kläder måste vämjas vid mig.
Ty han är ej min like, så att jag vågar svara honom, ej en sådan, att vi kunna gå till doms med varandra;
ingen skiljeman finnes mellan oss, ingen som har myndighet över oss båda.
Må han blott vända av från mig sitt ris, och må fruktan för honom ej förskräcka mig;
då skall jag tala utan att rädas för honom, ty jag vet med min själv att jag icke är en sådan.
Min själ är led vid livet.
Jag vill giva fritt lopp åt min klagan, jag vill tala i min själs bedrövelse.
Jag vill säga till Gud: Döm mig icke skyldig; låt mig veta varför du söker sak mot mig.
Anstår det dig att öva våld, att förkasta dina händers verk, medan du låter ditt ljus lysa över de ogudaktigas rådslag?
Har du då ögon som en varelse av kött, eller ser du såsom människor se?
Är din ålder som en människas ålder, eller äro dina år såsom en mans tider,
eftersom du letar efter missgärning hos mig och söker att hos mig finna synd,
du som dock vet att jag icke är skyldig, och att ingen finnes, som kan rädda ur din hand?
Dina händer hava danat och gjort mig, helt och i allo; och nu fördärvar du mig!
Tänk på huru du formade mig såsom lera; och nu låter du mig åter varda till stoft!
Ja, du utgöt mig såsom mjölk, och såsom ostämne lät du mig stelna.
Med hud och kött beklädde du mig, av ben och senor vävde du mig samman.
Liv och nåd beskärde du mig, och genom din vård bevarades min ande.
Men därvid gömde du i ditt hjärta den tanken, jag vet att du hade detta i sinnet:
om jag syndade, skulle du vakta på mig och icke lämna min missgärning ostraffad.
Ve mig, om jag befunnes vara skyldig!
Men vore jag än oskyldig, så finge jag ej lyfta mitt huvud, jag skulle mättas av skam och skåda min ofärd.
Höjde jag det likväl, då skulle du såsom ett lejon jaga mig och alltjämt bevisa din undermakt på mig.
Nya vittnen mot mig skulle du då föra fram och alltmer låta mig känna din förtörnelse; med skaror efter skaror skulle du ansätta mig.
Varför lät du mig då komma ut ur modersskötet?
Jag borde hava förgåtts, innan något öga såg mig,
hava blivit såsom hade jag aldrig varit till; från moderlivet skulle jag hava förts till graven.
Kort är ju min tid; må han då låta mig vara, lämna mig i fred, så att jag får en flyktig glädje,
innan jag går hädan, för att aldrig komma åter, bort till mörkrets och dödsskuggans land,
till det land vars dunkel är såsom djupa vatten, dit där dödsskugga och förvirring råder, ja, där dagsljuset självt är såsom djupa vatten.
Därefter tog Sofar från Naama till orda och sade:
Skall sådant ordflöde bliva utan svar och en så stortalig man få rätt?
Skall ditt lösa tal nödga män till tystnad, så att du får bespotta, utan att någon kommer dig att blygas?
Och skall du så få säga: »Vad jag lär är rätt, och utan fläck har jag varit inför dina ögon»?
Nej, om allenast Gud ville tala och upplåta sina läppar till att svara dig,
om han ville uppenbara dig sin visdoms lönnligheter, huru han äger förstånd, ja, i dubbelt mått, då insåge du att Gud, dig till förmån, har lämnat åt glömskan en del av din missgärning.
Men kan väl du utrannsaka Guds djuphet eller fatta den Allsmäktiges fullkomlighet?
Hög såsom himmelen är den -- vad kan du göra? djupare än dödsriket -- vad kan du förstå?
Dess längd sträcker sig vidare än jorden, och i bredd överträffar den havet.
När han vill fara fram och spärra någon inne eller kalla någon till doms, vem kan då hindra honom?
Han är ju den som känner lögnens män, fördärv upptäcker han, utan att leta därefter.
Men lika lätt kan en dåraktig man få förstånd, som en vildåsnefåle kan födas till människa.
Om du nu rätt bereder ditt hjärta och uträcker dina händer till honom,
om du skaffar bort det fördärv som kan låda vid din hand och ej låter orättfärdighet bo i dina hyddor,
ja, då får du upplyfta ditt ansikte utan skam, du står fast och har intet att frukta.
Ja, då skall du förgäta din olycka, blott minnas den såsom vatten som har förrunnit.
Ditt liv skall då stråla klarare än middagens sken; och kommer mörker på, så är det som en gryning till morgon.
Du kan då vara trygg, ty du äger ett hopp; du spanar omkring dig och går sedan trygg till vila.
Ja, du får då ligga i ro, utan att någon förskräcker dig, och många skola söka din ynnest.
Men de ogudaktigas ögon skola försmäkta; ingen tillflykt skall mer finnas för dem, och deras hopp skall vara att få giva upp andan.
Därefter tog Job till orda och sade:
Ja, visst ären I det rätta folket, och med eder kommer visheten att dö ut!
Dock, jämväl jag har förstånd så gott som I, icke står jag tillbaka för eder; ty vem är den som ej begriper slikt?
Så måste jag då vara ett åtlöje för min vän, jag som fick svar, så snart jag ropade till Gud; man ler åt en som är rättfärdig och ostrafflig!
Ja, med förakt ses olyckan av den som står säker; förakt väntar dem vilkas fötter vackla.
Men förhärjares hyddor åtnjuta frid, och trygghet få sådana som trotsa Gud, de som hava sin gud i sin hand.
Men fråga du boskapen, den må undervisa dig, och fåglarna under himmelen, de må upplysa dig;
eller tala till jorden, hon må undervisa dig, fiskarna i havet må giva dig besked.
Vem kan icke lära genom allt detta att det är HERRENS hand som har gjort det?
I hans han är ju allt levandes själ och alla mänskliga varelsers anda.
Skall icke öra pröva orden, likasom munnen prövar matens smak?
Vishet tillkommer ju de gamle och förstånd dem som länge hava levat.
Hos Honom finnes vishet och makt, hos honom råd och förstånd.
Se, vad han river ned, det bygges ej upp; för den han spärrar inne kan ingen upplåta.
Han håller vattnen tillbaka -- se, se då bliver där torrt, han släpper dem lösa, då fördärva de landet.
Hos honom är kraft och klokhet, den förvillade och förvillaren äro båda i hans hand.
Rådsherrar utblottar han, han för dem i landsflykt, och domare gör han till dårar.
Han upplöser konungars välde och sätter fångbälte om deras höfter.
Präster utblottar han, han för dem i landsflykt, och de säkrast rotade kommer han på fall.
Välbetrodda män berövar han målet och avhänder de äldste deras insikt.
Han utgjuter förakt över furstar och lossar de starkes gördel.
Han blottar djupen, så att de ej höljas av mörker, dödsskuggan drager han fram i ljuset.
Han låter folkslag växa till -- och förgör dem; han utvidgar deras gränser, men för dem sedan bort.
Stamhövdingar i landet berövar han förståndet, han leder dem vilse i väglösa ödemarker.
De famla i mörkret och hava intet ljus, han kommer dem att ragla såsom druckna.
Ja, alltsammans har mitt öga sett, mitt öra har hört det och nogsamt givit akt.
Vad I veten, det vet också jag; icke står jag tillbaka för eder.
Men till den Allsmäktige vill jag nu tala, det lyster mig att gå till rätta med Gud.
Dock, I ären män som spinna ihop lögn, allasammans hopsätten I fåfängligt tal.
Om I ändå villen alldeles tiga!
Det kunde tillräknas eder som vishet.
Hören nu likväl mitt klagomål, och akten på mina läppars gensagor.
Viljen I försvara Gud med orättfärdigt tal och honom till förmån bruka oärligt tal?
Skolen I visa eder partiska för honom eller göra eder till sakförare för Gud?
Icke kan sådant ändas väl, när han håller räfst med eder?
Eller kunnen I gäckas med honom, såsom man kan gäckas med en människa?
Nej, förvisso skall han straffa eder, om I visen en hemlig partiskhet.
Sannerligen, hans majestät skall då förskräcka eder, och fruktan för honom skall falla över eder.
Edra tänkespråk skola då bliva visdomsord av aska, edra försvarsverk varda såsom vallar av ler.
Tigen nu för min, så skall jag tala, gånge så över mig vad det vara må.
Ja, huru det än går, vill jag fatta mitt kött mellan tänderna och taga min själ i min hand.
Må han dräpa mig, jag hoppas intet annat; min vandel vill jag ändå hålla fram inför honom.
Redan detta skall lända mig till frälsning, ty ingen gudlös dristar komma inför honom.
Hören, hören då mina ord, och låten min förklaring tränga in i edra öron.
Se, här lägger jag saken fram; jag vet att jag skall befinnas hava rätt.
Eller gives det någon som kan vederlägga mig?
Ja, då vill jag tiga -- och dö.
Allenast två ting må du ej göra mot mig, så behöver jag ej dölja mig inför ditt ansikte:
din hand må du ej låta komma mig när, och fruktan för dig må icke förskräcka mig.
Sedan må du åklaga, och jag vill svara, eller ock skall jag tala, och du må gendriva mig.
Huru är det alltså med mina missgärningar och synder?
Låt mig få veta min överträdelse och synd.
Varför döljer du ditt ansikte och aktar mig såsom din fiende?
Vill du skrämma ett löv som drives av vinden, vill du förfölja ett borttorkat strå?
Du skriver ju bedrövelser på min lott och giver mig till arvedel min ungdoms missgärningar;
du sätter mina fötter i stocken, du vaktar på alla vägar, för mina fotsulor märker du ut stegen.
Och detta mot en som täres bort lik murket trä, en som liknar en klädnad sönderfrätt av mal!
Människan, av kvinna född, lever en liten tid och mättas av oro;
lik ett blomster växer hon upp och vissnar bort, hon flyr undan såsom skuggan och har intet bestånd.
Och till att vakta på en sådan upplåter du dina ögon, ja, du drager mig till doms inför dig.
Som om en ren skulle kunna framgå av en oren!
Sådant kan ju aldrig ske.
Äro nu människans dagar oryggligt bestämda, hennes månaders antal fastställt av dig, har du utstakat en gräns som hon ej kan överskrida,
vänd då din blick ifrån henne och unna henne ro, låt henne njuta en dagakarls glädje av sin dag.
För ett träd finnes ju kvar något hopp; hugges det än ned, kan det åter skjuta skott, och telningar behöva ej fattas därpå.
Om än dess rot tynar hän i jorden och dess stubbe dör bort i mullen,
så kan det grönska upp genom vattnets ångor och skjuta grenar lik ett nyplantat träd.
Men om en man dör, så ligger han där slagen; om en människa har givit upp andan, var finnes hon då mer?
Såsom när vattnet har förrunnit ur en sjö, och såsom när en flod har sinat bort och uttorkat,
så ligger mannen där och står ej mer upp, han vaknar icke åter, så länge himmelen varar; aldrig väckes han upp ur sin sömn.
Ack, att du ville gömma mig i dödsriket, fördölja mig, till dess din vrede hade upphört, staka ut för mig en tidsgräns och sedan tänka på mig --
fastän ju ingen kan få liv, när han en gång är död!
Då skulle jag hålla min stridstid ut, ända till dess att min avlösning komme.
Du skulle då ropa på mig, och jag skulle svara dig; efter dina händers verk skulle du längta;
ja, du skulle då räkna mina steg, du skulle ej akta på min synd.
I en förseglad pung låge då min överträdelse, och du överskylde min missgärning.
Men såsom själva berget faller och förvittrar, och såsom klippan flyttas ifrån sin plats,
såsom stenar nötas sönder genom vattnet, och såsom mullen sköljes bort av dess flöden, så gör du ock människans hopp om intet.
Du slår henne ned för alltid, och hon far hädan; du förvandlar hennes ansikte och driver henne bort.
Om hennes barn komma till ära, så känner hon det icke; om de sjunka ned till ringhet, så aktar hon dock ej på dem.
Hennes kropp känner blott sin egen plåga, hennes själ blott den sorg hon själv får förnimma.
Därefter tog Elifas från Teman till orda och sade:
Skall en vis man tala så i vädret och fylla upp sitt bröst med östanvind?
Skall han försvara sin sak med haltlöst tal, med ord som ingenting bevisa?
Än mer, du gör gudsfruktan om intet och kommer med klagolåt inför Gud.
Ty din ondska lägger dig orden i munnen, och ditt behag står till illfundigt tal.
Så dömes du nu skyldig av din mun, ej av mig, dina egna läppar vittna emot dig.
Var du den första människa som föddes, och fick du liv, förrän höjderna funnos?
Blev du åhörare i Guds hemliga råd och fick så visheten i ditt våld?
Vad vet du då, som vi icke veta?
Vad förstår du, som ej är oss kunnigt?
Gråhårsman och åldring finnes också bland oss, ja, en som övergår din fader i ålder.
Försmår du den tröst som Gud har att bjuda, och det ord som i saktmod talas med dig?
Vart föres du hän av ditt sinne, och varför välva dina ögon så,
i det du vänder ditt raseri mot Gud och öser ut ord ur din mun?
Vad är en människa, att hon skulle vara ren?
Vad en av kvinna född, att han skulle vara rättfärdig?
Se, ej ens på sina heliga kan han förlita sig, och himlarna äro icke rena inför hans ögon;
huru mycket mindre då den som är ond och fördärvad, den man som läskar sig med orättfärdighet såsom med vatten!
Jag vill kungöra dig något, så hör nu mig; det som jag har skådat vill jag förtälja,
vad visa män hava gjort kunnigt, lagt fram såsom ett arv ifrån sina fäder,
ifrån dem som allena fingo landet till gåva, och bland vilka ingen främling ännu hade trängt in:
Den ogudaktige har ångest i alla sina dagar, under de år, helt få, som beskäras en våldsverkare.
Skräckröster ljuda i hans öron; när han är som tryggast, kommer förhärjaren över honom.
Han har intet hopp om räddning ur mörkret, ty svärdet lurar på honom.
Såsom flykting söker han sitt bröd: var är det?
Han förnimmer att mörkrets dag är för handen.
Ångest och trångmål förskräcka honom, han nedslås av dem såsom av en stridsrustad konung.
Ty mot Gud räckte han ut sin hand, och mot den Allsmäktige förhävde han sig;
han stormade mot honom med trotsig hals, med sina sköldars ryggar i sluten hop;
han höljde sitt ansikte med fetma och samlade hull på sin länd;
han bosatte sig i städer, dömda till förstöring, i hus som ej fingo bebos, ty till stenhopar voro de bestämda.
Därför bliver han ej rik, och hans gods består ej, hans skördar luta ej tunga mot jorden.
Han kan icke undslippa mörkret; hans telningar skola förtorka av hetta, och själv skall han förgås genom Guds muns anda.
I sin förvillelse må han ej lita på vad fåfängligt är, ty fåfänglighet måste bliva hans lön.
I förtid skall hans mått varda fyllt, och hans krona skall ej grönska mer.
Han bliver lik ett vinträd som i förtid mister sina druvor, lik ett olivträd som fäller sina blommor.
Ty den gudlöses hus förbliver ofruktsamt, såsom eld förtär hyddor där mutor tagas.
Man går havande med olycka och föder fördärv; den livsfrukt man alstrar är ett sviket hopp.
Därefter tog Job till orda och sade:
Över nog har jag fått höra av sådant; usla tröstare ären I alla.
Är det nu slut på detta tal i vädret, eller eggar dig ännu något till gensvar?
Jag kunde väl ock tala, jag såsom I; ja, jag ville att I voren i mitt ställe!
Då kunde jag hopsätta ord mot eder och skaka mot eder mitt huvud till hån.
Med munnen kunde jag då styrka eder och med läpparnas ömkan bereda eder lindring.
Om jag nu talar, så lindras därav ej min plåga; och tiger jag, icke släpper den mig ändå.
Nej, nu har all min kraft blivit tömd; du har ju förött hela mitt hus.
Och att du har hemsökt mig, det gäller såsom vittnesbörd; min sjukdom får träda upp och tala mot mig.
I vrede söndersliter och ansätter man mig, man biter sina tänder samman emot mig; ja, min ovän vässer mot mig sina blickar.
Man spärrar upp munnen mot mig, smädligt slår man mig på mina kinder; alla rota sig tillsammans emot mig.
Gud giver mig till pris åt orättfärdiga människor och kastar mig i de ogudaktigas händer.
Jag satt i god ro, då krossade han mig; han grep mig i nacken och slog mig i smulor.
Han satte mig upp till ett mål för sina skott;
från alla sidor träffa mig hans pilar, han genomborrar mina njurar utan förskoning, min galla gjuter han ut på jorden.
Han bryter ned mig med stöt på stöt, han stormar emot mig såsom en kämpe.
Säcktyg bär jag hopfäst över min hud, och i stoftet har jag måst sänka mitt horn,
Mitt anlete är glödande rött av gråt, och på mina ögonlock är dödsskugga lägrad.
Och detta, fastän våld ej finnes i mina händer, och fastän min bön är ren!
Du jord, överskyl icke mitt blod, och låt för mitt rop ingen vilostad finnas.
Se, redan nu har jag i himmelen mitt vittne, och i höjden den som skall tala för mig.
Mina vänner hava mig nu till sitt åtlöje, därför skådar mitt öga med tårar till Gud,
Ja, må han här skaffa rätt åt en man mot Gud och åt ett människobarn mot dess nästa.
Ty få äro de år som skola upprinna, innan jag vandrar den väg där jag ej mer kommer åter.
Min livskraft är förstörd, mina dagar slockna ut, bland gravar får jag min lott.
Ja, i sanning är jag omgiven av gäckeri, och avoghet får mitt öga ständigt skåda hos dessa!
Så ställ nu säkerhet och borgen för mig hos dig själv; vilken annan vill giva mig sitt handslag?
Dessas hjärtan har du ju tillslutit för förstånd, därför skall du icke låta dem triumfera.
Den som förråder sina vänner till plundring, på hans barn skola ögonen försmäkta.
Jag är satt till ett ordspråk bland folken; en man som man spottar i ansiktet är jag.
Därför är mitt öga skumt av grämelse, och mina lemmar äro såsom en skugga allasammans.
De redliga häpna över sådant, och den oskyldige uppröres av harm mot den gudlöse.
Men den rättfärdige håller fast vid sin väg, och den som har rena händer bemannar sig dess mer.
Ja, gärna mån I alla ansätta mig på nytt, jag lär ändå bland eder ej finna någon vis.
Mina dagar äro förlidna, sönderslitna äro mina planer, vad som var mitt hjärtas begär.
Men natten vill man göra till dag, ljuset skulle vara nära, nu då mörker bryter in.
Nej, huru jag än bidar, bliver dödsriket min boning, i mörkret skall jag bädda mitt läger;
till graven måste jag säga: »Du är min fader», till förruttnelsens maskar: »Min moder», »Min syster».
Vad bliver då av mitt hopp, ja, mitt hopp, vem får skåda det?
Till dödsrikets bommar far det ned, då jag nu själv går till vila i stoftet.
Därefter tog Bildad från Sua till orda och sade:
Huru länge skolen I gå på jakt efter ord?
Kommen till förstånd; sedan må vi talas vid.
Varför skola vi aktas såsom oskäliga djur, räknas i edra ögon såsom ett förstockat folk?
Du som i din vrede sliter sönder dig själv, menar du att dör din skull jorden skall bliva öde och klippan flyttas bort från sin plats?
Nej, den ogudaktiges ljus skall slockna ut, och lågan av hans eld icke giva något sken.
Ljuset skall förmörkas i hans hydda, och lampan slockna ut för honom.
Hans väldiga steg skola stäckas, hans egna rådslag bringa honom på fall.
Ty han rusar med sina fötter in i nätet, försåten lura, där han vandrar fram;
snaran griper honom om hälen, och gillret tager honom fatt;
garn till att fånga honom äro lagda på marken och snärjande band på hans stig.
Från alla sidor ängsla honom förskräckelser, de jaga honom, varhelst han går fram.
Olyckan vill uppsluka honom, och ofärd står redo, honom till fall.
Under hans hud frätas hans lemmar bort, ja, av dödens förstfödde bortfrätas hans lemmar.
Ur sin hydda, som han förtröstar på, ryckes han bort, och till förskräckelsernas konung vandrar han hän.
I hans hydda får främlingar bo, och svavel utströs över hans boning.
Nedantill förtorkas hans rötter, och ovantill vissnar hans krona bort.
Hans åminnelse förgås ifrån jorden, hans namn lever icke kvar i världen.
Från ljus stötes han ned i mörker och förjagas ifrån jordens krets.
Utan barn och avkomma bliver han i sitt folk, och ingen i hans boningar skall slippa undan.
Över hans ofärdsdag häpna västerns folk, och österns män gripas av rysning.
Ja, så sker det med den orättfärdiges hem, så går det dens hus, som ej vill veta av Gud.
Därefter tog Job till orda och sade:
Huru länge skolen I bedröva min själ och krossa mig sönder med edra ord?
Tio gånger haven I nu talat smädligt mot mig och kränkt mig utan all försyn.
Om så är, att jag verkligen har farit vilse, då är förvillelsen min egen sak.
Men viljen I ändå verkligen förhäva eder mot mig, och påstån I att smäleken har drabbat mig med skäl,
så veten fastmer att Gud har gjort mig orätt och att han har omsnärjt mig med sitt nät.
Se, jag klagar över våld, men får intet svar; jag ropar, men får icke rätt.
Min väg har han spärrat, så att jag ej kommer fram, och över mina stigar breder han mörker.
Min ära har han avklätt mig, och från mitt huvud har han tagit bort kronan.
Från alla sidor bryter han ned mig, så att jag förgås; han rycker upp mitt hopp, såsom vore det ett träd.
Sin vrede låter han brinna mot mig och aktar mig såsom sina ovänners like.
Hans skaror draga samlade fram och bereda sig väg till anfall mot mig; de lägra sig runt omkring min hydda.
Långt bort ifrån mig har han drivit mina fränder; mina bekanta äro idel främlingar mot mig.
Mina närmaste hava dragit sig undan, och mina förtrogna hava förgätit mig.
Mitt husfolk och mina tjänstekvinnor akta mig såsom främling; en främmande man har jag blivit i deras ögon.
Kallar jag på min tjänare, så svarar han icke; ödmjukt måste jag bönfalla hos honom.
Min andedräkt är vidrig för min hustru, jag väcker leda hos min moders barn.
Till och med de små barnen visa mig förakt; så snart jag står upp, tala de ohöviskt emot mig.
Ja, en styggelse är jag för alla dem jag umgicks med; de som voro mig kärast hava vänt sig emot mig.
Benen i min kropp tränga ut i hud och hull; knappt tandköttet har jag fått behålla kvar.
Haven misskund, haven misskund med mig, I mina vänner, då nu Guds hand så har hemsökt mig.
Varför skolen I förfölja mig, I såsom Gud, och aldrig bliva mätta av mitt kött?
Ack att mina ord skreves upp, ack att de bleve upptecknade i en bok,
ja, bleve med ett stift av järn och med bly för evig tid inpräglade i klippan!
Dock, jag vet att min förlossare lever, och att han till slut skall stå fram över stoftet.
Och sedan denna min sargade hud är borta, skall jag fri ifrån mitt kött få skåda Gud.
Ja, honom skall jag få skåda, mig till hjälp, för mina ögon skall jag se honom, ej såsom en främling; därefter trånar jag i mitt innersta.
Men när I tänken: »huru skola vi icke ansätta honom!» -- såsom vore skulden att finna hos mig --
då mån I taga eder till vara för svärdet, ty vreden hör till de synder som straffas med svärd; så mån I då besinna att en dom skall komma.
Därefter tog Sofar från Naama till orda och sade:
På sådant tal giva mina tankar mig ett svar, än mer, då jag nu är så upprörd i mitt inre.
Smädlig tillrättavisning måste jag höra, och man svarar mig med munväder på förståndigt tal.
Vet du då icke att så har varit från evig tid, från den stund då människor sattes på jorden:
att de ogudaktigas jubel varar helt kort och den gudlöses glädje ett ögonblick?
Om än hans förhävelse stiger upp till himmelen och hans huvud når intill molnen,
Så förgås han dock för alltid och aktas lik sin träck; de som sågo honom måste fråga: »Var är han?»
Lik en dröm flyger han bort, och ingen finner honom mer; han förjagas såsom en syn om natten.
Det öga som såg honom ser honom icke åter, och hans plats får ej skåda honom mer.
Hans barn måste gottgöra hans skulder till de arma, hans händer återbära hans vinning.
Bäst ungdomskraften fyller hans ben, skall den ligga i stoftet med honom.
Om än ondskan smakar ljuvligt i hans mun, så att han gömmer den under sin tunga,
är rädd om den och ej vill gå miste därom, utan håller den förvarad inom sin gom,
så förvandlas denna kost i hans inre, bliver huggormsetter i hans liv.
Den rikedom han har slukat måste han utspy; av Gud drives den ut ur hans buk.
Ja, huggormsgift kommer han att dricka, av etterormens tunga bliver han dräpt.
Ingen bäck får vederkvicka hans syn, ingen ström med flöden av honung och gräddmjölk.
Sitt fördärv måste han återbära, han får ej njuta därav; hans fröjd svarar ej mot den rikedom han har vunnit.
Ty mot de arma övade han våld och lät dem ligga där; han rev till sig hus som han ej kan hålla vid makt.
Han visste ej av någon ro för sin buk, men han skall icke rädda sig med sina skatter.
Intet slapp undan hans glupskhet, därför äger och hans lycka intet bestånd.
Mitt i hans överflöd påkommer honom nöd, och envar eländig vänder då mot honom sin hand.
Ja, så måste ske, för att hans buk må bliva fylld; sin vredes glöd skall Gud sända över honom och låta den tränga såsom ett regn in i hans kropp.
Om han flyr undan för vapen av järn, så genomborras han av kopparbågens skott.
När han då drager i pilen och den kommer ut ur hans rygg, när den ljungande udden kommer fram ur hans galla, då falla dödsfasorna över honom.
Idel mörker är förvarat åt hans skatter; till mat gives honom eld som brinner utan pust, den förtär vad som är kvar i hans hydda.
Himmelen lägger hans missgärning i dagen, och jorden reser sig upp emot honom.
Vad som har samlats i hans hus far åter sin kos, likt förrinnande vatten, på vredens dag.
Sådan lott får en ogudaktig människa av Gud, sådan arvedel har av Gud blivit bestämd åt henne.
Därefter tog Job till orda och sade:
Hören åtminstone på mina ord; låten det vara den tröst som I given mig.
Haven fördrag med mig, så att jag får tala; sedan jag har talat, må du bespotta.
Är då min klagan, såsom när människor eljest klaga?
Eller huru skulle jag kunna vara annat än otålig?
Akten på mig, så skolen I häpna och nödgas lägga handen på munnen.
Ja, när jag tänker därpå, då förskräckes jag själv, och förfäran griper mitt kött.
Varför få de ogudaktiga leva, ja, med åldern växa till i rikedom?
De se sina barn leva kvar hos sig, och sin avkomma hava de inför sina ögon.
Deras hus stå trygga, ej hemsökta av förskräckelse; Gud låter sitt ris icke komma vid dem.
När deras boskap parar sig, är det icke förgäves; lätt kalva deras kor, och icke i otid.
Sina barn släppa de ut såsom en hjord, deras piltar hoppa lustigt omkring.
De stämma upp med pukor och harpor, och glädja sig vid pipors ljud.
De förnöta sina dagar i lust, och ned till dödsriket fara de i frid.
Och de sade dock till Gud: »Vik ifrån oss, dina vägar vilja vi icke veta av.
Vad är den Allsmäktige, att vi skulle tjäna honom? och vad skulle det hjälpa oss att åkalla honom?»
Det är sant, i deras egen hand står ej deras lycka, och de ogudaktigas rådslag vare fjärran ifrån mig!
Men huru ofta utslocknar väl de ogudaktigas lampa, huru ofta händer det att ofärd kommer över dem, och att han tillskiftar dem lotter i vrede?
De borde ju bliva såsom halm för vinden, lika agnar som stormen rycker bort.
»Gud spar åt hans barn att lida för hans ondska.»
Ja, men honom själv borde han vedergälla, så att han finge känna det.
Med egna ögon borde han se sitt fall, och av den Allsmäktiges vrede borde han få dricka.
Ty vad frågar han efter sitt hus, när han själv är borta, när hans månaders antal har nått sin ände?
»Skall man då lära Gud förstånd, honom som dömer över de högsta?»
Ja, den ene får dö i sin välmaktstid, där han sitter i allsköns frid och ro;
hans stävor hava fått stå fulla med mjölk, och märgen i hans ben har bevarat sin saft.
Den andre måste dö med bedrövad själ, och aldrig fick han njuta av någon lycka.
Tillsammans ligga de så i stoftet, och förruttnelsens maskar övertäcka dem.
Se, jag känner väl edra tankar och de funder med vilka I viljen nedslå mig.
I spörjen ju: »Vad har blivit av de höga herrarnas hus, av hyddorna när de ogudaktiga bodde?»
Haven I då ej frågat dem som vida foro, och akten I ej på deras vittnesbörd:
att den onde bliver sparad på ofärdens dag och bärgad undan på vredens dag?
Vem vågar ens förehålla en sådan hans väg?
Vem vedergäller honom, vad han än må göra?
Och när han har blivit bortförd till graven, så vakar man sedan där vid kullen.
Ljuvligt får han vilja under dalens torvor.
I hans spår drager hela världen fram; före honom har och otaliga gått.
Huru kunnen I då bjuda mig så fåfänglig tröst?
Av edra svar står allenast trolösheten kvar.
Därefter tog Elifas från Teman till orda och sade:
Kan en man bereda Gud något gagn, så att det länder honom till gagn, om någon är förståndig?
Har den Allsmäktige någon båtnad av att du är rättfärdig, eller någon vinning av att du vandrar ostraffligt?
Är det för din gudsfruktans skull som han straffar dig, och som han går med dig till doms?
Har då icke din ondska varit stor, och voro ej dina missgärningar utan ände?
Jo, du tog pant av din broder utan sak, du plundrade de utblottade på deras kläder.
Åt den försmäktande gav du intet vatten att dricka, och den hungrige nekade du bröd.
För den väldige ville du upplåta landet, och den myndige skulle få bo däri,
men änkor lät du gå med tomma händer, och de faderlösas armar blevo krossade.
Därför omgives du nu av snaror och förfäras av plötslig skräck.
ja, av ett mörker där du intet ser, och av vattenflöden som övertäcka dig.
I himmelens höjde är det ju Gud som har sin boning, och du ser stjärnorna däruppe, huru högt de sitta;
därför tänker du: »Vad kan Gud veta?
Skulle han kunna döma, han som bor bortom töcknet?
Molnen äro ju ett täckelse, så att han intet ser; och på himlarunden är det han har sin gång.»
Vill du då hålla dig på forntidens väg, där fördärvets män gingo fram,
de män som bortrycktes, innan deras tid var ute, och såsom en ström flöt deras grundval bort,
de män som sade till Gud: »Vik ifrån oss», ty vad skulle den Allsmäktige kunna göra dem?
Det var ju dock han som uppfyllde deras hus med sitt goda.
De ogudaktigas rådslag vare fjärran ifrån mig!
De rättfärdiga skola se det och glädja sig, och den oskyldige skall få bespotta dem:
»Ja, nu äro förvisso våra motståndare utrotade, och deras överflöd har elden förtärt.»
Men sök nu förlikning och frid med honom; därigenom skall lycka falla dig till.
Tag emot undervisning av hans mun, och förvara hans ord i ditt hjärta.
Om du omvänder dig till den Allsmäktige, så bliver du upprättad; men orättfärdighet må du skaffa bort ur din hydda.
Ja kasta din gyllene skatt i stoftet och Ofirs-guldet ibland bäckens stenar,
så bliver den Allsmäktige din gyllene skatt, det ädlaste silver varder han för dig.
Ja, då skall du hava din lust i den Allsmäktige och kunna upplyfta ditt ansikte till Gud.
När du då beder till honom, skall han höra dig, och de löften du gör skall du få infria.
Allt vad du besluter skall då lyckas för dig, och ljus skall skina på dina vägar.
Om de leda mot djupet och du då beder: »Uppåt!», så frälsar han mannen som har ödmjukat sig.
Ja han räddar och den som ej är fri ifrån skuld; genom dina händers renhet räddas en sådan.
Därefter tog Job till orda och sade:
Också i dag vill min klaga göra uppror.
Min hand kännes matt för min suckans skull.
Om jag blott visste huru jag skulle finna honom, huru jag kunde komma dit där han bor!
Jag skulle då lägga fram för honom min sak och fylla min mun med bevis.
Jag ville väl höra vad han kunde svara mig, och förnimma vad han skulle säga till mig.
Icke med övermakt finge han bekämpa mig, nej, han borde allenast lyssna till mig.
Då skulle hans motpart stå här såsom en redlig man, ja, då skulle jag för alltid komma undan min domare.
Men går jag mot öster, så är han icke där; går jag mot väster, så varsnar jag honom ej;
har han något att skaffa i norr, jag skådar honom icke; döljer han sig i söder, jag ser honom ej heller där.
Han vet ju vilken väg jag har vandrat; han har prövat mig, och jag har befunnits lik guld.
Vid hans spår har min for hållit fast, hans väg har jag följt, utan att vika av.
Från hans läppars bud har jag icke gjort något avsteg; mer än egna rådslut har jag aktat hans muns tal.
Men hans vilja är orygglig; vem kan hindra honom?
Vad honom lyster, det gör han ock.
Ja, han giver mig fullt upp min beskärda del, och mycket av samma slag har han ännu i förvar.
Därför gripes jag av förskräckelse för hans ansikte; när jag betänker det, fruktar jag för honom.
Det är Gud som har gjort mitt hjärta försagt, den Allsmäktige är det som har vållat min förskräckelse,
ty jag fick icke förgås, innan mörkret kom, dödsnatten undanhöll han mig.
Varför har den Allsmäktige inga räfstetider i förvar? varför få hans vänner ej skåda hans hämndedagar?
Se, råmärken flyttar man undan, rövade hjordar driver man i bet;
de faderlösas åsna för man bort och tager änkans ko i pant.
Man tränger de fattiga undan från vägen, de betryckta i landet måste gömma sig med varandra.
Ja, såsom vildåsnor måste de leva i öknen; dit gå de och möda sig och söka något till täring; hedmarken är det bröd de hava åt sina barn.
På fältet få de till skörd vad boskap plägar äta, de hämta upp det sista i den ogudaktiges vingård.
Nakna ligga de om natten, berövade sina kläder; de hava intet att skyla sig med i kölden.
Av störtskurar från bergen genomdränkas de; de famna klippan, ty de äga ej annan tillflykt.
Den faderlöse slites från sin moders bröst, och den betryckte drabbas av utpantning.
Nakna måste de gå omkring, berövade sina kläder, hungrande nödgas de bära på kärvar.
Inom sina förtryckares murar måste de bereda olja, de få trampa vinpressar och därvid lida törst.
Utstötta ur människors samfund jämra de sig, ja, från dödsslagnas själar uppstiger ett rop.
Men Gud aktar ej på vad förvänt som sker.
Andra hava blivit fiender till ljuset; de känna icke dess vägar och hålla sig ej på dess stigar.
Vid dagningen står mördaren upp för att dräpa den betryckte och fattige; och om natten gör han sig till tjuvars like.
Äktenskapsbrytarens öga spejar efter skymningen, han tänker: »Intet öga får känna igen mig», och sätter så ett täckelse framför sitt ansikte.
När det är mörkt, bryta sådana sig in i husen, men under dagen stänga de sig inne; ljuset vilja de icke veta av.
Ty det svarta mörkret räknas av dem alla såsom morgon, med mörkrets förskräckelser äro de ju förtrogna.
»Men hastigt», menen I, »ryckes en sådan bort av strömmen, förbannad bliver hans del i landet; till vingårdarna får han ej mer styra sina steg.
Såsom snövatten förtäres av torka och hetta, så förtär dödsriket den som har syndat.
Hans moders liv förgäter honom, maskar frossa på honom, ingen finnes, som bevarar hans minne; såsom ett träd brytes orättfärdigheten av.
Så går det, när någon plundrar den ofruktsamma, som intet föder, och när någon icke gör gott mot änkan.»
Ja, men han uppehåller ock våldsmännen genom sin kraft, de få stå upp, när de redan hade förlorat hoppet om livet;
han giver dem trygghet, så att de få vila, och hans ögon vaka över deras vägar.
När de hava stigit till sin höjd, beskäres dem en snar hädanfärd, de sjunka då ned och dö som alla andra; likasom axens toppar vissna de bort.
Är det ej så, vem vill då vederlägga mig, vem kan göra mina ord om intet?
Därefter tog Bildad från Sua till orda och sade:
Hos honom är väldighet och förskräckande makt, hos honom, som skapar frid i sina himlars höjd.
Vem finnes, som förmår räkna hans skaror?
Och vem överstrålas ej av hans ljus?
Huru skulle då en människa kunna hava rätt mot Gud eller en av kvinna född kunna befinnas ren?
Se, ej ens månen skiner nog klart, ej ens stjärnorna äro rena i hans ögon;
huru mycket mindre då människan, det krypet, människobarnet, den masken!
Därefter tog Job till orda och sade:
Vilken hjälp har du ej skänkt den vanmäktige, huru har du ej stärkt den maktlöses arm!
Vilka råd har du ej givit den ovise, och vilket överflöd av klokhet har du ej lagt i dagen!
Vem gav dig kraft att tala sådana ord, och vems ande var det som kom till orda ur dig?
Dödsrikets skuggor gripas av ångest, djupets vatten och de som bo däri.
Dödsriket ligger blottat för honom, och avgrunden har intet täckelse.
Han spänner ut nordanrymden över det tomma och hänger upp jorden på intet.
Han samlar vatten i sina moln såsom i ett knyte, och skyarna brista icke under bördan.
Han gömmer sin tron för vår åsyn, han omhöljer den med sina skyar.
En rundel har han välvt såsom gräns för vattnen, där varest ljus ändas i mörker.
Himmelens pelare skälva, de gripas av förfäran vid hans näpst.
Med sin kraft förskräckte han havet, och genom sitt förstånd sönderkrossade han Rahab.
Blott han andades, blev himmelen klar; hans hand genomborrade den snabba ormen.
Se, detta är allenast utkanterna av hans verk; en sakta viskning är allt vad vi förnimma därom.
Hans allmakts dunder, vem skulle kunna fatta det?
Åter hov Job upp sin röst och kvad:
Så sant Gud lever, han som har förhållit mig min rätt, den Allsmäktige, som har vållat min själs bedrövelse:
aldrig, så länge ännu min ande är i mig och Guds livsfläkt är kvar i min näsa,
aldrig skola mina läppar tala vad orättfärdigt är, och min tunga bära fram oärligt tal.
Bort det, att jag skulle giva eder rätt!
Intill min död låter jag min ostrafflighet ej tagas ifrån mig.
Vid min rättfärdighet håller jag fast och släpper den icke, mitt hjärta förebrår mig ej för någon av mina dagar.
Nej, såsom ogudaktig må min fiende stå där och min motståndare såsom orättfärdig.
Ty vad hopp har den gudlöse när hans liv avskäres, när hans själ ryckes bort av Gud?
Månne Gud skall höra hans rop, när nöden kommer över honom?
Eller kan en sådan hava sin lust i den Allsmäktige, kan han åkalla Gud alltid?
Jag vill undervisa eder om huru Gud går till väga; huru den Allsmäktige tänker, vill jag icke fördölja.
Dock, I haven ju själva allasammans skådat det; huru kunnen I då hängiva eder åt så fåfängliga tankar?
Hören vad den ogudaktiges lott bliver hos Gud, vilken arvedel våldsverkaren får av den Allsmäktige:
Om hans barn bliva många, så är vinningen svärdets; hans avkomlingar få ej bröd att mätta sig med.
De som slippa undan läggas i graven genom pest, och hans änkor kunna icke hålla sin klagogråt.
Om han ock hopar silver såsom stoft och lägger kläder på hög såsom lera,
så är det den rättfärdige som får kläda sig i vad han lägger på hög, och den skuldlöse kommer att utskifta silvret.
Det hus han bygger bliver så förgängligt som malen, det skall likna skjulet som vaktaren gör sig.
Rik lägger han sig och menar att intet skall tagas bort; men när han öppnar sina ögon, är ingenting kvar.
Såsom vattenfloder taga förskräckelser honom fatt, om natten rövas han bort av stormen.
Östanvinden griper honom, så att han far sin kos, den rycker honom undan från hans plats.
Utan förskoning skjuter Gud sina pilar mot honom; för hans hand måste han flykta med hast.
Då slår man ihop händerna, honom till hån; man visslar åt honom på platsen där han var.
Silvret har ju sin gruva, sin fyndort har guldet, som man renar;
järn hämtas upp ur jorden, och stenar smältas till koppar.
Man sätter då gränser för mörkret, och rannsakar ned till yttersta djupet,
Där spränger man schakt långt under markens bebyggare, där färdas man förgäten djupt under vandrarens fot, där hänger man svävande, fjärran ifrån människor.
Ovan ur jorden uppväxer bröd, men därnere omvälves den såsom av eld.
Där, bland dess stenar, har safiren sitt fäste, guldmalm hämtar man ock där.
Stigen ditned är ej känd av örnen, och falkens öga har ej utspanat den;
den har ej blivit trampad av stolta vilddjur, intet lejon har gått därfram.
Ja, där bär man hand på hårda stenen; bergen omvälvas ända ifrån rötterna.
In i klipporna bryter man sig gångar, där ögat får se allt vad härligt är.
Vattenådror täppas till och hindras att gråta.
Så dragas dolda skatter fram i ljuset.
Men visheten, var finnes hon, och var har förståndet sin boning?
Priset för henne känner ingen människa; hon står ej att finna i de levandes land.
Djupet säger: »Hon är icke här», och havet säger: »Hos mig är hon icke.»
Hon köper icke för ädlaste metall, med silver gäldas ej hennes värde.
Hon väges icke upp med guld från Ofir, ej med dyrbar onyx och safir.
Guld och glas kunna ej liknas vid henne; hon får ej i byte mot gyllene klenoder.
Koraller och kristall må icke ens nämnas; svårare är förvärva vishet än pärlor.
Etiopisk topas kan ej liknas vid henne; hon väges icke upp med renaste guld.
Ja, visheten, varifrån kommer väl hon, och var har förståndet sin boning?
Förborgad är hon för alla levandes ögon, för himmelens fåglar är hon fördold;
avgrunden och döden giva till känna; »Blott hörsägner om henne förnummo våra öron.»
Gud, han är den som känner vägen till henne, han är den som vet var hon har sin boning.
Ty han förmår skåda till jordens ändar, allt vad som finnes under himmelen ser han.
När han mätte ut åt vinden dess styrka och avvägde vattnen efter mått,
när han stadgade en lag för regnet och en väg för tordönets stråle,
då såg han och uppenbarade henne, då lät han henne stå fram, då utforskade han henne.
Och till människorna sade han så: »Se Herrens fruktan, det är vishet, och att fly det onda är förstånd.»
Åter hov Job upp sin röst och kvad:
Ack att jag vore såsom i forna månader, såsom i de dagar då Gud gav mig sitt beskydd,
då hans lykta sken över mitt huvud och jag vid hans ljus gick fram genom mörkret!
Ja, vore jag såsom i min mognads dagar, då Guds huldhet vilade över min hydda,
då ännu den Allsmäktige var med mig och mina barn stodo runt omkring mig,
då mina fötter badade i gräddmjölk och klippan invid mig göt ut bäckar av olja!
När jag då gick upp till porten i staden och intog mitt säte på torget,
då drogo de unga sig undan vid min åsyn, de gamla reste sig upp och blevo stående.
Då höllo hövdingar tillbaka sina ord och lade handen på munnen;
furstarnas röst ljöd då dämpad, och deras tunga lådde vid gommen.
Ja, vart öra som hörde prisade mig då säll, och vart öga som såg bar vittnesbörd om mig;
ty jag räddade den betryckte som ropade, och den faderlöse, den som ingen hjälpare hade.
Den olyckliges välsignelse kom då över mig, och änkans hjärta uppfyllde jag med jubel.
I rättfärdighet klädde jag mig, och den var såsom min klädnad; rättvisa bar jag såsom mantel och huvudbindel.
Ögon blev jag då åt den blinde, och fötter var jag åt den halte.
Jag var då en fader för de fattiga, och den okändes sak redde jag ut.
Jag krossade den orättfärdiges käkar och ryckte rovet undan hans tänder.
Jag tänkte då: »I mitt näste skall jag få dö, mina dagar skola bliva många såsom sanden.
Min rot ligger ju öppen för vatten, och i min krona faller nattens dagg.
Min ära bliver ständigt ny, och min båge föryngras i min hand.»
Ja, på mig hörde man då och väntade, man lyssnade under tystnad på mitt råd.
Sedan jag hade talat, talade ingen annan; såsom ett vederkvickande flöde kommo mina ord över dem.
De väntade på mig såsom på regn, de spärrade upp sina munnar såsom efter vårregn.
När de misströstade, log jag emot dem, och mitt ansiktes klarhet kunde de icke förmörka.
Täcktes jag besöka dem, så måste jag sitta främst; jag tronade då såsom en konung i sin skara, lik en man som har tröst för de sörjande.
Och nu le de åt mig, människor som äro yngre till åren än jag, män vilkas fäder jag aktade ringa, ja, ej ens hade velat sätta bland mina vallhundar.
Vad skulle de också kunna gagna mig med sin hjälp, dessa människor som sakna all manlig kraft?
Utmärglade äro de ju av brist och svält; de gnaga sin föda av torra öknen, som redan i förväg är öde och ödslig.
Saltörter plocka de där bland snåren, och ginströtter är vad de hava till mat.
Ur människors samkväm drives de ut, man ropar efter dem såsom efter tjuvar.
I gruvliga klyftor måste de bo, i hålor under jorden och i bergens skrevor.
Bland snåren häva de upp sitt tjut, under nässlor ligga de skockade,
en avföda av dårar och ärelöst folk, utjagade ur landet med hugg och slag.
Och för sådana har jag nu blivit en visa, de hava mig till ämne för sitt tal;
med avsky hålla de sig fjärran ifrån mig, de hava ej försyn för att spotta åt mig.
Nej, mig till plåga, lossa de alla band, alla tyglar kasta de av inför mig.
Invid min högra sida upphäver sig ynglet; mina fötter vilja de stöta undan.
De göra sig vägar som skola leda till min ofärd.
Stigen framför mig hava de rivit upp.
De göra sitt bästa till att fördärva mig, de som dock själva äro hjälplösa.
Såsom genom en bred rämna bryta de in; de vältra sig fram under murarnas brak.
Förskräckelser välvas ned över mig.
Såsom en storm bortrycka de min ära, och såsom ett moln har min välfärd farit bort.
Och nu utgjuter sig min själ inom mig, eländesdagar hålla mig fast.
Natten bortfräter benen i min kropp, och kvalen som gnaga mig veta ej av vila.
Genom övermäktig kraft har mitt kroppshölje blivit vanställt, såsom en livklädnad hänger det omkring mig.
I orenlighet har jag blivit nedstjälpt, och själv är jag nu lik stoft och aska.
Jag ropar till dig, men du svarar mig icke; jag står här, men de bespejar mig allenast.
Du förvandlas för mig till en grym fiende, med din starka hand ansätter du mig.
Du lyfter upp mig i stormvinden och för mig hän, och i bruset låter du mig försmälta av ångest.
Ja, jag förstår att du vill föra mig till döden, till den boning dit allt levande församlas.
Men skulle man vid sitt fall ej få sträcka ut handen, ej ropa efter hjälp, när ofärd har kommit?
Grät jag ej själv över den som hade hårda dagar, och ömkade sig min själ ej över den fattige?
Se, jag väntade mig lycka, men olycka kom; jag hoppades på ljus, men mörker kom.
Därför sjuder mitt innersta och får ingen ro, eländesdagar hava ju mött mig.
Med mörknad hud går jag, fastän ej bränd av solen; mitt i församlingen står jag upp och skriar.
En broder har jag blivit till schakalerna, och en frände är jag vorden till strutsarna.
Min hud har svartnat och lossnat från mitt kött, benen i min kropp äro förbrända av hetta.
I sorgelåt är mitt harpospel förbytt, mina pipors klang i högljudd gråt.
Ett förbund slöt jag med mina ögon: aldrig skulle jag skåda efter någon jungfru.
Vilken lott finge jag eljest av Gud i höjden, vilken arvedel av den Allsmäktige därovan?
Ofärd kommer ju över de orättfärdiga, och olycka drabbar ogärningsmän.
Ser icke han mina vägar, räknar han ej alla mina steg?
Har jag väl umgåtts med lögn, och har min fot varit snar till svek?
Nej, må jag vägas på en riktig våg, så skall Gud förnimma min ostrafflighet.
Hava mina steg vikit av ifrån vägen, har mitt hjärta följt efter mina ögon, eller låder vid min händer en fläck?
Då må en annan äta var jag har sått, och vad jag har planterat må ryckas upp med roten.
Har mitt hjärta låtit dåra sig av någon kvinna, så att jag har stått på lur vid min nästas dörr?
Då må min hustru mala mjöl åt en annan, och främmande män må då famntaga henne.
Ja, sådant hade varit en skändlighet, en straffbar missgärning hade det varit,
en eld som skulle förtära intill avgrunden och förhärja till roten all min gröda.
Har jag kränkt min tjänares eller tjänarinnas rätt, när de hade någon tvist med mig?
Vad skulle jag då göra, när Gud stode upp, och när han hölle räfst, vad kunde jag då svara honom?
Han som skapade mig skapade ju och dem i moderlivet, han, densamme, har berett dem i modersskötet.
Har jag vägrat de arma vad de begärde eller låtit änkans ögon försmäkta?
Har jag ätit mitt brödstycke allena, utan att den faderlöse och har fått äta därav?
Nej, från min ungdom fostrades han hos mig såsom hos en fader, och från min moders liv var jag änkors ledare.
Har jag kunnat se en olycklig gå utan kläder, se en fattig ej äga något att skyla sig med?
Måste ej fastmer hans länd välsigna mig, och fick han ej värma sig i ull av mina lamm?
Har jag lyft min hand mot den faderlöse, därför att jag såg mig hava medhåll i porten?
Då må min axel lossna från sitt fäste och min arm brytas av ifrån sin led.
Jag måste då frukta ofärd ifrån Gud och skulle stå maktlös inför hans majestät.
Har jag satt mitt hopp till guldet och kallat guldklimpen min förtröstan?
Var det min glädje att min rikedom blev så stor, och att min hand förvärvade så mycket?
Hände det, när jag såg solljuset, huru det sken, och månen, huru härligt den gick fram,
att mitt hjärta hemligen lät dåra sig, så att jag med handkyss gav dem min hyllning?
Nej, också det hade varit en straffbar missgärning; därmed hade jag ju förnekat Gud i höjden.
Har jag glatt mig åt min fiendes ofärd och fröjdats, när olycka träffade honom?
Nej, jag tillstadde ej min mun att synda så, ej att med förbannelse begära hans liv.
Och kan mitt husfolk icke bevittna att envar fick mätta sig av kött vid mitt bord?
Främlingen behövde ej stanna över natten på gatan, mina dörrar lät jag stå öppna utåt vägen.
Har jag på människovis skylt mina överträdelser och gömt min missgärning i min barm,
av fruktan för den stora hopen och av rädsla för stamfränders förakt, så att jag teg och ej gick utom min dörr?
Ack att någon funnes, som ville höra mig!
Jag har sagt mitt ord.
Den Allsmäktige må nu svara mig; ack att jag finge min vederparts motskrift!
Sannerligen, jag skulle då bära den högt på min skuldra, såsom en krona skulle jag fästa den på mig.
Jag ville då göra honom räkenskap för alla mina steg, lik en furste skulle jag då träda inför honom.
Har min mark höjt rop över mig, och hava dess fåror gråtit med varandra?
Har jag förtärt dess gröda obetald eller utpinat dess brukares liv?
Då må törne växa upp för vete, och ogräs i stället för korn.
Slut på Jobs tal.
De tre männen upphörde nu att svara Job, eftersom han höll sig själv för rättfärdig.
Då blev Elihu, Barakels son, från Bus, av Rams släkt, upptänd av vrede.
Mot Job upptändes han av vrede, därför att denne menade sig hava rätt mot Gud;
och mot hans tre vänner upptändes hans vrede, därför att de icke funno något svar varmed de kunde vederlägga Job.
Hittills hade Elihu dröjt att tala till Job, därför att de andra voro äldre till åren än han.
Men då nu Elihu såg att de tre männen icke mer hade något att svara, upptändes hans vrede.
Så tog då Elihu, Barakels son, från Bus, till orda och sade; Ung till åren är jag, I däremot ären gamla.
Därför höll jag mig tillbaka och var försagd och lade ej fram för eder min mening.
Jag tänkte: »Må åldern tala, och må årens mängd förkunna visdom.»
Dock, på anden i människorna kommer det an, den Allsmäktiges livsfläkt giver dem förstånd.
Icke de åldriga äro alltid visast, icke de äldsta förstå bäst vad rätt är.
Därför säger jag nu: Hör mig; jag vill lägga fram min mening, också jag.
Se, jag väntade på vad I skullen tala, jag lyssnade efter förstånd ifrån eder, efter skäl som I skullen draga fram.
Ja, noga aktade jag på eder.
Men se, ingen fanns, som vederlade Job, ingen bland eder, som kunde svara på hans ord.
Nu mån I icke säga: »Vi möttes av vishet; Gud, men ingen människa, kan nedslå denne.»
Skäl mot min mening har han icke lagt fram, ej heller skall jag bemöta honom med edra bevis.
Se, nu stå de bestörta och svara ej mer, målet i munnen hava de mist.
Och jag skulle vänta, då de nu intet kunna säga, då de stå där och ej mer hava något svar!
Nej, också jag vill svara i min ordning, jag vill lägga fram min mening, också jag.
Ty, fullt upp har jag av skäl, anden i mitt inre vill spränga mig sönder.
Ja, mitt inre är såsom instängt vin, likt en lägel med nytt vin är det nära att brista.
Så vill jag då tala och skaffa mig luft, jag vill upplåta mina läppar och svara.
Jag får ej hava anseende till personen, och jag skall ej till någon tala inställsamma ord.
Nej, jag förstår ej att tala inställsamma ord; huru lätt kunde ej eljest min skapare rycka mig bort!
Men hör nu, Job, mina ord, och lyssna till allt vad jag vill säga.
Se, jag upplåter nu mina läppar, min tunga tager till orda i min mun.
Ur ett redbart hjärta framgår mitt tal, och vad mina läppar förstå säga de ärligt ut.
Guds ande är det som har gjort mig, den Allsmäktiges fläkt beskär mig liv.
Om du förmår, så må du nu svara mig; red dig till strid mot mig, träd fram.
Se, jag är likställd med dig inför Gud, jag är danad av en nypa ler, också jag.
Ja, fruktan för mig behöver ej förskräcka dig, ej heller kan min myndighet trycka dig ned.
Men nu sade du så inför mina öron, så ljödo de ord jag hörde:
»Ren är jag och fri ifrån överträdelse, oskyldig är jag och utan missgärning;
men se, han finner på sak mot mig, han aktar mig såsom sin fiende.
Han sätter mina fötter i stocken, vaktar på alla mina vägar.»
Nej, häri har du orätt, svarar jag dig.
Gud är ju förmer än en människa.
Huru kan du gå till rätta med honom, såsom gåve han aldrig svar i sin sak?
Både på ett sätt och på två talar Gud, om man också ej aktar därpå.
I drömmen, i nattens syn, när sömnen har fallit tung över människorna och de vila i slummer på sitt läger,
då öppnar han människornas öron och sätter inseglet på sina varningar till dem,
när han vill avvända någon från en ogärning eller hålla högmodet borta ifrån en människa.
Så bevarar han hennes själ från graven och hennes liv ifrån att förgås genom vapen.
Hon bliver ock agad genom plågor på sitt läger och genom ständig oro, allt intill benen.
Hennes sinne får leda vid maten, och hennes själ vid den föda hon älskade.
Hennes hull förtvinar, till dess intet är att se, ja, hennes ben täras bort intill osynlighet.
Så nalkas hennes själ till graven och hennes liv hän till dödens makter.
Men om en ängel då finnes, som vakar över henne, en medlare, någon enda av de tusen, och denne får lära människan hennes plikt,
då förbarmar Gud sig över henne och säger; »Fräls henne, så att hon slipper fara ned i graven; lösepenningen har jag nu fått.»
Hennes kropp får då ny ungdomskraft, hon bliver åter såsom under sin styrkas dagar.
När hon då beder till Gud, är han henne nådig och låter henne se sitt ansikte med jubel; han giver så den mannen hans rättfärdighet åter.
Så får denne då sjunga inför människorna och säga: »Väl syndade jag, och väl kränkte jag rätten, dock vederfors mig ej vad jag hade förskyllt;
ty han förlossade min själ, så att den undslapp graven, och mitt liv får nu med lust skåda ljuset.»
Se, detta allt kommer Gud åstad, både två gånger och tre, för den mannen,
till att rädda hans själ från graven, så att han får njuta av de levandes ljus.
Akta nu härpå, du Job, och hör mig; tig, så att jag får tala.
Dock, har du något att säga, så svara mig; tala, ty gärna gåve jag dig rätt.
Varom icke, så är det du som må höra på mig; du må tiga, så att jag får lära dig vishet.
Och Elihu tog till orda och sade:
Hören, I vise, mina ord; I förståndige, lyssnen till mig.
Örat skall ju pröva orden, och munnen smaken hos det man vill äta.
Må vi nu utvälja åt oss vad rätt är, samfällt söka förstå vad gott är.
Se, Job har sagt: »Jag är oskyldig.
Gud har förhållit mig min rätt.
Fastän jag har rätt, måste jag stå såsom lögnare; dödsskjuten är jag, jag som intet har brutit.»
Var finnes en man som är såsom Job?
Han läskar sig med bespottelse såsom med vatten,
han gör sig till ogärningsmäns stallbroder och sällar sig till ogudaktiga människor.
Ty han säger: »Det gagnar en man till intet, om han håller sig väl med Gud.»
Hören mig därför, I förståndige män: Bort det, att Gud skulle begå någon orätt, att den Allsmäktige skulle göra vad orättfärdigt är!
Nej, han vedergäller var människa efter hennes gärningar och lönar envar såsom hans vandel har förtjänat.
Ty Gud gör i sanning intet som är orätt, den Allsmäktige kan icke kränka rätten.
Vem har bjudit honom att vårda sig om jorden, och vem lade på honom bördan av hela jordens krets?
Om han ville tänka allenast på sig själv och åter draga till sig sin anda och livsfläkt,
då skulle på en gång allt kött förgås, och människorna skulle vända åter till stoft.
Men märk nu väl och hör härpå, lyssna till vad mina ord förkunna.
Skulle den förmå regera, som hatade vad rätt är?
Eller fördömer du den som är den störste i rättfärdighet?
Får man då säga till en konung: »Du ogärningsman», eller till en furste: »Du ogudaktige»?
Gud har ju ej anseende till någon hövdings person, han aktar den rike ej för mer än den fattige, ty alla äro de hans händers verk.
I ett ögonblick omkomma de, mitt i natten: folkhopar gripas av bävan och förgås, de väldige ryckas bort, utan människohand.
Ty hans ögon vakta på var mans vägar, och alla deras steg, dem ser han.
Intet mörker finnes och ingen skugga så djup, att ogärningsmän kunna fördölja sig däri.
Ty länge behöver Gud ej vakta på en människa, innan hon måste stå till doms inför honom.
Han krossar de väldige utan rannsakning och låter så andra träda fram i deras ställe.
Ja, han märker väl vad de göra, han omstörtar dem om natten och låter dem förgås.
Såsom ogudaktiga tuktar han dem öppet, inför människors åsyn,
eftersom de veko av ifrån honom och ej aktade på alla hans vägar.
De bragte så den armes rop inför honom, och rop av betryckta fick han höra.
Vem vågar då fördöma, om han stillar larmet?
Ja, vem vill väl skåda honom, om han döljer sitt ansikte, för ett folk eller för en enskild man,
när han vill rycka makten ifrån gudlösa människor och hindra dem att bliva snaror för folket?
Kan man väl säga till Gud: »Jag måste lida, jag som ändå intet har förbrutit.
Visa mig du vad som går över mitt förstånd; om jag har gjort något orätt, vill jag då ej göra så mer.»
Skall då han, för ditt klanders skull, giva vedergällning såsom du vill?
Du själv, och icke jag, må döma därom; ja, tala du ut vad du menar.
Men kloka män skola säga så till mig, visa män, när de få höra mig:
»Job talar utan någon insikt, hans ord äro utan förstånd.»
Så må nu Job utstå prövningar allt framgent, då han vill försvara sig på ogärningsmäns sätt.
Till sin synd lägger han ju uppenbar ondska, oss till hån slår han ihop sina händer och talar stora ord mot Gud.
Och Elihu tog till orda och sade:
Menar du att sådant är riktigt?
Kan du påstå att du har rätt mot Gud,
du som frågar vad rättfärdighet gagnar dig, vad den båtar dig mer än synd?
Svar härpå vill jag giva dig, jag ock dina vänner med dig.
Skåda upp mot himmelen och se, betrakta skyarna, som gå där högt över dig.
Om du syndar, vad gör du väl honom därmed?
Och om dina överträdelser äro många, vad skadar du honom därmed?
Eller om du är rättfärdig, vad giver du honom, och vad undfår han av din hand?
Nej, för din like kunde din ogudaktighet något betyda och för en människoson din rättfärdighet.
Väl klagar man, när våldsgärningarna äro många, man ropar om hjälp mot de övermäktigas arm;
men ingen frågar: »Var är min Gud, min skapare, han som låter lovsånger ljuda mitt i natten,
han som giver oss insikt framför markens djur och vishet framför himmelens fåglar?»
Därför är det man får ropa utan svar om skydd mot de ondas övermod.
Se, på fåfängliga böner hör icke Gud, den Allsmäktige aktar icke på slikt;
allra minst, när du påstår att du icke får skåda honom, att du måste vänta på honom, fastän saken är uppenbar.
Och nu menar du att hans vrede ej håller någon räfst, och att han föga bekymrar sig om människors övermod?
Ja, till fåfängligt tal spärrar Job upp sin mun, utan insikt talar han stora ord.
Vidare sade Elihu:
Bida ännu litet, så att jag får giva dig besked, ty ännu något har jag att säga till Guds försvar.
Min insikt vill jag hämta vida ifrån, och åt min skapare vill jag skaffa rätt.
Ja, förvisso skola mina ord icke vara lögn; en man med fullgod insikt har du framför dig.
Se, Gud är väldig, men han försmår dock ingen, han som är så väldig i sitt förstånds kraft.
Den ogudaktige låter han ej bliva vid liv, men åt de arma skaffar han rätt.
Han tager ej sina ögon från de rättfärdiga; de få trona i konungars krets, för alltid låter han dem sitta där i höghet.
Och om de läggas bundna i kedjor och fångas i eländets snaror,
så vill han därmed visa dem vad de hava gjort, och vilka överträdelser de hava begått i sitt högmod;
han vill då öppna deras öra för tuktan och mana dem att vända om ifrån fördärvet.
Om de då höra på honom och underkasta sig, så få de framleva sina dagar i lycka och sina år i ljuvlig ro.
Men höra de honom ej, så förgås de genom vapen och omkomma, när de minst tänka det.
Ja, de som med gudlöst hjärta hängiva sig åt vrede och icke anropa honom, när han lägger dem i band,
deras själ skall i deras ungdom ryckas bort av döden, och deras liv skall dela tempelbolares lott.
Genom lidandet vill han rädda den lidande, och genom betrycket vill han öppna hans öra.
Så sökte han ock draga dig ur nödens gap, ut på en rymlig plats, där intet trångmål rådde; och ditt bord skulle bliva fullsatt med feta rätter.
Men nu bär du till fullo ogudaktighetens dom; ja, dom och rättvisa hålla dig nu fast.
Ty vrede borde ej få uppegga dig under din tuktans tid, och huru svårt du än har måst plikta, borde du ej därav ledas vilse.
Huru kan han lära dig bedja, om icke genom nöd och genom allt som nu har prövat din kraft?
Du må ej längta så ivrigt efter natten, den natt då folken skola ryckas bort ifrån sin plats.
Tag dig till vara, så att du ej vänder dig till vad fördärvligt är; sådant behagar dig ju mer än att lida.
Se, Gud är upphöjd genom sin kraft.
Var finnes någon mästare som är honom lik?
Vem har föreskrivit honom hans väg, och vem kan säga: »Du gör vad orätt är?»
Tänk då på att upphöja hans gärningar, dem vilka människorna besjunga
och som de alla skåda med lust, de dödliga, om de än blott skönja dem i fjärran.
Ja, Gud är för hög för vårt förstånd, hans år äro flera än någon kan utrannsaka.
Se, vattnets droppar drager han uppåt, och de sila ned såsom regn, där hans dimma går fram;
skyarna gjuta dem ut såsom en ström, låta dem drypa ned över talrika människor.
Ja, kan någon fatta molnens utbredning, braket som utgår från hans hydda?
Se, sitt ljungeldsljus breder han ut över molnen, och själva havsgrunden höljer han in däri.
Ty så utför han sina domar över folken; så bereder han ock näring i rikligt mått.
I ljungeldsljus höljer han sina händer och sänder det ut mot dem som begynna strid.
Budskap om honom bär hans dunder; själva boskapen bebådar hans antåg.
Ja, vid sådant förskräckes mitt hjärta, bävande spritter det upp.
Hören, hören huru hans röst ljuder vred, hören dånet som går ut ur hans mun.
Han sänder det åstad, så långt himmelen når, och sina ljungeldar bort till jordens ändar.
Efteråt ryter så dånet, när han dundrar med sin väldiga röst; och på ljungeldarna spar han ej, då hans röst låter höra sig.
Ja, underbart dundrar Gud med sin röst, stora ting gör han, utöver vad vi förstå.
Se, åt snön giver han bud: »Fall ned till jorden», så ock åt regnskuren, åt sitt regnflödes mäktiga skur.
Därmed fjättrar han alla människors händer, så att envar som han har skapat kan lära därav.
Då draga sig vilddjuren in i sina gömslen, och i sina kulor lägga de sig till ro.
Från Stjärngemaket kommer då storm och köld genom nordanhimmelens stjärnor;
med sin andedräkt sänder Gud frost, och de vida vattnen betvingas.
Skyarna lastar han ock med väta och sprider omkring sina ljungeldsmoln.
De måste sväva än hit, än dit, alltefter hans rådslut och de uppdrag de få, vadhelst han ålägger dem på jordens krets.
Än är det som tuktoris, än med hjälp åt hans jord, än är det med nåd som han låter dem komma.
Lyssna då härtill, du Job; stanna och betänk Guds under.
Förstår du på vad sätt Gud styr deras gång och låter ljungeldarna lysa fram ur sina moln?
Förstår du lagen för skyarnas jämvikt, den Allvises underbara verk?
Förstår du huru kläderna bliva dig så heta, när han låter jorden domna under sunnanvinden?
Kan du välva molnhimmelen så som han, så fast som en spegel av gjuten metall?
Lär oss då vad vi skola säga till honom; för vårt mörkers skull hava vi intet att lägga fram.
Ej må det bebådas honom att jag vill tala.
Månne någon begär sitt eget fördärv?
Men synes icke redan skenet?
Strålande visar han sig ju mellan skyarna, där vinden har gått fram och sopat dem undan.
I guldglans kommer han från norden.
Ja, Gud är höljd i fruktansvärt majestät;
den Allsmäktige kunna vi icke fatta, honom som är så stor i kraft, honom som ej kränker rätten, ej strängaste rättfärdighet.
Fördenskull frukta människorna honom; men de självkloka -- dem alla aktar han ej på.
Och HERREN svarade Job ur stormvinden och sade:
Vem är du som stämplar vishet såsom mörker, i det att du talar så utan insikt?
Omgjorda nu såsom ej man dina länder; jag vill fråga dig, och du må giva mig besked.
Var var du, när jag lade jordens grund?
Säg det, om du har ett så stort förstånd.
Vem har fastställt hennes mått -- du vet ju det?
Och vem spände sitt mätsnöre ut över henne?
Var fingo hennes pelare sina fästen, och vem var det som lade hennes hörnsten,
medan morgonstjärnorna tillsammans jublade och alla Guds söner höjde glädjerop?
Och vem satte dörrar för havet, när det föddes och kom ut ur moderlivet,
när jag gav det moln till beklädnad och lät töcken bliva dess linda,
när jag åt det utstakade min gräns och satte bom och dörrar därför,
och sade: »Härintill skall du komma, men ej vidare, här skola dina stolta böljor lägga sig»?
Har du i din tid bjudit dagen att gry eller anvisat åt morgonrodnaden dess plats,
där den skulle fatta jorden i dess flikar, så att de ogudaktiga skakades bort därifrån?
Då ändrar den form såsom leran under signetet, och tingen stå fram såsom klädda i skrud;
då berövas de ogudaktiga sitt ljus, och den arm som lyftes för högt brytes sönder.
Har du stigit ned till havets källor och vandrat omkring på djupets botten?
Hava dödens portar avslöjat sig för dig, ja, såg du dödsskuggans portar?
Har du överskådat jordens vidder?
Om du känner allt detta, så låt höra.
Vet du vägen dit varest ljuset bor, eller platsen där mörkret har sin boning,
så att du kan hämta dem ut till deras gräns och finna stigarna som leda till deras hus?
Visst kan du det, ty så tidigt blev du ju född, så stort är ju dina dagars antal!
Har du varit framme vid snöns förrådshus?
Och haglets förrådshus, du såg väl dem
-- de förråd som jag har sparat till hemsökelsens tid, till stridens och drabbningens dag?
Vet du vägen dit varest ljuset delar sig, dit där stormen sprider sig ut över jorden?
Vem har åt regnflödet öppnat en ränna och banat en väg för tordönets stråle,
till att sända regn över länder där ingen bor, över öknar, där ingen människa finnes,
till att mätta ödsliga ödemarker och giva växt åt gräsets brodd?
Säg om regnet har någon fader, och vem han är, som födde daggens droppar?
Ur vilken moders liv är det isen gick fram, och vem är hon som födde himmelens rimfrost?
Se, vattnet tätnar och bliver likt sten, så ytan sluter sig samman över djupet.
Knyter du tillhopa Sjustjärnornas knippe?
Och förmår du att lossa Orions band?
Är det du som, när tid är, för himmelstecknen fram, och som leder Björninnan med hennes ungar?
Ja, förstår du himmelens lagar, och ordnar du dess välde över jorden?
Kan du upphöja din röst till molnen och förmå vattenflöden att övertäcka dig?
Kan du sända ljungeldar åstad, så att de gå, så att de svara dig: »Ja vi äro redo»?
Vem har lagt vishet i de mörka molnen, och vem gav förstånd åt järtecknen i luften?
Vem håller med sin vishet räkning på skyarna?
Och himmelens läglar, vem häller ut dem,
medan mullen smälter såsom malm och jordkokorna klibbas tillhopa?
Är det du som jagar upp rov åt lejoninnan och stillar de unga lejonens hunger,
när de trycka sig ned i sina kulor eller ligga på lur i snåret?
Vem är det som skaffar mat åt korpen, när hans ungar ropar till Gud, där de sväva omkring utan föda?
Vet du tiden för stengetterna att föda, vakar du över när hindarna bör kalva?
Räknar du månaderna som de skola gå dräktiga, ja, vet du tiden för dem att föda?
De böja sig ned, de avbörda sig sina foster, hastigt göra de sig fria ifrån födslovåndan.
Deras ungar frodas och växa till på marken, så springa de sin väg och vända ej tillbaka.
Vem har skänkt vildåsnan hennes frihet, vem har lossat den skyggas band?
Se, hedmarken gav jag henne till hem, och saltöknen blev hennes boning.
Hon ler åt larmet i staden, hon hör ingen pådrivares rop.
Vad hon spanar upp på berget har hon till bete, hon letar efter allt som är grönt.
Skall vildoxen finnas hågad att tjäna dig och att stanna över natten invid din krubba?
Kan du tvinga vildoxen att gå i fåran efter töm och förmå honom att i ditt spår harva markerna jämna?
Kan du lita på honom, då ju hans kraft är så stor, kan du betro åt honom ditt arbetes frukt?
Överlåter du åt honom att föra hem din säd och att hämta den tillhopa till din loge?
Strutshonans vingar flaxa med fröjd, men vad modersömhet visa väl hennes pennor, hennes fjädrar?
Åt jorden överlåter hon ju sina ägg och ruvar dem ovanpå sanden.
Hon bryr sig ej om att en fot kan krossa dem, att ett vilddjur kan trampa dem sönder.
Hård är hon mot sin avkomma, såsom vore den ej hennes; att hennes avel kan gå under, det bekymrar henne ej.
Ty Gud har gjort henne glömsk för vishet, han har ej tilldelat henne förstånd.
Men när det gäller, piskar hon sig själv upp till språng; då ler hon åt både häst och man.
Är det du som giver åt hästen hans styrka och kläder hans hals med brusande man?
Är det du som lär honom gräshoppans språng?
Hans stolta frustning, en förskräckelse är den!
Han skrapar marken och fröjdar sig i sin kraft och rusar så fram mot väpnade skaror.
Han ler åt fruktan och känner ej förfäran, han ryggar icke tillbaka för svärd.
Omkring honom ljuder ett rassel av koger, av ljungande spjut och lans.
Han skakas och rasar och uppslukar marken, han kan icke styra sig, när basunen har ljudit.
För var basunstöt frustar han: Huj!
Ännu i fjärran vädrar han striden, anförarnas rop och larmet av härskrin.
Är det ett verk av ditt förstånd, att falken svingar sig upp och breder ut sina vingar till flykt mot söder?
Eller är det på ditt bud som örnen stiger så högt och bygger sitt näste i höjden?
På klippan bor han, där har han sitt tillhåll, på klippans spets och på branta berget.
Därifrån spanar han efter sitt byte, långt bort i fjärran skådar hans ögon.
Hans ungar frossa på blod, och där slagna ligga, där finner man honom.
Så svarade nu HERREN Job och sade:
Vill du tvista med den Allsmäktige, du mästare?
Svara då, du som så klagar på Gud!
Job svarade HERREN och sade:
Nej, därtill är jag för ringa; vad skulle jag svara dig?
Jag måste lägga handen på munnen.
En gång har jag talat, och nu säger jag intet mer; ja, två gånger, men jag gör det icke åter.
Och HERREN talade till Job ur stormvinden och sade:
Omgjorda såsom en man dina länder; jag vill fråga dig, och du må giva mig besked.
Vill du göra min rätt om intet och döma mig skyldig, för att själv stå såsom rättfärdig?
Har du en sådan arm som Gud, och förmår du dundra med din röst såsom han?
Pryd dig då med ära och höghet, kläd dig i majestät och härlighet.
Gjut ut din vredes förgrymmelse, ödmjuka med en blick allt vad högt är.
Ja, kuva med en blick allt vad högt är, slå ned de ogudaktiga på stället.
Göm dem i stoftet allasammans, ja, fjättra deras ansikten i mörkret.
Då vill jag prisa dig, också jag, för segern som din högra hand har berett dig.
Se, Behemot, han är ju mitt verk såväl som du.
Han lever av gräs såsom en oxe.
Och se vilken kraft han äger i sina länder, vilken styrka han har i sin buks muskler.
Han bär sin svans så styv som en ceder, ett konstrikt flätverk äro senorna i hans lår.
Hans benpipor äro såsom rör av koppar, benen i hans kropp likna stänger av järn.
Förstlingen är han av vad Gud har gjort; hans skapare själv har givit honom hans skära.
Ty foder åt honom frambära bergen, där de vilda djuren alla hava sin lek.
Under lotusträd lägger han sig ned, i skygdet av rör och vass.
Lotusträd giva honom tak och skugga, pilträd hägna honom runt omkring.
Är floden än så våldsam, så ängslas han dock icke; han är trygg, om ock en Jordan bryter fram mot hans gap.
Vem kan fånga honom, när han är på sin vakt, vem borrar en snara genom hans nos?
Kan du draga upp Leviatan med krok och med en metrev betvinga hans tunga?
Kan du sätta en sävhank i hans nos eller borra en hake genom hans käft?
Menar du att han skall slösa på dig många böner eller tala till dig med mjuka ord?
Att han skall vilja sluta fördrag med dig, så att du finge honom till din träl för alltid?
Kan du hava honom till leksak såsom en fågel och sätta honom i band åt dina tärnor?
Pläga fiskarlag köpslå om honom och stycka ut hans kropp mellan krämare?
Kan du skjuta hans hud full med spjut och hans huvud med fiskharpuner?
Ja, försök att bära hand på honom du skall minnas den striden och skall ej föra så mer.
Nej, den sådant vågar, hans hopp bliver sviket, han fälles till marken redan vid hans åsyn.
Så oförvägen är ingen, att han törs reta denne.
Vem vågar då sätta sig upp mot mig själv?
Vem har först givit mig något, som jag alltså bör betala igen?
Mitt är ju allt vad som finnes under himmelen.
Jag vill ej höra upp att tala om hans lemmar, om huru väldig han är, och huru härligt han är danad.
Vem mäktar rycka av honom hans pansar?
Vem vågar sig in mellan hans käkars par?
Hans gaps dörrar, vem vill öppna dem?
Runtom hans tänder bor ju förskräckelse.
Stolta sitta på honom sköldarnas rader; hopslutna äro de med fast försegling.
Tätt fogar sig den ena intill den andra, icke en vindfläkt tränger in mellan dem.
Var och en håller ihop med den nästa, de gripa in i varandra och skiljas ej åt.
När han fnyser, strålar det av ljus; hans blickar äro såsom morgonrodnadens ögonbryn.
Bloss fara ut ur hans gap, eldgnistor springa fram därur.
Från hans näsborrar utgår rök såsom ur en sjudande panna på bränslet.
Hans andedräkt framgnistrar eldkol, och lågor bryta fram ur hans gap.
På hans hals har kraften sin boning, och framför honom stapplar försagdhet.
Själva det veka på hans buk är ett stadigt fogverk, det sitter orubbligt, såsom gjutet på honom.
Hans hjärta är fast såsom sten, fast såsom bottenstenen i kvarnen.
När han reser sig, bäva hjältar, av ångest mista de all sans.
Angripes han med ett svärd, så håller det ej stånd, ej heller spjut eller pil eller pansar.
Han aktar järn såsom halm och koppar såsom murket trä.
Bågskott skrämma honom ej bort, slungstenar förvandlas för honom till strå;
ja, stridsklubbor aktar han såsom strå, han ler åt rasslet av lansar.
På sin buk bär han skarpa eggar, spår såsom av en tröskvagn ristar han i dyn.
Han gör djupet sjudande som en gryta, likt en salvokokares kittel förvandlar han vattnet.
Bakom honom strålar vägen av ljus, djupet synes bära silverhår.
Ja, på jorden finnes intet som är honom likt, otillgänglig för fruktan skapades han.
På allt vad högt är ser han med förakt, konung är han över alla stolta vilddjur.
Job svarade HERREN och sade:
Ja, jag vet att du förmår allt, och att intet som du besluter är dig för svårt.
Vem var då jag som i oförstånd gav vishet namn av mörker?
Jag ordade ju om vad jag icke begrep, om det som var mig för underbart och det jag ej kunde förstå.
Men hör nu, så vill jag tala; jag vill fråga dig, och du må giva mig besked.
Blott hörsägner hade jag förnummit om dig, men nu har jag fått se dig med egna ögon.
Därför tager jag det tillbaka och ångrar mig, i stoft och aska.
Sedan HERREN hade talat så till Job, sade han till Elifas från Teman: »Min vrede är upptänd mot dig och dina båda vänner, därför att I icke haven talat om mig vad rätt är, såsom min tjänare Job har gjort.
Så tagen eder nu sju tjurar och sju vädurar, och gån till min tjänare Job och offren dem såsom brännoffer för eder; ock låten min tjänare Job bedja för eder.
Till äventyrs skall jag då, av nåd mot honom, avstå från att göra något förskräckligt mot eder, till straff därför att I icke haven talat om mig vad rätt är, såsom min tjänare Job har gjort.»
Då gingo Elifas från Teman, Bildad från Sua och Sofar från Naaman åstad och gjorde såsom HERREN hade tillsagt dem; och HERREN tog nådigt emot Jobs bön.
Och då nu Job bad för sina vänner, upprättade HERREN åter honom själv; HERREN gav Job dubbelt igen mot vad han förut hade haft.
Och alla hans bröder och systrar och alla hans forna bekanta kommo till honom och höllo måltid med honom i hans hus, och ömkade honom för alla de olyckor som HERREN hade låtit komma över honom.
Och de gåvo honom vardera en kesita och en guldring.
Och HERREN välsignade slutet av Jobs levnad ännu mer än begynnelsen, så att han fick fjorton tusen får, sex tusen kameler, ett tusen par oxar och ett tusen åsninnor.
Och han fick sju söner och tre döttrar.
Den första dottern kallade han Jemima, den andra Kesia och den tredje Keren-Happuk.
Och så sköna kvinnor som Jobs döttrar funnos icke i hela landet; och deras fader gav dem arvedel bland deras bröder.
Och Job levde därefter ett hundra fyrtio år, och fick se sina barn och barnbarn i fyra led.
Sedan dog Job, gammal och mätt på att leva.
Säll är den man som icke vandrar i de ogudaktigas råd och icke träder in på syndares väg, ej heller sitter där bespottare sitta,
utan har sin lust i HERRENS lag och tänker på hans lag både dag och natt.
Han är såsom ett träd, planterat vid vattenbäckar, vilket bär sin frukt i sin tid, och vars löv icke vissna; och allt vad han gör, det lyckas väl.
Icke så de ogudaktiga, utan de äro såsom agnar som vinden bortför.
Därför skola de ogudaktiga icke bestå i domen, ej heller syndarna i de rättfärdigas församling.
Ty HERREN känner de rättfärdigas väg, men de ogudaktigas väg förgås.
Varför larma hedningarna och tänka folken fåfänglighet?
Jordens konungar resa sig upp, och furstarna rådslå med varandra, mot HERREN och hans smorde:
»Låt oss slita sönder deras bojor och kasta deras band ifrån oss.»
Han som bor i himmelen ler, HERREN bespottar dem.
Då talar han till dem i sin vrede, och i sin förgrymmelse förskräcker han dem:
»Jag själv har insatt min konung på Sion, mitt heliga berg.»
Jag vill förtälja om vad beslutet är; HERREN sade till mig: »Du är min son, jag har i dag fött dig.
Begär av mig, så skall jag giva dig hedningarna till arvedel och jordens ändar till egendom.
Du skall sönderslå dem med järnspira, såsom lerkärl skall du krossa dem.»
Så kommen nu till förstånd, I konungar; låten varna eder, I domare på jorden.
Tjänen HERREN med fruktan, och fröjden eder med bävan.
Hyllen sonen, så att han icke vredgas och I förgåns på eder väg; ty snart kunde hans vrede upptändas.
Saliga äro alla de som taga sin tillflykt till honom.
En psalm av David, när han flydde för sin son Absalom.
HERRE, huru många äro icke mina ovänner!
Ja, många resa sig upp mot mig.
Många säga om mig: »Det finnes ingen frälsning för honom hos Gud.»
Men du, HERRE, är en sköld för mig; du är min ära och den som upplyfter mitt huvud.
Jag höjer min röst och ropar till HERREN, och han svarar mig från sitt heliga berg.
Sela.
Jag lade mig och somnade in; jag har åter vaknat upp, ty HERREN uppehåller mig.
Jag fruktar icke för skaror av många tusen, som lägra sig mot mig runt omkring.
Stå upp, HERRE, fräls mig, min Gud; ty du slår alla mina fiender på kinden, du krossar de ogudaktigas tänder.
Hos HERREN är frälsningen; över ditt folk komme din välsignelse.
Sela.
För sångmästaren, med strängaspel; en psalm av David.
När jag ropar, så svara mig, du min rättfärdighets Gud, du som i trångmål skaffar mig rum; var mig nådig och hör min bön.
I herrar, huru länge skall min ära vara vänd i smälek, huru länge skolen I älska fåfänglighet och fara efter lögn?
Sela.
Besinnen dock att HERREN har utvalt åt sig den fromme; HERREN hör, när jag ropar till honom.
Vredgens, men synden icke; eftersinnen i edra hjärtan, på edra läger, och varen stilla.
Sela.
Offren rätta offer, och förtrösten på HERREN.
Många säga: »Vem skall låta oss se det gott är?»
Upplyft du över oss ditt ansiktes ljus, o HERRE.
Du giver mig glädje i hjärtat, större än andras, när de få säd och vin i myckenhet.
I frid vill jag lägga mig ned, och i frid skall jag somna in, ty du, HERRE, låter mig bo avskild och i trygghet.
För sångmästaren, till Nehilót; en psalm av David.
Lyssna till mina ord, HERRE; förnim min suckan.
Akta på mitt klagorop, du min konung och min Gud; ty till dig vill jag ställa min bön.
HERRE, bittida hör du nu min röst, bittida frambär jag mitt offer till dig och skådar efter dig.
Ty du är icke en Gud som har behag till ogudaktighet; den som är ond får icke bo hos dig.
De övermodiga bestå icke inför dina ögon; du hatar alla ogärningsmän.
Du förgör dem som tala lögn; de blodgiriga och falska äro en styggelse för HERREN.
Men jag får gå in i ditt hus, genom din stora nåd; jag får tillbedja i din fruktan, vänd mot ditt heliga tempel.
HERRE, led mig genom din rättfärdighet, för mina förföljares skull; gör din väg jämn för mig.
Ty i deras mun är intet visst, deras innersta är fördärv, en öppen grav är deras strupe, sin tunga göra de hal.
Döm dem, o Gud; må de komma på fall med sina anslag.
Driv bort dem för deras många överträdelsers skull, eftersom de äro gensträviga mot dig.
Men låt alla dem glädjas, som taga sin tillflykt till dig; evinnerligen må de jubla, ty du beskärmar dem; i dig må de fröjda sig, som hava ditt namn kärt.
Ty du, HERRE, välsignar den rättfärdige; du betäcker honom med nåd såsom med en sköld.
För sångmästaren, med strängaspel, till Seminit; en psalm av David.
HERRE, straffa mig icke i din vrede, och tukta mig icke i din förtörnelse.
Var mig nådig, HERRE, ty jag försmäktar; hela mig, HERRE, ty ända in i mitt innersta är jag förskräckt.
Ja, min själ är storligen förskräckt; ack HERRE, huru länge?
Vänd åter, HERRE, rädda min själ, fräls mig för din nåds skull.
Ty i döden tänker man icke på dig; vem tackar dig i dödsriket?
Jag är så trött av suckande; var natt fuktar jag min säng och väter mitt läger med mina tårar.
Av sorg är mitt öga förmörkat; det har åldrats för alla mina ovänners skull.
Viken bort ifrån mig, alla I ogärningsmän; ty HERREN har hört min högljudda gråt.
HERREN har hört min åkallan, min bön upptager HERREN.
Alla mina fiender skola komma på skam och storligen förskräckas; de skola vika tillbaka och komma på skam med hast.
En sång av David, som han sjöng till HERREN för benjaminiten Kus' ords skull.
HERRE, min Gud, till dig tager jag min tillflykt; fräls mig från alla mina förföljare och rädda mig,
så att de icke, såsom lejon, sönderslita min själ och rycka bort henne utan räddning.
HERRE, min Gud, har jag gjort sådant, och är orätt i mina händer,
har jag med ont vedergällt ned som höll frid med mig eller plundrat den som var min ovän utan sak,
så förfölje fienden min själ och tage henne fatt och trampe mitt liv till jorden och lägge min ära i stoftet.
Sela.
Stå upp, HERRE, i din vrede, res dig mot mina ovänners raseri och vakna upp till min hjälp, du som har påbjudit dom.
Må folkens församling omgiva dig, och må du över den vända åter till höjden.
HERREN håller dom över folken; skaffa mig rätt, HERRE, efter min rättfärdighet och ostrafflighet.
Låt de ogudaktigas ondska få en ände, men håll den rättfärdige vid makt; ty du, som prövar hjärtan och njurar, är en rättfärdig Gud.
Min sköld är i Guds hand; han frälsar de rättsinniga.
Gud är en rättfärdig domare och en Gud som dagligen vredgas.
Om någon icke vill omvända sig, så vässer han sitt svärd, sin båge spänner han och gör den redo;
och han riktar mot honom dödande skott, sina pilar gör han brinnande.
Se, denne är i födsloarbete med fördärv, han går havande med olycka, men han föder ett intet.
Han gräver en grop och gör den djup, men han faller själv i den grav som han gräver.
Den olycka han tänkte vålla vänder tillbaka på hans huvud, och över hans hjässa kommer hans ondska.
Jag vill tacka HERREN efter hans rättfärdighet och lovsjunga HERRENS, den Högstes, namn.
För sångmästaren, till Gittít; en psalm av David.
HERRE, vår Herre, huru härligt är icke ditt namn över hela jorden, du som har satt ditt majestät på himmelen!
Av barns och spenabarns mun har du upprättat en makt, för dina ovänners skull, till att nedslå fienden och den hämndgirige.
När jag ser din himmel, dina fingrars verk, månen och stjärnorna, som du har berett,
vad är då en människa, att du tänker på henne, eller en människoson, att du låter dig vårda om honom.
Dock gjorde du honom nästan till ett gudaväsen; med ära och härlighet krönte du honom.
Du satte honom till herre över dina händers verk; allt lade du under hans fötter:
får och oxar, allasammans, så ock vildmarkens djur,
fåglarna under himmelen och fiskarna i havet, vad som vandrar havens vägar.
HERRE, vår Herre, huru härligt är icke ditt namn över hela jorden!
För sångmästaren, till Mutlabbén; en psalm av David.
Jag vill tacka HERREN av allt mitt hjärta; jag vill förtälja alla dina under.
Jag vill vara glad och fröjdas i dig, jag vill lovsjunga ditt namn, du den Högste.
Ty mina fiender vika tillbaka, de falla och förgås för ditt ansikte.
Ja, du har utfört min rätt och min sak; du sitter på din tron såsom en rättfärdig domare.
Du har näpst hedningarna och förgjort de ogudaktiga; deras namn har du utplånat för alltid och evinnerligen.
Fienderna äro nedgjorda, utrotade för alltid; deras städer har du omstörtat, deras åminnelse har förgåtts.
Men HERREN tronar evinnerligen, sin stol har han berett till doms;
och han skall döma jordens krets med rättfärdighet, han skall skipa lag bland folken med rättvisa.
Så vare då HERREN en borg för den förtryckte, en borg i nödens tider.
Och må de som känna ditt namn förtrösta på dig; ty du övergiver icke dem som söka dig, HERRE.
Lovsjungen HERREN, som bor i Sion, förkunnen bland folken hans gärningar.
Ty han som utkräver blodskulder har kommit ihåg dem; han har icke förgätit de betrycktas klagorop.
Var mig nådig, HERRE; se huru jag plågas av dem som hata mig, du som lyfter mig upp från dödens portar;
på det att jag må förtälja allt ditt lov och i dottern Sions portar fröjda mig över din frälsning.
Hedningarna hava sjunkit ned i den grav som de grävde; i det nät som de lade ut har deras fot blivit fångad.
HERREN har gjort sig känd, han har hållit dom; han snärjer den ogudaktige i hans händers verk.
Higgajón.
Sela.
DE ogudaktiga vika tillbaka, ned i dödsriket, alla hedningar, de som förgäta Gud.
Ty icke för alltid skall den fattige vara förgäten, de betrycktas hopp skall ej varda om intet evinnerligen.
Stå upp, HERRE; låt icke människor få överhanden, låt hedningarna bliva dömda inför ditt ansikte.
Låt, o HERRE, förskräckelse komma över dem; må hedningarna förnimma att de äro människor.
Sela.
Varför, HERRE, står du så långt ifrån och fördöljer dig i nödens tider?
Genom de ogudaktigas övermod måste den arme lida.
Må de fångas i de ränker som de hava uttänkt!
Ty den ogudaktige berömmer sig av sin själs lystnad, och den rovgirige talar förgripligt och föraktar HERREN.
Den ogudaktige säger i sitt högmod: »Han frågar icke därefter.» »Det finnes ingen Gud», så äro alla hans tankar.
Trygga äro alltid hans vägar, dina domar gå högt över hans blickar; alla sina ovänner räknar han för intet.
Han säger i sitt hjärta: »Jag skall icke vackla, över mig skall i evighet ingen olycka komma.»
Hans mun är full av förbannelse, av svek och förtryck; hans tunga gömmer olycka och fördärv.
Han lägger sig i försåt vid gårdarna, i lönndom vill han dräpa den oskyldige; hans ögon lura på den olycklige.
Han ligger i försåt på lönnligt ställe, såsom ett lejon i sitt snår, han ligger i försåt för att gripa den arme; han griper den arme, i det han drager honom in i sitt nät.
Han trycker sig ned, han ligger på lur, och de olyckliga falla i hans klor.
Han säger i sitt hjärta: »Gud förgäter det, han har dolt sitt ansikte, han ser det aldrig.»
Stå upp, HERRE; Gud, upplyft din hand, förgät icke de arma.
Varför skall den ogudaktige få förakta Gud och säga i sitt hjärta att du icke frågar därefter?
Du har ju sett det, ty du giver akt på olycka och jämmer, för att taga det i din hand.
Åt dig överlämnar den olycklige sin sak; du blev den faderlöses hjälpare.
Bryt sönder den ogudaktiges arm, och hemsök de ondas ogudaktighet, så att du icke mer finner den.
Ja, HERREN är konung alltid och evinnerligen; hedningarna utrotas ur hans land.
De ödmjukas trängtan hör du, HERRE; du gör deras hjärtan ståndaktiga; du låter ditt öra giva akt
för att skaffa den faderlöse och förtryckte rätt, så att människor, komna av jord, ej längre vålla skräck.
För sångmästaren; av David.
Till HERREN Har jag tagit min tillflykt.
Huru kunnen I då säga till mig: »Flyn såsom fåglar till edert berg;
ty se, de ogudaktiga spänna bågen, de hava lagt sin pil på strängen, för att i mörkret skjuta på de rättsinniga.
När grundvalarna upprivas, vad kan då den rättfärdige uträtta?»
HERREN är i sitt heliga tempel, HERRENS tron är i himmelen; hans ögon skåda, hans blickar pröva människors barn.
HERREN prövar den rättfärdige; men den ogudaktige och den som älskar våld, dem hatar hans själ.
Han skall låta ljungeldssnaror regna över de ogudaktiga; eld och svavel och glödande vind, det är den kalk som bliver dem beskärd.
Ty HERREN är rättfärdig, han älskar rättfärdigheten; de redliga skola skåda hans ansikte.
För sångmästaren, till Seminít; en psalm av David.
Fräls, HERRE; ty de fromma äro borta, de trogna äro försvunna ifrån människors barn.
De tala lögn, den ene med den andre; med hala läppar tala de, och med dubbelt hjärta.
HERREN utrote alla hala läppar, den tunga som talar stora ord,
dem som säga: »Genom vår tunga äro vi starka, våra läppar stå oss bi; vem är herre över oss?»
»Eftersom de arma lida övervåld och de fattiga klaga, vill jag nu stå upp», säger HERREN; »jag vill skaffa frälsning åt den som längtar därefter.»
HERRENS tal är ett rent tal, likt silver som rinner ned mot jorden, luttrat i degeln, renat sju gånger.
Du, HERRE, skall bevara dem, du skall beskydda dem för detta släkte evinnerligen.
Ty runt omkring dem vandra de ogudaktiga, då nu uselheten är rådande bland människors barn.
För sångmästaren; en psalm av David.
Huru länge, HERRE; skall du så alldeles förgäta mig?
Huru länge skall du fördölja ditt ansikte för mig?
Huru länge skall jag bekymras i min själ och ängslas i mitt hjärta dagligen?
Huru länge skall min fiende förhäva sig över mig?
Skåda ned, svara mig, HERRE, min Gud; upplys mina ögon, så att jag icke somnar in i döden;
på det att min fiende icke må säga: »Jag blev honom övermäktig», och på att mina ovänner ej må fröjda sig, när jag vacklar.
Jag förtröstar på din nåd, mitt hjärta fröjde sig över din frälsning.
Jag vill sjunga till HERRENS ära, ty han har gjort väl mot mig.
För sångmästaren; av David.
Dårarna säga i sina hjärtan: »Det finnes ingen Gud.»
Fördärv och styggelse är deras verk; ingen finnes, som gör vad gott är.
HERREN skådar ned från himmelen på människors barn, för att se om det finnes någon förståndig, någon som söker Gud.
Nej, alla äro de avfälliga, allasammans äro de fördärvade; ingen finnes, som gör vad gott är, det finnes icke en enda.
Hava de då intet fått förnimma, alla dessa ogärningsmän, dessa som uppäta mitt folk, likasom åte de bröd, och som icke åkalla HERREN?
Jo, där överföll dem förskräckelse -- ty Gud är hos de rättfärdigas släkte.
Den betrycktes rådslag mån I söka bringa på skam, HERREN är ju ändå hans tillflykt.
Ack att från Sion komme frälsning för Israel!
När HERREN vill åter upprätta sitt folk, då skall Jakob fröjda sig, då skall Israel vara glad.
En psalm av David.
HERRE, vem får bo i din hydda?
Vem får dväljas på ditt heliga berg?
Den som vandrar ostraffligt och gör vad rätt är och talar sanning av hjärtat;
den som icke bär förtal på sin tunga, den som icke gör sin broder något ont och icke drager smälek över sin nästa;
den som aktar den förkastlige för intet, men ärar dem som frukta HERREN; den som svär sig till skada, men ej bryter sin ed;
den som icke driver ocker med sina penningar och icke tager mutor för att fälla den oskyldige.
Den som så handlar, han skall icke vackla till evig tid.
En sång av David.
Bevara mig, Gud, ty jag tager min tillflykt till dig.
Jag säger till HERREN: »Du är ju Herren; för mig finnes intet gott utom dig;
de heliga som finnas i landet, de äro de härliga till vilka jag har allt mitt behag.»
Men de som taga sig en annan gud, de hava stora vedermödor; jag vill icke offra deras drickoffer av blod eller taga deras namn på mina läppar.
HERREN är min beskärda del och bägare; du är den som uppehåller min arvedel.
En lott har tillfallit mig i det ljuvliga, ja, ett arv som behagar mig väl.
Jag vill lova HERREN, ty han giver mig råd; ännu om natten manar mig mitt innersta.
Jag har haft HERREN för mina ögon alltid; ja, han är på min högra sida, jag skall icke vackla.
Fördenskull gläder sig mitt hjärta, och min ära fröjdar sig; jämväl min kropp får bo i trygghet.
Ty du skall icke lämna min själ åt dödsriket, du skall icke låta din fromme få se graven.
Du skall kungöra mig livets väg; inför ditt ansikte är glädje till fyllest, ljuvlighet i din högra hand evinnerligen.
En bön av David.
Hör, o HERRE, en rättfärdig sak, akta på mitt rop, lyssna till min bön; den kommer icke ifrån falska läppar.
Av dig må jag få min rätt; dina ögon må skåda vad rättvist är.
Du prövar mitt hjärta, du utrannsakar mig, men du finner intet; ingen ond tanke går ut ur min mun.
Efter dina läppars ord, och vad människor än må göra, tager jag mig till vara för våldsverkares stigar.
Mina steg hålla sig stadigt på dina vägar, mina fötter vackla icke.
Så åkallar jag nu dig, ty du, Gud, skall svara mig; böj ditt öra till mig, hör mitt tal.
Bevisa din underbara nåd, du som frälsar undan motståndarna dem som taga sin tillflykt till din högra hand.
Bevara mig såsom en ögonsten, beskärma mig under dina vingars skugga
för de ogudaktiga, som vilja fördärva mig, för mina dödsfiender, som omringa mig.
Sitt hjärta förstocka de; med sin mun tala de stora ord.
Nu äro de omkring mig, var vi gå, deras ögon speja efter huru de skola böja mig till jorden.
Ja, denne är lik ett lejon som längtar efter rov, lik ett ungt lejon som ligger i försåt.
Stå upp, HERRE; träd emot honom, slå honom ned, rädda med ditt svärd min själ från den ogudaktige,
ja, med din hand, från människorna, HERRE, från denna världens människor, som hava sin del i detta livet, och vilkas buk du fyller med dina håvor, som hava söner i mängd och lämna sitt överflöd åt sina barn.
Men jag skall skåda ditt ansikte i rättfärdighet; när jag uppvaknar, vill jag mätta mig av din åsyn.
För sångmästaren; av HERRENS tjänare David, som talade till HERREN denna sångs ord, när HERREN hade räddat honom från alla hans fienders hand och ur Sauls våld.
Han sade: Hjärtligen kär har jag dig, HERRE, min starkhet,
HERRE, mitt bergfäste, min borg och min räddare, min Gud, min klippa, till vilken jag tager min tillflykt, min sköld och min frälsnings horn, mitt värn.
HERREN, den högtlovade, åkallar jag, och från mina fiender bliver jag frälst.
Dödens band omvärvde mig, och fördärvets strömmar förskräckte mig.
Dödsrikets band omslöto mig, dödens snaror föllo över mig.
Men jag åkallade HERREN i min nöd och ropade till min Gud.
Han hörde från sin himmelska boning min röst, och mitt rop inför honom kom till hans öron.
Då skalv jorden och bävade, och bergens grundvalar darrade; de skakades, ty hans vrede var upptänd.
Rök steg upp från hans näsa och förtärande eld från hans mun; eldsglöd ljungade från honom.
Och han sänkte himmelen och for ned, och töcken var under hans fötter.
Han for på keruben och flög, han svävade på vindens vingar.
Han gjorde mörker till sitt täckelse, till en hydda som omslöt honom; mörka vatten, tjocka moln.
Av glansen framför honom veko molnen undan; hagel föll, och eldsglöd for ned.
Och HERREN dundrade i himmelen, den Högste lät höra sin röst; hagel föll, och eldsglöd for ned.
Han sköt sina pilar och förskingrade dem, ljungeldar i mängd och förvirrade dem.
Vattnens bäddar kommo i dagen, och jordens grundvalar blottades, för din näpst, o HERRE, för din vredes stormvind.
Han räckte ut sin hand från höjden och fattade mig, han drog mig upp ur de stora vattnen.
Han räddade mig från min starke fiende och från mina ovänner, ty de voro mig övermäktiga.
De överföllo mig på min olyckas dag, men HERREN blev mitt stöd.
Han förde mig ut på rymlig plats; han räddade mig, ty han hade behag till mig.
HERREN lönar mig efter min rättfärdighet; efter mina händers renhet vedergäller han mig.
Ty jag höll mig på HERRENS vägar och avföll icke från min Gud i ogudaktighet;
nej, alla hans rätter hade jag för ögonen, och hans stadgar lät jag icke vika ifrån mig.
Så var jag ostrafflig inför honom och tog mig till vara för missgärning.
Därför vedergällde mig HERREN efter min rättfärdighet, efter mina händers renhet inför hans ögon.
Mot den fromme bevisar du dig from, mot en ostrafflig man bevisar du dig ostrafflig.
Mot den rene bevisar du dig ren, men mot den vrånge bevisar du dig avog.
Ty du frälsar ett betryckt folk, men stolta ögon ödmjukar du.
Ja, du låter min lampa brinna klart; HERREN, min Gud, gör mitt mörker ljuset.
Ja, med dig kan jag nedslå härskaror, och med min Gud stormar jag murar.
Guds väg är ostrafflig; HERRENS tal är luttrat.
En sköld är han för alla som taga sin tillflykt till honom.
Ty vem är Gud förutom HERREN, och vem är en klippa utom vår Gud?
Gud, du som omgjordade mig med kraft och lät min väg vara lyckosam,
du som gjorde mina fötter såsom hindens och ställde mig på mina höjder,
du som lärde mina händer att strida och mina armar att spänna kopparbågen!
Du gav mig din frälsnings sköld, och din högra hand stödde mig, och ditt saktmod gjorde mig stor;
du skaffade rum för mina steg, där jag gick, och mina fötter vacklade icke.
Jag förföljde mina fiender och hann upp dem; jag vände icke tillbaka, förrän jag hade gjort ände på dem.
Jag slog dem, så att de icke mer kunde resa sig; de föllo under mina fötter.
Du omgjordade mig med kraft till striden, du böjde mina motståndare under mig.
Mina fiender drev du på flykten för mig, och dem som hatade mig förgjorde jag.
De ropade, men det fanns ingen som frälste; till HERREN, men han svarade dem icke.
Och jag stötte dem sönder till stoft för vinden, jag kastade ut dem såsom orenlighet på gatan.
Du räddade mig ur folkets strider, du satte mig till ett huvud över hedningar; folkslag som jag ej kände blevo mina tjänare.
Vid blotta ryktet hörsammade de mig; främlingar visade mig underdånighet.
Ja, främlingarnas mod vissnade bort; med bävan övergåvo de sina borgar.
HERREN lever!
Lovad vare min klippa, och upphöjd vare min frälsnings Gud!
Gud, som har givit mig hämnd och tvingat folken under mig;
du som har befriat mig från mina fiender och upphöjt mig över mina motståndare, räddat mig från våldets man!
Fördenskull vill jag tacka dig bland hedningarna, HERRE, och lovsjunga ditt namn.
Ty du giver din konung stor seger och gör nåd mot din smorde, mot David och hans säd till evig tid.
För sångmästaren; en psalm av David.
Himlarna förtälja Guds ära, och fästet förkunnar hans händers verk;
den ena dagen talar därom till den andra, och den ena natten kungör det för den andra;
det är ej ett tal eller språk vars ljud icke höres.
De sträcka sig ut över hela jorden, och deras ord gå till världens ändar.
Åt solen har han gjort en hydda i dem;
och den är såsom en brudgum som går ut ur sin kammare, den fröjdar sig, såsom en hjälte, att löpa sin bana.
Vid himmelens ända är det den går upp, och dess omlopp når intill himmelens gränser, och intet är skylt för dess hetta.
HERRENS lag är utan brist och vederkvicker själen; HERRENS vittnesbörd är fast och gör den enfaldige vis.
HERRENS befallningar äro rätta och giva glädje åt hjärtat; HERRENS bud är klart och upplyser ögonen.
HERRENS fruktan är ren och består evinnerligen; HERRENS rätter äro sanning, allasammans rättfärdiga.
De äro dyrbarare än guld, ja, än fint guld i mängd; de äro sötare än honung, ja, än renaste honung.
Av dem hämtar ock din tjänare varning; den som håller dem har stor lön.
Vem märker själv huru ofta han felar?
Förlåt mig mina hemliga brister.
Bevara ock din tjänare för fräcka människor; låt dem icke få makt med mig, så bliver jag ostrafflig och varder fri ifrån svår överträdelse.
Låt min muns tal täckas dig och mitt hjärtas tankar, HERRE, min klippa och min förlossare.
För sångmästaren; en psalm av David.
HERREN bönhöre dig på nödens dag, Jakobs Guds namn beskydde dig.
Han sände dig hjälp från helgedomen, och stödje dig från Sion.
Han tänke på alla dina spisoffer och upptage med välbehag ditt brännoffer.
Sela.
Han give dig vad ditt hjärta begär och fullborde alla dina rådslag.
Må vi få jubla över din seger och i vår Guds namn resa upp baneret; HERREN uppfylle alla dina böner.
Nu vet jag att HERREN giver seger åt sin smorde; han svarar honom från sin heliga himmel, genom väldiga gärningar giver hans högra hand seger.
De andra prisa vagnar, de prisa hästar, men vi prisa HERRENS, vår Guds, namn.
De sjunka ned och falla, men vi resa oss upp och bliva beståndande.
HERRE, giv seger; ja, konungen svare oss på den tid då vi ropa.
För sångmästaren; en psalm av David.
HERRE, över din makt gläder sig konungen; huru fröjdas han icke högeligen över din seger!
Vad hans hjärta önskar har du givit honom, och hans läppars begäran har du icke vägrat honom.
Sela.
Ty du kommer honom till mötes med välsignelser av vad gott är; du sätter på hans huvud en gyllene krona.
Han bad dig om liv, och du gav honom det, ett långt liv alltid och evinnerligen.
Stor är hans ära genom din seger; majestät och härlighet beskär du honom.
Ja, du låter honom bliva till välsignelse evinnerligen; du fröjdar honom med glädje inför ditt ansikte.
Ty konungen förtröstar på HERREN, och genom den Högstes nåd skall han icke vackla.
Din hand skall nå alla dina fiender; din högra hand skall träffa dem som hata dig.
Du skall låta dem känna det såsom i en glödande ugn, när du låter se ditt ansikte.
HERREN skall fördärva dem i sin vrede; eld skall förtära dem.
Deras livsfrukt skall du utrota från jorden och deras avkomma från människors barn.
Ty de ville draga ont över dig; de tänkte ut ränker, men de förmå intet.
Nej, du skall driva dem tillbaka; med din båge skall du sikta mot deras anleten.
Upphöjd vare du, HERREN, i din makt; vi vilja besjunga och lovsäga din hjältekraft.
För sångmästaren, efter »Morgonrodnadens hind»; en psalm av David.
Min Gud, min Gud, varför har du övergivit mig?
Jag brister ut och klagar, men min frälsning är fjärran.
Men Gud, jag ropar om dagen, men du svarar icke, så ock om natten, men jag får ingen ro.
Och dock är du den Helige, den som tronar på Israels lovsånger.
På dig förtröstade våra fäder; de förtröstade, och du räddade dem.
Till dig ropade de och blevo hulpna; på dig förtröstade de och kommo icke på skam.
Men jag är en mask, och icke en människa, till smälek bland män, föraktad av folket.
Alla som se mig bespotta mig; de spärra upp munnen, de skaka huvudet:
»Befall dig åt HERREN!
Han befrie honom, han rädde honom, ty han har ju behag till honom.»
Ja, det var du som hämtade mig ut ur moderlivet och lät mig vila trygg vid min moders bröst.
På dig är jag kastad allt ifrån modersskötet; du är min Gud allt ifrån min moders liv.
Var icke långt ifrån mig, ty nöd är nära, och det finnes ingen hjälpare.
Tjurar i mängd omgiva mig, Basans oxar omringa mig.
Såsom glupande och rytande lejon spärrar man upp gapet mot mig.
Jag är lik vatten som utgjutes, alla mina leder hava skilts åt; mitt hjärta är såsom vax, det smälter i mitt liv.
Min kraft är förtorkad och lik en lerskärva, min tunga låder vid min gom, och du lägger mig i dödens stoft.
Ty hundar omgiva mig; de ondas hop har kringränt mig, mina händer och fötter hava de genomborrat.
Jag kan räkna alla mina ben; de skåda därpå, de se med lust på mig.
De dela mina kläder mellan sig och kasta lott om min klädnad.
Men du, HERRE, var icke fjärran; du min starkhet, skynda till min hjälp.
Rädda min själ från svärdet, mitt liv ur hundarnas våld.
Fräls mig från lejonets gap.
Ja, du bönhör mig och räddar mig undan vildoxarnas horn.
Då skall jag förkunna ditt namn för mina bröder, mitt i församlingen skall jag prisa dig:
I som frukten HERREN, loven honom; ären honom, alla Jakobs barn, och bäven för honom, alla Israels barn.
Ty han föraktade icke den betrycktes elände och höll det icke för en styggelse; han fördolde icke sitt ansikte för honom, och när han ropade, lyssnade han till honom.
Genom dig skall min lovsång ljuda i den stora församlingen; mina löften får jag infria inför dem som frukta honom.
De ödmjuka skola äta och bliva mätta, de som söka HERREN skola få lova honom; ja, edra hjärtan skola leva evinnerligen.
Alla jordens ändar skola betänka det och omvända sig till HERREN.
Hedningarnas alla släkter skola tillbedja inför dig.
Ty riket är HERRENS, och han råder över hedningarna.
Ja, alla mäktiga på jorden skola äta och tillbedja; inför honom skola knäböja alla de som måste fara ned i graven, de som icke kunna behålla sin själv vid liv.
Kommande ättled skola tjäna honom; man skall förtälja om Herren för ett annat släkte.
Man skall träda upp och förkunna hans rättfärdighet, ja, bland folk som skola födas att han har gjort det.
En psalm av David.
HERREN är min herde, mig skall intet fattas,
han låter mig vila på gröna ängar; han för mig till vatten där jag finner ro,
han vederkvicker min själ; han leder mig på rätta vägar, för sitt namns skull.
Om jag ock vandrar i dödsskuggans dal, fruktar jag intet ont, ty du är med mig; din käpp och stav, de trösta mig.
Du bereder för mig ett bord i mina ovänners åsyn; du smörjer mitt huvud med olja och låter min bägare flöda över.
Godhet allenast och nåd skola följa mig i alla mina livsdagar, och jag skall åter få bo i HERRENS hus, evinnerligen.
Av David; en psalm.
Jorden är HERRENS och allt vad därpå är, jordens krets och de som bo därpå.
Ty han är den som har lagt hennes grund på haven, den som på strömmarna har berett henne fäste.
Vem får gå upp på HERRENS berg, och vem får träda in i hans helgedom?
Den som har oskyldiga händer och rent hjärta, den som icke vänder sin själ till lögn och den som icke svär falskt.
Han skall undfå välsignelse av HERREN och rättfärdighet av sin frälsnings Gud.
Sådant är det släkte som frågar efter honom; de som söka ditt ansikte, de äro Jakobs barn.
Sela.
Höjen, I portar, edra huvuden, höjen eder, I eviga dörrar, för att ärans konung må draga därin.
Vem är då ärans konung?
Det är HERREN, stark och väldig, HERREN, väldig i strid.
Höjen, I portar, edra huvuden, höjen dem, I eviga dörrar, för att ärans konung må draga därin.
Vem är då denne ärans konung?
Det är HERREN Sebaot; han är ärans konung.
Sela.
Av David.
Till dig, HERRE, upplyfter jag min själ.
Min Gud, på dig förtröstar jag; låt mig icke komma på skam, låt icke mina fiender fröjda sig över mig.
Nej, ingen kommer på skam, som förbidar dig; på skam kommer de som, utan sak, handla trolöst.
HERRE, kungör mig dina vägar, lär mig dina stigar.
Led mig i din sanning, och lär mig, ty du är min frälsnings Gud; dig förbidar jag alltid.
Tänk, HERRE, på din barmhärtighet och din nåd, ty de äro av evighet.
Tänk icke på min ungdoms synder och på mina överträdelser, utan tänk på mig efter din nåd, för din godhets skull, HERRE.
HERREN är god och rättfärdig, därför undervisar han syndare om vägen.
Han leder de ödmjuka rätt, han lär de ödmjuka sin väg.
Alla HERRENS vägar äro nåd och trofasthet för dem som hålla hans förbund och vittnesbörd.
För ditt namns skull, HERRE, förlåt min missgärning, ty den är stor.
Finnes det en man som fruktar HERREN, då undervisar han honom om den väg han bör välja.
Han själv skall leva i lycka, och hans efterkommande skola besitta landet.
HERREN har sin umgängelse med dem som frukta honom, och sitt förbund vill han kungöra för dem.
Mina ögon se alltid till HERREN, ty han drager mina fötter ur nätet.
Vänd dig till mig och var mig nådig; ty jag är ensam och betryckt.
Mitt hjärtas ångest är stor; för mig ut ur mitt trångmål.
Se till mitt lidande och min vedermöda, och förlåt mig alla mina synder.
Se därtill att mina fiender äro så många och hata mig med orätt.
Bevara min själ och rädda mig; låt mig icke komma på skam, ty jag tager min tillflykt till dig.
Ostrafflighet och redlighet bevare mig, ty jag förbidar dig.
Förlossa Israel, o Gud, ur all dess nöd.
Av David.
Skaffa mig rätt, HERRE, ty jag vandrar i ostrafflighet, och jag förtröstar på HERREN utan att vackla.
Pröva mig, HERRE, och försök mig; rannsaka mina njurar och mitt hjärta.
Ty din nåd är inför mina ögon, och jag vandrar i din sanning.
Jag sitter icke hos lögnens män, och med hycklare har jag icke min umgängelse.
Jag hatar de ondas församling, och hos de ogudaktiga sitter jag icke.
Jag tvår mina händer i oskuld, och kring ditt altare, HERRE, vill jag vandra,
för att höja min röst till tacksägelse och förtälja alla dina under.
HERRE, jag har din boning kär och den plats där din härlighet bor.
Ryck icke min själ bort med syndare, icke mitt liv med de blodgiriga,
i vilkas händer är skändlighet, och vilkas högra hand är full av mutor.
Jag vandrar ju i ostrafflighet; förlossa mig och var mig nådig.
Ja, min fot står på jämn mark; i församlingarna skall jag lova HERREN.
Av David.
HERREN är mitt ljus och min frälsning; för vem skulle jag frukta?
HERREN är mitt livs värn; för vem skulle jag rädas?
När de onda draga emot mig och vilja uppsluka mig, då stappla de själva och falla, mina motståndare och fiender.
Om ock en här lägrar sig mot mig, så fruktar ändå icke mitt hjärta; om krig uppstår mot mig, så är jag dock trygg.
Ett har jag begärt av HERREN, därefter traktar jag: att jag må få bo i HERRENS hus i alla mina livsdagar, för att skåda HERRENS ljuvlighet och betrakta hans tempel.
Ty han döljer mig i sin hydda på olyckans dag, han beskärmar mig i sitt tjäll, han för mig upp på en klippa.
Och nu skall mitt huvud resa sig över mina fiender runt omkring mig, och jag vill offra i hans hydda jublets offer, jag vill sjunga till HERRENS ära och lovsäga honom.
Hör, o HERRE!
Jag höjer min röst och ropar, var mig nådig och svara mig.
Mitt hjärta förehåller dig ditt ord: »Söken mitt ansikte.»
Ja, ditt ansikte, HERRE, söker jag;
fördölj icke ditt ansikte för mig.
Driv icke bort din tjänare i vrede, du som har varit min hjälp; förskjut mig icke, övergiv mig icke, du min frälsnings Gud.
Nej, om än min fader och min moder övergiva mig, skall HERREN upptaga mig.
Visa mig, HERRE, din väg, och led mig på en jämn stig, för mina förföljares skull.
Överlämna mig icke åt mina ovänners vilja; ty mot mig uppstå falska vittnen och män som andas våld.
Ja, jag tror förvisso att jag skall få se HERRENS goda i de levandes land.
Förbida HERREN, var frimodig och oförfärad i ditt hjärta; ja, förbida HERREN.
Av David.
Till dig, HERRE, ropar jag; min klippa, var icke stum mot mig.
Ja, var icke tyst mot mig, så att jag bliver lik dem som fara ned i graven.
Hör mina böners ljud, när jag ropar till dig, när jag upplyfter mina händer mot det allraheligaste i din helgedom.
Tag mig icke bort med de ogudaktiga och med ogärningsmännen, som tala vänligt med sin nästa men hava ondska i sina hjärtan.
Giv dem efter deras gärningar och efter deras onda väsende, giv dem efter deras händers verk, vedergäll dem vad de hava gjort.
Ty de akta icke på HERRENS gärningar, icke på hans händer verk; därför skall han slå dem ned och ej mer bygga upp dem.
Lovad vare HERREN, ty han har hört mina böners ljud!
HERREN är min starkhet och min sköld; på honom förtröstade mitt hjärta.
Och jag vart hulpen, därför fröjdar sig mitt hjärta, och med min sång vill jag tacka honom.
HERREN är sitt folks starkhet, och ett frälsningens värn är han för sin smorde.
Fräls ditt folk och välsigna din arvedel, och var deras herde och bär dem till evig tid.
En psalm av David.
Given åt HERREN, I Guds sönder, given åt HERREN ära och makt;
given åt HERREN hans namns ära, tillbedjen HERREN i helig skrud.
HERRENS röst går ovan vattnen; Gud, den härlige, dundrar, ja, HERREN, ovan de stora vattnen.
HERRENS röst ljuder med makt, HERRENS röst ljuder härligt.
HERRENS röst bräcker cedrar, HERREN bräcker Libanons cedrar.
Han kommer dem att hoppa likasom kalvar, Libanon och Sirjon såsom unga vildoxar.
HERRENS röst sprider ljungeldslågor.
HERRENS röst kommer öknen att bäva, HERREN kommer Kades' öken att bäva.
HERRENS röst bringar hindarna att föda; skogarnas klädnad rycker den bort.
I hans himmelska boning förkunnar allting hans ära.
HERREN på sin tron bjöd floden komma, och HERREN tronar såsom konung evinnerligen.
HERREN skall giva makt åt sitt folk, HERREN skall välsigna sitt folk med frid.
En psalm, en sång av David, vid templets invigning.
Jag vill upphöja dig, HERRE, ty du har dragit mig ur djupet, du har icke låtit mina fiender glädja sig över mig.
HERRE, min Gud, jag ropade till dig, och du helade mig.
HERRE, du förde min själ upp ur dödsriket, du tog mig levande ut från dem som foro ned i graven.
Lovsjungen HERREN, I hans fromme, och prisen hans heliga namn.
Ty ett ögonblick varar hans vrede, men hela livet hans nåd; om aftonen gästar gråt, men om morgonen kommer jubel.
Jag sade, när det gick mig väl: »Jag skall aldrig vackla.»
HERRE, i din nåd hade du gjort mitt berg starkt; men du fördolde ditt ansikte, då förskräcktes jag.
Till dig, HERRE, ropade jag, och till Herren bad jag:
»Vad vinning har du av mitt blod, eller därav att jag far ned i graven?
Kan stoftet tacka dig, kan det förkunna din trofasthet?
Hör, o HERRE, och var mig nådig; HERRE, var min hjälpare.»
Då förvandlade du min klagan i fröjdesprång; du klädde av mig sorgens dräkt och omgjordade mig med glädje.
Därför skall min ära lovsjunga dig, utan att tystna; HERRE, min Gud, jag vill tacka dig evinnerligen.
För sångmästaren; en psalm av David.
Till dig, HERRE, tager jag min tillflykt; låt mig aldrig komma på skam, befria mig genom din rättfärdighet.
Böj ditt öra till mig, rädda mig snarligen; var mig en fast klippa, en bort till min frälsning.
Ty du är mitt bergfäste och min bort, och du skall, för ditt namns skull, leda och föra mig.
Du skall draga mig ur det nät som de lade ut för mig; ty du är mitt värn.
I din hand befaller jag min ande; du förlossar mig, HERRE, du trofaste Gud.
Jag hatar dem som hålla sig till fåfängliga avgudar, men jag förtröstar på HERREN.
Jag vill fröjda mig och vara glad över din nåd, att du ser till mitt lidande, att du låter dig vårda om min själ i nöden
och icke överlämnar mig i fiendens hand, utan ställer mina fötter på rymlig plats.
Var mig nådig, HERRE, ty jag är i nöd; av sorg är mitt öga förmörkat, ja, min själ såväl som min kropp.
Ty mitt liv har försvunnit i bedrövelse och mina år i suckan; min kraft är bruten genom min missgärning, och benen i min kropp äro maktlösa.
För alla mina ovänners skull har jag blivit till smälek, ja, till stor smälek för mina grannar och till skräck för mina förtrogna; de som se mig på gatan fly undan för mig.
Jag är bortglömd ur hjärtat, såsom vore jag död; jag har blivit såsom ett sönderslaget kärl.
Ty jag hör mig förtalas av många; skräck från alla sidor!
De rådslå med varandra mot mig och stämpla för att taga mitt liv.
Men jag förtröstar på dig, HERRE; jag säger: »Du är min Gud.»
Min tid står i dina händer; rädda mig från mina fienders hand och mina förföljare.
Låt ditt ansikte lysa över din tjänare; fräls mig genom din nåd.
HERRE, låt mig icke komma på skam, ty jag åkallar dig; låt de ogudaktiga komma på skam och varda tystade i dödsriket.
Må lögnaktiga läppar förstummas, de som tala vad fräckt är mot den rättfärdige, med högmod och förakt.
Huru stor är icke din godhet, den du förvarar åt dem som frukta dig, och den du bevisar inför människors barn mot dem som taga sin tillflykt till dig!
Du beskärmar dem i ditt ansiktes beskärm mot människors sammangaddning; du döljer dem i din hydda mot tungors angrepp.
Lovad vare HERREN, ty han har bevisat mig sin underbara nåd genom att beskära mig en fast stad!
Ty väl sade jag i min ångest: »Jag är bortdriven från dina ögon.»
Likväl hörde du mina böners ljud, när jag ropade till dig.
Älsken HERREN, alla I hans fromme.
HERREN bevarar de trogna, men han vedergäller i fullt mått den som över högmod.
Varen frimodiga och oförfärade i edra hjärtan, alla I som sätten edert hopp till HERREN.
Av David; en sång.
Säll är den vilkens överträdelse är förlåten, vilkens synd är överskyld.
Säll är den människa som HERREN icke tillräknar missgärning, och i vilkens ande icke är något svek.
Så länge jag teg, försmäktade mina ben vid min ständiga klagan.
Ty dag och natt var din hand tung över mig; min livssaft förtorkades såsom av sommarhetta.
Sela.
Då uppenbarade jag min synd för dig och överskylde icke min missgärning.
Jag sade: »Jag vill bekänna för HERREN mina överträdelser»; då förlät du mig min synds missgärning.
Sela.
Därför skola alla fromma bedja till dig på den tid då du är att finna; sannerligen, om ock stora vattenfloder komma, skola de icke nå till dem.
Du är mitt beskärm, för nöd bevarar du mig; med räddningens jubel omgiver du mig.
Sela.
Jag vill lära dig och undervisa dig om den väg du skall vandra; jag vill giva dig råd och låta mitt öga vaka över dig.
Varen icke såsom hästar och mulåsnor utan förstånd, på vilka man lägger töm och betsel för att tämja dem, eljest får man dem ej fram.
Den ogudaktige har många plågor; men den som förtröstar på HERREN, honom omgiver han med nåd.
Varen glada i HERREN och fröjden eder, I rättfärdige, och jublen, alla I rättsinnige.
Jublen i HERREN, I rättfärdige; lovsång höves de redliga.
Tacken HERREN på harpa, lovsjungen honom till tiosträngad psaltare.
Sjungen honom en ny sång, spelen skönt med jubelklang.
Ty HERRENS ord är rätt, och allt vad han gör är gjort i trofasthet.
Han älskar rättfärdighet och rätt; jorden är full av HERRENS nåd.
Himmelen är gjord genom HERRENS ord och all dess här genom hans muns anda.
Han samlar havets vatten såsom i en hög; han lägger djupen i deras förvaringsrum.
Hela jorden frukte HERREN; för honom bäve alla som bo på jordens krets.
Ty han sade, och det vart; han bjöd, och det stod där.
HERREN gjorde hedningarnas råd om intet, han lät folkens tankar komma på skam.
Men HERRENS råd består evinnerligen, hans hjärtas tankar från släkte till släkte.
Saligt är det folk vars Gud HERREN är, det folk som han har utvalt till arvedel åt sig.
Ja, från himmelen skådade HERREN ned, han såg alla människors barn.
Från sin boning blickade han ned till alla dem som bo på jorden,
han som har danat allas deras hjärtan, han som aktar på alla deras verk.
En konung segrar icke genom sin stora styrka, en hjälte räddas icke genom sin stora kraft.
Förgäves väntar man sig seger genom hästar, med all sin styrka rädda de icke.
Se, HERRENS öga är vänt till dem som frukta honom, till dem som hoppas på hans nåd;
han vill rädda deras själ från döden och behålla dem vid liv i hungerns tid.
Vår själ väntar efter HERREN; han är vår hjälp och sköld.
Ty i honom gläder sig vårt hjärta, vi förtrösta på hans heliga namn.
Din nåd, HERRE, vare över oss, såsom vi hoppas på dig.
Av David, här han ställde sig vansinnig inför Abimelek, och denne drev honom ifrån sig, och han gick sin väg.
Jag vill lova HERREN alltid; hans pris skall ständigt vara i min mun.
Min själ skall berömma sig av HERREN; de ödmjuka skola höra det och glädja sig.
Loven med mig HERREN, låtom oss med varandra upphöja hans namn.
Jag sökte HERREN, och han svarade mig, och ur all min förskräckelse räddade han mig.
De som skåda upp till honom stråla av fröjd, och deras ansikten behöva icke rodna av blygsel.
Här är en betryckt som ropade, och HERREN hörde honom och frälste honom ur all hans nöd.
HERRENS ängel slår sitt läger omkring dem som frukta honom, och han befriar dem.
Smaken och sen att HERREN är god; säll är den som tager sin tillflykt till honom.
Frukten HERREN, I hans helige; ty de som frukta honom lida ingen brist.
Unga lejon lida nöd och hungra, men de som söka HERREN hava icke brist på något gott.
Kommen, barn, hören mig; jag skall lära eder HERRENS fruktan.
Är du en man som älskar livet och önskar att se goda dagar?
Avhåll då din tunga från det som är ont och dina läppar från att tala svek.
Vänd dig bort ifrån det som är ont, och gör vad gott är, sök friden och trakta därefter.
HERRENS ögon äro vända till de rättfärdiga och hans öron till deras rop.
Men HERRENS ansikte är emot dem som göra det onda, han vill utrota deras åminnelse från jorden.
När de rättfärdiga ropa, då hör HERREN och räddar dem ur all deras nöd.
HERREN är nära dem som hava ett förkrossat hjärta och frälsar dem som hava en bedrövad ande.
Den rättfärdige måste lida mycket, men HERREN räddar honom ur allt.
Han bevarar alla hans ben; icke ett enda av dem skall sönderslås.
Den ogudaktige skall dödas av olyckan, och de som hata den rättfärdige skola stå med skuld.
Men sina tjänares själar förlossar HERREN, och ingen skall stå med skuld, som tager sin tillflykt till honom.
Av David.
Gå till rätta, HERRE, med dem som gå till rätta med mig; strid mot dem som strida mot mig.
Fatta sköld och skärm, och stå upp till min hjälp;
drag fram spjutet, och spärra vägen för mina förföljare.
Säg till min själ: »Jag är din frälsning.»
Må de komma på skam och blygas, som stå efter mitt liv; må de vika tillbaka och varda utskämda, som hava ont i sinnet mot mig.
Må de bliva såsom agnar för vinden, och HERRENS ängel drive dem bort.
Deras väg blive mörk och slipprig, och HERRENS ängel drive dem bort.
Ty utan sak hava de försåtligen tillrett sin nätgrop för mig, utan sak hava de grävt en grav för mitt liv.
Fördärv komme över den mannen oförtänkt, det nät han har utlagt må fånga honom; ja, till sitt fördärv falle han själv däri.
Men min själ skall fröjda sig i HERREN och vara glad över hans frälsning.
Alla ben i min kropp skola säga: »HERRE, vem är dig lik, du som räddar den betryckte från den som är honom för stark, den betryckte och fattige ifrån den som plundrar honom?»
Orättfärdiga vittnen träda fram; de utfråga mig om det jag icke vet.
De löna mig med ont för gott; övergiven är min själ.
Jag åter bar sorgdräkt, när de voro sjuka, jag späkte min själ med fasta, jag bad med nedsänkt huvud;
såsom gällde det min vän, min broder, så skickade jag mig; lik den som sörjer sin moder gick jag sorgklädd och lutande.
Men de glädja sig över mitt fall och rota sig samman; ja, eländiga människor, som jag icke känner, rota sig samman mot mig, de smäda mig utan uppehåll.
Dessa gudlösa, som driva gyckel för en kaka bröd, bita ihop tänderna mot mig.
Herre, huru länge skall du se härpå?
Ryck min själ undan det fördärv de bereda, och mitt liv undan lejonen.
Då skall jag tacka dig i den stora församlingen, och bland mycket folk skall jag lova dig.
Låt icke dem få glädja sig över mig, som utan skäl äro mina fiender; låt icke dem som utan sak hata mig få blinka med ögonen.
Ty det är icke frid som de tala; nej, svekets ord tänka de ut mot de stilla i landet.
De spärra upp munnen mot mig; de säga: »Rätt så, rätt så, nu se vi det med egna ögon!»
Du, HERRE, ser det; tig icke.
Herre, var icke långt ifrån mig.
Vakna och stå upp för att skaffa mig rätt, för att utföra min sak, du min Gud och Herre.
Skaffa mig rätt efter din rättfärdighet, HERRE, min Gud, och låt dem icke få glädja sig över mig.
Låt dem icke säga i sina hjärtan: »Rätt så, det gick såsom vi ville!»
Låt dem icke säga: »Vi hava fördärvat honom.»
Må alla komma på skam och blygas, som glädja sig över min ofärd.
Med skam och blygd må de varda klädda, som förhäva sig över mig.
Men må de jubla och glädja sig, som unna mig min rätt, och må de alltid kunna säga: »Lovad vare HERREN, han som unnar sin tjänare gott!»
Då skall min tunga förkunna din rättfärdighet och hela dagen ditt lov.
För sångmästaren; av HERRENS tjänare David.
I mitt hjärta betänker jag vad synden säger till den ogudaktige, till den för vilkens ögon Guds fruktan ej finnes.
Den intalar ju honom vad som är behagligt i hans ögon: att man icke skall finna hans missgärning och hata den.
Hans muns ord äro fördärv och svek; han vill icke göra vad förståndigt och gott är.
Fördärv tänker han ut på sitt läger, han träder på den väg som icke är god; han skyr icke för något ont.
HERRE, upp i himmelen räcker din nåd, och din trofasthet allt upp till skyarna.
Din rättfärdighet är såsom väldiga berg, dina rätter såsom det stora havsdjupet; både människor och djur hjälper du, HERRE.
Huru dyrbar är icke din nåd, o Gud!
Människors barn hava sin tillflykt under dina vingars skugga.
De varda mättade av ditt hus' rika håvor, och av din ljuvlighets ström giver du dem att dricka.
Ty hos dig är livets källa, i ditt ljus se vi ljus.
Låt din nåd förbliva över dem som känna dig och din rättfärdighet över de rättsinniga.
Låt icke de högmodigas fot komma över mig eller de ogudaktigas hand driva mig bort.
Ja, där ligga ogärningsmännen fallna; de äro nedstötta och kunna icke mer resa sig.
Av David.
Harmas icke över de onda, avundas icke dem som göra orätt.
Ty såsom gräs varda de snart avhuggna, och såsom gröna örter vissna de.
Förtrösta på HERREN, och gör vad gott är, förbliv i landet och beflita dig om redbarhet,
och hav din lust i HERREN: då skall han giva dig vad ditt hjärta begär.
Befall din väg åt HERREN och förtrösta på honom; han skall göra det.
Han skall låta din rättfärdighet gå fram såsom ljuset och din rätt såsom middagens sken.
Var stilla för HERREN och förbida honom, harmas icke över den vilkens väg är lyckosam, över den man som umgås med ränker.
Avhåll dig från vrede och låt förbittringen fara; harmas icke; därmed gör du blott illa.
Ty de onda skola varda utrotade, men de som vänta efter HERREN, de skola besitta landet.
Ännu en liten tid, så är den ogudaktige icke mer; och när du ser efter hans plats, då är han borta.
Men de ödmjuka skola besitta landet och hugnas av stor frid.
Den ogudaktige stämplar mot den rättfärdige och biter sina tänder samman mot honom;
men Herren ler åt honom, ty han ser att hans dag kommer.
De ogudaktiga draga ut svärdet och spänna sin båge, för att fälla den som är betryckt och fattig, för att slakta dem som vandra i redlighet.
Men deras svärd skall gå in i deras eget hjärta, och deras bågar skola brista sönder.
Det lilla som en rättfärdig har är bättre än många ogudaktigas stora håvor.
Ty de ogudaktigas armar skola sönderbrytas; men HERREN uppehåller de rättfärdiga.
HERREN känner de frommas dagar, och deras arvedel skall bestå evinnerligen.
De skola icke komma på skam i den onda tiden, och i hungerns dagar skola de varda mättade.
Ty de ogudaktiga skola förgås; HERRENS fiender äro såsom ängarnas prakt: de försvinna såsom rök, ja, de försvinna.
Den ogudaktige lånar och kan icke betala, men den rättfärdige är barmhärtig och givmild.
Ty HERRENS välsignade skola besitta landet, men de som han förbannar skola varda utrotade.
Genom HERREN bliva en mans steg fasta, när han har behag till hans väg.
Om han faller, störtar han dock icke till marken, ty HERREN håller honom vid handen.
Jag har varit ung och är nu gammal, men jag har icke sett den rättfärdige övergiven eller hans barn gå efter bröd.
Han är alltid barmhärtig och villig att låna och hans barn äro till välsignelse.
Vänd dig bort ifrån det som är ont, och gör vad gott är, så skall du få bo kvar evinnerligen.
Ty HERREN älskar vad rätt är och övergiver icke sina fromma, evinnerligen bliva de bevarade; men de ogudaktigas avkomma varder utrotad.
De rättfärdiga skola besitta landet och bo däri evinnerligen.
Den rättfärdiges mun talar visdom, och hans tunga säger vad rätt är.
Hans Guds lag är i hans hjärta; hans steg vackla icke.
Den ogudaktige vaktar på den rättfärdige och står efter att döda honom,
men HERREN överlämnar honom icke i hans hand och fördömer honom icke, när han dömes.
Förbida HERREN, och håll dig på hans väg, så skall han upphöja dig till att besitta landet; du skall se med lust huru de ogudaktiga varda utrotade.
Jag såg en ogudaktig som trotsade på sin makt; han utbredde sig såsom ett grönskande träd, väl rotat.
Men när man sedan gick där fram, se, då var han borta; jag sökte efter honom, men han fanns icke mer.
Giv akt på den ostrafflige, och se på den redlige, huru fridens man har en framtid.
Men överträdarna skola allasammans förgås, de ogudaktigas framtid varder avskuren.
Till de rättfärdiga kommer frälsning ifrån HERREN; han är deras värn i nödens tid.
HERREN hjälper dem och befriar dem; han befriar dem från de ogudaktiga och frälsar dem, ty de taga sin tillflykt till honom.
En psalm av David; till åminnelse.
HERRE, straffa mig icke i din förtörnelse, och tukta mig icke i din vrede.
Ty dina pilar hava träffat mig, och din hand drabbar mig.
Det finnes intet helt på min kropp för din vredes skull, intet helbrägda i mina ben för min synds skull.
Ty mina missgärningar gå mig över huvudet; såsom en svår börda äro de mig för tunga.
Mina sår stinka och flyta för min dårskaps skull.
Jag går krokig och mycket lutande; hela dagen går jag sörjande.
Ty mina länder äro fulla av brand, och intet helt finnes på min kropp.
Jag är vanmäktig och illa sönderslagen; jag klagar för mitt hjärtas jämmers skull.
Herre, du känner all min trängtan, och min suckan är dig icke fördold.
Mitt hjärta slår häftigt, min kraft har övergivit mig; mina ögons ljus, också det är borta.
Mina vänner och fränder hålla sig fjärran ifrån min plåga, och mina närmaste hava ställt sig långt ifrån.
Snaror lägga de ut, som stå efter mitt liv, och de som söka min ofärd tala vad fördärvligt är; på svek tänka de hela dagen.
Men jag är lik en döv, som intet hör, och lik en stum, som icke upplåter sin mun;
ja, jag är lik en man som intet hör, och som icke har något gensvar i sin mun.
Se, på dig, HERRE, hoppas jag; du skall svara, Herre, min Gud.
Ty jag fruktar att de annars få glädja sig över mig, att de skola förhäva sig över mig, när min fot vacklar.
Ty jag är nära att falla, och min plåga är alltid inför mig;
ja, jag måste bekänna min missgärning, och jag sörjer över min synd.
Men mina fiender få leva och äro mäktiga, och många äro de som hata mig utan sak,
de som löna gott med ont, och som stå mig emot, därför att jag far efter det goda.
Övergiv mig icke, HERRE; min Gud, var icke långt ifrån mig.
Skynda till min hjälp, Herre, du min frälsning.
För sångmästaren, till Jedutun; en psalm av David.
Jag sade: »Jag vill akta på vad jag gör, så att jag icke syndar med min tunga; jag vill akta på att tygla min mun, så länge den ogudaktige är för mina ögon.»
Jag blev stum och tyst, jag teg i min sorg; man jag upprördes av smärta.
Mitt hjärta blev brinnande i mitt bröst: när jag begrundade, upptändes en eld i mig; jag talade med min tunga.
HERRE, lär mig betänka att jag måste få en ände, och vad som är mina dagars mått, så att jag förstår huru förgänglig jag är.
Se, såsom en handsbredd har du gjort mina dagars mått, och min livslängd är såsom intet inför dig; fåfänglighet allenast äro alla människor, huru säkra de än stå.
Sela.
Såsom en drömbild allenast gå de fram, fåfänglighet allenast är deras ävlan; de samla tillhopa och veta icke vem som skall få det.
Och nu, vad förbidar jag, Herre?
Till dig står mitt hopp.
Befria mig från alla mina överträdelser, låt mig icke bliva till smälek för dåren.
Jag tiger och upplåter icke min mun; ty det är du som har gjort det.
Vänd av ifrån mig din plåga; för din hands aga försmäktar jag.
Om du tuktar någon med näpst för missgärning, så är det ute med hans härlighet, såsom när mal krossas.
Fåfänglighet allenast äro alla människor.
Sela.
Hör min bön, o HERRE, och lyssna till mitt rop, tig icke vid mina tårar; ty jag är en främling i ditt hägn, en gäst såsom alla mina fäder.
Vänd ifrån mig din blick, så att jag får vederkvickas, innan jag går hädan och icke mer är till.
För sångmästaren; av David; en psalm.
Stadigt förbidade jag HERREN, och han böjde sig till mig och hörde mitt rop.
Han drog mig upp ur fördärvets grop, ur den djupa dyn; han ställde mina fötter på en klippa, han gjorde mina steg fasta;
han lade i min mun en ny sång, en lovsång till vår Gud.
Det skola många se och varda häpna, och skola förtrösta på HERREN.
Säll är den man som sätter sin förtröstan till HERREN; och icke vänder sig till dem som äro stolta och vika av i lögn.
Stora äro de under du har gjort, HERRE, min Gud, och de tankar du har tänkt för oss; dig är intet likt.
Jag ville förkunna dem och tala om dem, men de stå icke till att räkna.
Till slaktoffer och spisoffer har du icke behag -- öppna öron har du givit mig -- brännoffer och syndoffer begär du icke.
Därför säger jag: »Se, jag kommer; i bokrullen är skrivet vad jag skall göra.
Att göra din vilja, min Gud, är min lust, och din lag är i mitt hjärta.»
Jag bådar glädje, jag förkunnar din rättfärdighet i den stora församlingen; se, jag tillsluter icke mina läppar; du, HERRE, vet det.
Din rättfärdighet fördöljer jag icke i mitt hjärta, om din trohet och din frälsning talar jag; jag förtiger icke din nåd och din trofasthet för den stora församlingen.
Du, HERRE, skall icke tillsluta din barmhärtighet för mig; din nåd och din trofasthet må alltid bevara mig.
Ty lidanden omvärva mig, flera än jag kan räkna; mina missgärningar hava tagit mig fatt, så att jag icke kan se; de äro flera än håren på mitt huvud, och mitt mod har övergivit mig.
Värdes, o HERRE, rädda mig; HERRE, skynda till min hjälp.
Må alla de komma på skam och varda utskämda, som stå efter mitt liv för att förgöra det; må de vika tillbaka och blygas, som önska min ofärd.
Må de häpna i sin skam, som säga till mig: »Rätt så, rätt så!»
Men alla de som söka dig må fröjdas och vara glada i dig; de som åstunda din frälsning säge alltid: »Lovad vare HERREN!»
Är jag ock betryckt och fattig, Herren sörjer dock för mig.
Min hjälp och min befriare är du; min Gud, dröj icke.
För sångmästaren; en psalm av David.
Säll är den som låter sig vårda om den arme; honom skall HERREN hjälpa på olyckans dag.
HERREN skall bevara honom och behålla honom vid liv, han skall prisas säll i landet.
Icke skall du överlämna honom åt hans fienders vilja!
HERREN skall på sjukbädden stå honom bi; vid hans krankhet förvandlar du alldeles hans läger.
Så säger jag då: HERRE; var du mig nådig; hela du min själ, ty jag har syndat mot dig.
Mina fiender tala vad ont är mot mig: »När skall han dö och hans namn förgås?»
Kommer någon och besöker mig, så talar han falskhet; hans hjärta samlar åt honom vad ondskefullt är; sedan går han ut och talar därom.
De som hata mig tassla alla med varandra mot mig; de tänka ut mot mig det som är mig till skada.
»Ohjälplig ofärd har drabbat honom, han som ligger där skall icke mer stå upp.»
Ja, också min vän, som jag litade på, han som åt mitt bröd, lyfter nu mot mig sin häl.
Men du, HERRE, var mig nådig och upprätta mig, så vill jag vedergälla dem.
Att du har behag till mig, det vet jag därav att min fiende icke får jubla över mig.
Ty mig uppehåller du, för min ostrafflighets skull, och låter mig stå inför ditt ansikte evinnerligen. ----
Lovad vare HERREN, Israels Gud, från evighet till evighet!
Amen, Amen.
Andra boken
För sångmästaren; en sång av Koras söner.
Såsom hjorten trängtar till vattenbäckar, så trängtar min själ efter dig, o Gud.
Min själ törstar efter Gud, efter den levande Guden.
När skall jag få träda fram inför Guds ansikte?
Mina tårar äro min spis både dag och natt, ty ständigt säger man till mig: »Var är nu din Gud?»
Men jag vill utgjuta inom mig min själ och hava i minne huru jag gick med hopen upp till Guds hus, under fröjderop och tacksägelse, i högtidsskaran.
Varför är du så bedrövad, min själ, och så orolig i mig?
Hoppas på Gud; ty jag skall åter få tacka honom för frälsning genom honom.
Min Gud, bedrövad är min själ i mig; därför tänker jag på dig i Jordans land och på Hermons höjder, på Misars berg.
Djup ropar till djup, vid dånet av dina vattenfall; alla dina svallande böljor gå fram över mig.
Om dagen må HERREN beskära sin nåd, och om natten vill jag sjunga till hans ära och bedja till mitt livs Gud.
Jag vill säga till Gud, min klippa: »Varför har du förgätit mig, varför måste jag gå sörjande, trängd av fiender?»
Det är såsom krossade man benen i min kropp, när mina ovänner smäda mig, när de beständigt säga till mig: »Var är nu din Gud?»
Varför är du så bedrövad, min själ, och varför så orolig i mig?
Hoppas på Gud; ty jag skall åter få tacka honom, min frälsning och min Gud.
Skaffa mig rätt, o Gud, och utför min sak mot ett folk utan fromhet; rädda mig ifrån falska och orättfärdiga människor.
Ty du är den Gud som är mitt värn; varför har du förkastat mig?
Varför måste jag gå sörjande, trängd av fiender?
Sänd ditt ljus och din sanning; må de leda mig, må de föra mig till ditt heliga berg och till dina boningar,
så att jag får gå in till Guds altare, till Gud, som är min glädje och fröjd, och tacka dig på harpa, Gud, min Gud.
Varför är du så bedrövad, min själ, och varför så orolig i mig?
Hoppas på Gud; ty jag skall åter få tacka honom, min frälsning och min Gud.
För sångmästaren; av Koras söner; en sång.
Gud, med våra öron hava vi hört, våra fäder hava förtäljt därom för oss: om den gärning du gjorde i deras dagar, i forntidens dagar.
Det var du som med din hand utrotade hedningarna, men planterade dem; du fördärvade andra folk, men dem lät du utbreda sig.
Ty icke med sitt svärd intogo de landet, och deras egen arm gav dem icke seger, utan din högra hand och din arm och ditt ansiktes ljus, ty du hade behag till dem.
Du, densamme, är min konung, o Gud; så tillsäg nu Jakob seger.
Med din hjälp kunna vi stöta ned våra ovänner och i ditt namn förtrampa våra motståndare.
Ty icke på min båge förlitar jag mig, och mitt svärd kan icke giva mig seger;
nej, du giver oss seger över våra ovänner, och dem som hata oss låter du komma på skam.
Gud lova vi alltid, och ditt namn prisa vi evinnerligen.
Sela.
Och dock har du nu förkastat oss och låtit oss varda till blygd, och du drager icke ut med våra härar.
Du låter oss vika tillbaka för ovånnen, och de som hata oss taga sig byte.
Du låter oss bliva uppätna såsom får, och bland hedningarna han du förstrött oss.
Du säljer ditt folk för ett ringa pris, stor är icke den vinst du har gjort därpå.
Du låter oss bliva till smälek för våra grannar, till spott och hån för dem som bo omkring oss.
Du gör oss till ett ordspråk bland hedningarna, du låter folken skaka huvudet åt oss.
Hela dagen är min smälek inför mig, och blygsel höljer mitt ansikte,
när jag hör smädarens och lastarens tal, när jag ser fienden och den hämndgirige.
Allt detta har kommit över oss, och vi hava dock icke förgätit dig, ej heller svikit ditt förbund.
Våra hjärtan avföllo icke, och våra steg veko ej av ifrån din väg,
så att du därför har krossat oss i schakalers land och övertäckt oss med dödsskugga.
Om vi hade förgätit vår Guds namn och uträckt våra händer till en främmande gud,
månne icke Gud skulle hava utrannsakat det, han som känner hjärtats lönnligheter?
Nej, för din skull varda vi dödade hela dagen och bliva aktade såsom slaktfår.
Vakna upp; varför sover du, Herre?
Vakna, förkasta oss icke för alltid.
Varför döljer du ditt ansikte och förgäter vårt lidande och trångmål?
Se, vår själ är nedböjd i stoftet, vår kropp ligger nedtryckt till jorden.
Stå upp till vår hjälp, och förlossa oss för din nåds skull.
För sångmästaren, efter »Liljor»; av Koras söner; en sång, ett kväde om kärlek.
Mitt hjärta flödar över av sköna ord; jag säger: min dikt gäller en konung; en snabb skrivares penna är min tunga.
Du är den skönaste bland människors barn, ljuvlighet är utgjuten över dina läppar; så se vi att Gud har välsignat dig evinnerligen.
Omgjorda din länd med ditt svärd, du hjälte, i ditt majestät och din härlighet.
Och drag så åstad, lyckosam i din härlighet, till försvar för sanning, för ödmjukhet och rättfärdighet, så skall din högra hand lära dig underbara gärningar.
Skarpa äro dina pilar; folk skola falla för dig; konungens fiender skola träffas i hjärtat.
Gud, din tron förbliver alltid och evinnerligen; ditt rikes spira är rättvisans spira.
Du älskar rättfärdighet och hatar orättfärdighet; därför har Gud, din Gud, smort dig med glädjens olja mer än dina medbröder.
Av myrra, aloe och kassia dofta alla dina kläder; från elfenbenspalatser gläder dig strängaspel.
Konungadöttrar har du såsom tärnor i ditt hov, en drottning står vid din högra sida, i guld från Ofir.
Hör, dotter, och giv akt, och böj ditt öra härtill: Förgät nu ditt folk och din faders hus,
och må konungen få hava sin lust i din skönhet; ty han är din herre, och för honom skall du falla ned.
Se, dottern Tyrus, ja, de rikaste folk söka nu att vinna din ynnest med skänker.
Idel härlighet är hon, konungadottern i gemaket: av guldvirkat tyg består hennes dräkt,
i brokigt vävda kläder föres hon till konungen; jungfrur, hennes väninnor, följa henne åt; de ledas in till dig.
Under glädje och fröjd föras de fram, de tåga in i konungens palats.
I dina fäders ställe skola dina söner träda; dem skall du sätta till furstar överallt i landet.
Ditt namn vill jag göra prisat bland alla kommande släkten; så skola ock folken lova dig, alltid och evinnerligen.
För sångmästaren; av Koras söner; till Alamót; en sång.
Gud är vår tillflykt och vår starkhet, en hjälp i nöden, väl beprövad.
Därför skulle vi icke frukta, om än jorden omvälvdes och bergen vacklade ned i havsdjupet;
om än dess vågor brusade och svallade, så att bergen bävade vid dess uppror.
Sela.
En ström går fram, vars flöden giva glädje åt Guds stad, åt den Högstes heliga boning.
Gud bor därinne, den vacklar icke; Gud hjälper den, när morgonen gryr.
Hedningarna larma, riken vackla; han låter höra sin röst, då försmälter jorden.
HERREN Sebaot är med oss, Jakobs Gud är vår borg.
Sela.
Kommen och skåden HERRENS verk: gärningar som väcka häpnad gör han på jorden.
Han stillar strider intill jordens ända, bågen bryter han sönder och bräcker spjutet, i eld bränner han upp stridsvagnarna.
»Bliven stilla och besinnen att jag är Gud; hög varder jag bland hedningarna, hög på jorden.»
HERREN Sebaot är men oss, Jakobs Gud är vår borg.
Sela.
För sångmästaren; av Koras söner; en psalm.
Klappen i händerna, alla folk, höjen jubel till Gud med fröjderop.
Ty HERREN är den Högste, fruktansvärd är han, en stor konung över hela jorden.
Han tvingar folk under oss och folkslag under våra fötter.
Han utväljer åt oss vår arvedel, Jakobs, hans älskades, stolthet.
Sela.
Gud har farit upp under jubel, HERREN, under basuners ljud.
Lovsjungen Gud, lovsjungen; lovsjungen vår konung, lovsjungen.
Ty Gud är konung över hela jorden; lovsjungen honom med en sång.
Gud är nu konung över hedningarna, Gud har satt sig på sin heliga tron.
Folkens ypperste hava församlat sig till att bliva ett Abrahams Guds folk.
Ty Gud tillhöra de som äro jordens sköldar; högt är han upphöjd.
En sång, en psalm av Koras söner.
Stor är HERREN och högt lovad, i vår Guds stad, på sitt heliga berg.
Skönt höjer det sig, hela jordens fröjd, berget Sion längst uppe i norr, den store konungens stad.
Gud har i dess palatser gjort sig känd såsom ett värn.
Ty se, konungarna församlade sig, tillhopa drogo de fram.
De sågo det, då häpnade de; de förskräcktes, de flydde.
Bävan grep dem där, ångest lik en barnaföderskas.
Så krossar du Tarsis-skepp med östanvinden.
Såsom vi hade hört, så fingo vi se det, i HERREN Sebaots stad, i vår Guds stad; Gud håller den vid makt till evig tid.
Sela.
Vi tänka, o Gud, på din nåd, när vi stå i ditt tempel.
Såsom ditt namn, o Gud, så når ock ditt lov intill jordens ändar; din högra hand är full av rättfärdighet.
Sions berg glädje sig, Juda döttrar fröjde sig, för dina domars skull.
Gån omkring Sion och vandren runt därom, räknen dess torn;
given akt på dess murar, skriden genom dess palatser, så att I kunnen förtälja därom för ett kommande släkte.
Ty sådan är Gud, vår Gud, alltid och evinnerligen; intill döden skall han ledsaga oss.
För sångmästaren; av Koras söner; en psalm.
Hören detta, alla folk, lyssnen härtill, I alla som leven i världen,
både låga och höga, rika såväl som fattiga.
Hin mun skall tala visdom, och mitt hjärtas tanke skall vara förstånd.
Jag vill böja mitt öra till lärorikt tal, jag vill yppa vid harpan min förborgade kunskap.
Varför skulle jag frukta i olyckans dagar, när mina förföljares ondska omgiver mig?
De förlita sig på sina ägodelar och berömma sig av sin stora rikedom.
Men sin broder kan ingen förlossa eller giva Gud lösepenning för honom.
För dyr är lösen för hans själ och kan icke betalas till evig tid,
så att han skulle få leva för alltid och undgå att se graven.
Nej, man skall se att visa män dö, att dårar och oförnuftiga förgås likasom de; de måste lämna sina ägodelar åt andra.
De tänka att deras hus skola bestå evinnerligen, deras boningar från släkte till släkte; de uppkalla jordagods efter sina namn.
Men en människa har, mitt i sin härlighet, intet bestånd, hon är lik fänaden, som förgöres.
Den vägen gå de, dårar som de äro, och de följas av andra som finna behag i deras tal.
Sela.
Såsom en fårhjord drivas de ned till dödsriket, där döden bliver deras herde.
Så få de redliga makt över dem, när morgonen gryr, medan deras skepnader förtäras av dödsriket och ej få annan boning.
Men min själ skall Gud förlossa ifrån dödsrikets våld, ty han skall upptaga mig.
Sela.
Frukta icke, när en man bliver rik, när hans hus växer till i härlighet.
Ty av allt detta får han vid sin död intet med sig, och hans härlighet följer honom icke ditned.
Om han ock prisar sig välsignad under sitt liv, ja, om man än berömmer dig, när du gör goda dagar, så skall dock vars och ens själ gå till hans fäders släkte, till dem som aldrig mer se ljuset.
En människa som, mitt i sin härlighet, är utan förstånd, hon är lik fänaden, som förgöres.
En psalm av Asaf.
Gud, HERREN Gud, talar och kallar jorden, allt mellan öster och väster.
Från Sion, skönhetens fullhet, träder Gud fram i glans.
Vår Gud kommer, och han skall icke tiga.
Förtärande eld går framför honom, och omkring honom stormar det med makt.
Han kallar på himmelen därovan och på jorden, för att döma sitt folk:
»Församlen till mig mina fromma, som sluta förbund med mig vid offer.»
Och himlarna förkunna att han är rättfärdig, att Gud är den som skipar rätt.
Sela.
Hör, mitt folk, jag vill tala; Israel, låt mig varna dig.
Gud, din Gud, är jag.
Icke för dina slaktoffer vill jag gå till rätta med dig; dina brännoffer har jag alltid inför mig.
Jag vill icke taga tjurar ur ditt hus eller bockar ur dina fållor;
ty mina äro alla skogens djur, boskapen på de tusende bergen;
jag känner alla fåglar på bergen, och vad som rör sig på marken är mig bekant.
Om jag hungrade, skulle jag icke säga dig det; ty min är jordens krets med allt vad därpå är.
Skulle jag äta tjurars kött, och skulle jag dricka bockars blod?
Nej, offra lovets offer åt Gud, så skall du få infria dina löften till den Högste.
Och åkalla mig i nöden, så vill jag hjälpa dig, och du skall prisa mig.»
Men till den ogudaktige säger Gud: »Huru kan du tala om mina stadgar och föra mitt förbund på tungan,
du som hatar tuktan och kastar mina ord bakom dig?
Om du ser en tjuv, så håller du med honom, och med äktenskapsbrytare giver du dig i lag.
Din mun släpper du lös till vad ont är, och din tunga hopspinner svek.
Du sitter där och förtalar din broder, din moders son lastar du!
Så gör du, och jag tiger, och nu tror du att jag är såsom du.
Nej, jag vill straffa dig och ställa dig det för ögonen.
I som förgäten Gud, märken detta, för att jag icke må sönderriva eder utan räddning:
den som offrar lovets offer, han ärar mig; och den som aktar på sin väg, honom skall jag låta se Guds frälsning.»
För sångmästaren; en psalm av David,
när profeten Natan kom till honom, då han hade gått in till Bat-Seba.
Gud, var mig nådig efter din godhet, utplåna mina överträdelser efter din stora barmhärtighet.
Två mig väl från min missgärning, och rena mig från synd.
Ty jag känner mina överträdelser, och min synd är alltid inför mig.
Mot dig allena har jag syndat och gjort vad ont är i dina ögon; på det att du må finnas rättfärdig i dina ord och rättvis i dina domar.
Se, i synd är jag född, och i synd har min moder avlat mig.
Du har ju behag till sanning i hjärtegrunden; så lär mig då vishet i mitt innersta.
Skära mig med isop, så att jag varder ren; två mig, så att jag bliver vitare än snö.
Låt mig förnimma fröjd och glädje, låt de ben som du har krossat få fröjda sig.
Vänd bort ditt ansikte från mina synder, och utplåna alla mina missgärningar.
Skapa i mig, Gud, ett rent hjärta, och giv mig på nytt en frimodig ande.
Förkasta mig icke från ditt ansikte, och tag icke din helige Ande ifrån mig.
Låt mig åter få fröjdas över din frälsning, och uppehåll mig med villighetens ande.
Då skall jag lära överträdarna dina vägar, och syndarna skola omvända sig till dig.
Rädda mig undan blodstider, Gud, du min frälsnings Gud, så skall min tunga jubla över din rättfärdighet.
Herre, upplåt mina läppar, så att min mun kan förkunna ditt lov.
Ty du har icke behag till offer, eljest skulle jag giva dig sådana; till brännoffer har du icke lust.
Det offer som behagar Gud är en förkrossad ande; ett förkrossat och bedrövat hjärta skall du, Gud, icke förakta.
Gör väl mot Sion i din nåd, bygg upp Jerusalems murar.
Då skall du undfå rätta offer, som behaga dig, brännoffer och heloffer; då skall man offra tjurar på ditt altare.
För sångmästaren; en sång av David,
när edoméen Doeg kom och berättade för Saul och sade till honom: »David har gått in i Ahimeleks hus.»
Varför berömmer du dig av vad ont är, du våldsverkare?
Guds nåd varar ju beständigt.
Din tunga far efter fördärv, den är lik en skarp rakkniv, du arglistige.
Du älskar ont mer än gott, lögn mer än att tala vad rätt är.
Sela.
Ja, du älskar allt fördärvligt tal, du falska tunga.
Därför skall ock Gud störta dig ned för alltid, han skall gripa dig och rycka dig ut ur din hydda och utrota dig ur de levandes land.
Sela.
Och de rättfärdiga skola se det och frukta, de skola le åt honom:
»Se där är den man som icke gjorde Gud till sitt värn, utan förlitade sig på sin stora rikedom, trotsig i sin lystnad!»
Men jag skall vara såsom ett grönskande olivträd i Guds hus; jag förtröstar på Guds nåd alltid och evinnerligen.
Jag skall evinnerligen tacka dig för att du har gjort det; och inför dina fromma skall jag förbida ditt namn, ty det är gott.
För sångmästaren, till Mahalát; en sång av David.
Dårarna säga i sina hjärtan: »Det finnes ingen Gud.»
Fördärv och styggelse är deras onda verk; ingen finnes, som gör vad gott är.
Gud skådar ned från himmelen på människors barn, för att se om det finnes någon förståndig, någon som söker Gud.
Nej, alla hava de avfallit, allasammans äro de fördärvade; ingen finnes, som gör vad gott är, det finnes icke en enda.
Hava de då intet fått förnimma, dessa ogärningsmän, dessa som uppäta mitt folk, likasom åte de bröd, och som icke åkalla Gud?
Jo, där överföll dem förskräckelse, varest intet förskräckligt var; ty Gud förströdde deras ben, när de lägrade sig mot dig.
Så lät du dem komma på skam, ja, Gud förkastade dem.
Ack att från Sion komme frälsning för Israel!
När Gud vill åter upprätta sitt folk, då skall Jakob fröjda sig, då skall Israel vara glad.
För sångmästaren, med strängaspel; en sång av David,
när sifiterna kommo och sade till Saul: »David håller sig nu gömd hos oss.»
Gud, fräls mig genom ditt namn, och skaffa mig rätt genom din makt.
Gud, hör min bön, lyssna till min muns tal.
Ty främlingar resa sig upp mot mig, och våldsverkare stå efter mitt liv; de hava icke Gud för ögonen.
Sela.
Se, Gud är min hjälpare, Herren uppehåller min själ.
Må det onda falla tillbaka på mina förföljare, förgör dem, du som är trofast.
Då skall jag offra åt dig med villigt hjärta; jag skall prisa ditt namn, o HERRE, ty det är gott.
Ja, ur all nöd räddar det mig, och mitt öga får se med lust på mina fiender.
För sångmästaren, med strängaspel; en sång av David.
Lyssna, Gud, till min bön, och fördölj dig icke för min åkallan.
Akta på mig och svara mig.
I mitt bekymmer är jag utan ro och måste klaga,
vid fiendens rop, vid den ogudaktiges skri.
Ty de vilja draga fördärv över mig, och i vrede ansätta de mig.
Mitt hjärta ängslas i mitt bröst, och dödens fasor hava fallit över mig.
Fruktan och bävan kommer över mig, och förfäran övertäcker mig.
Därför säger jag: Ack att jag hade vingar såsom duvan!
Då skulle jag flyga bort och söka mig ett bo.
Ja, långt bort skulle jag fly, jag skulle taga härbärge i öknen.
Sela.
Jag skulle skynda att söka mig en tillflykt undan stormvind och oväder.
Fördärva dem, Herre; gör deras tungor oense.
Ty våld och genstridighet ser jag i staden.
Dag och natt gå de omkring den, ovanpå dess murar, ondska och olycka råda därinne;
ja, fördärv råder därinne, och från dess torg vika icke förtryck och svek.
Se, det är icke en fiende som smädar mig, det kunde jag fördraga; det är icke min ovän som förhäver sig mot mig, för honom kunde jag gömma mig undan.
Nej, du gör det, du som var min jämlike, min vän och förtrogne,
du som levde med mig i ljuvlig förtrolighet, du som i Guds hus gick med mig i högtidsskaran.
Döden komme över dem oförtänkt, levande fare de ned i dödsriket; ty ondska råder i deras boning, i deras hjärtan.
Men jag ropar till Gud; HERREN skall frälsa mig.
Afton och morgon och middag vill jag utgjuta mitt bekymmer och klaga, och han skall höra min röst.
Han förlossar min själ och skaffar henne ro, så att de icke komma vid mig; ty de äro många, som stå mig emot.
Gud skall höra det och giva dem svar, han som sitter på sin tron av ålder.
Sela.
Ty de vilja icke ändra sig, och de frukta ej Gud.
Den mannen bär händer på sin vän; han bryter sitt förbund.
Orden i hans mun äro hala såsom smör, men stridslust fyller hans hjärta; hans ord äro lenare än olja, dock äro de dragna svärd.
Kasta din börda på HERREN, han skall uppehålla dig; han skall i evighet icke tillstädja att den rättfärdige vacklar.
Gud, du skall störta dem ned i gravens djup; de blodgiriga och falska skola ej nå sin halva ålder.
Men jag förtröstar på dig.
För sångmästaren, efter »Den stumma duvan i fjärran»; en sång av David, når filistéerna grepo honom i Gat.
Var mig nådig, o Gud, ty människor stå mig efter livet; beständigt tränga mig stridsmän.
Mina förföljare stå mig beständigt efter livet; ja, de äro många, som i högmod strida mot mig.
Men när fruktan kommer över mig, sätter jag min förtröstan på dig.
Med Guds hjälp skall jag få prisa hans ord, på Gud förtröstar jag och skall icke frukta; vad kan det som är kött göra mig?
Beständigt förbittra de livet för mig, alla deras tankar gå ut på att skada mig.
De rota sig samman, de lägga försåt, de vakta på mina steg, ty de stå efter mitt liv.
Skulle de räddas med all sin ondska?
Nej, slå ned folken, Gud, i din vrede.
Du har räknat min flykts dagar.
Samla mina tårar i din lägel; de stå ju i din bok.
Så måste då mina fiender vika tillbaka på den dag då jag ropar; det vet jag, att Gud står mig bi.
Med Guds hjälp skall jag få prisa hans ord; med HERRENS hjälp skall jag få prisa hans ord.
På Gud förtröstar jag och skall icke frukta; vad kunna människor göra mig?
Jag har löften att infria till dig, o Gud; jag vill betala dig lovoffer.
Ty du har räddat min själ från döden, ja, mina fötter ifrån fall, så att jag kan vandra inför Gud i de levandes ljus.
För sångmästaren; »Fördärva icke»; en sång av David, när han flydde för Saul och var i grottan.
Var mig nådig, o Gud, var mig nådig; ty till dig tager min själ sin tillflykt.
Ja, under dina vingars skugga vill jag taga min tillflykt, till dess att det onda är förbi.
Jag ropar till Gud den Högste, till Gud, som fullbordar sitt verk för mig.
Han skall sända från himmelen och frälsa mig, när jag smädas av människor som stå mig efter livet.
Sela.
Gud skall sända sin nåd och sin trofasthet.
Min själ är omgiven av lejon, jag måste ligga bland eldsprutare, bland människor vilkas tänder äro spjut och pilar, och vilkas tungor äro skarpa svärd.
Upphöjd vare du, Gud, över himmelen; över hela jorden sträcke sig din ära.
De lägga ut nät för mina fötter, min själ böjes ned, de gräva för mig en grop, men de falla själva däri.
Sela.
Mitt hjärta är frimodigt, o Gud, mitt hjärta är frimodigt; jag vill sjunga och lova.
Vakna upp, min ära; upp, psaltare och harpa!
Jag vill väcka morgonrodnaden.
Jag vill tacka dig bland folken, Herre; jag vill lovsjunga dig bland folkslagen.
Ty din nåd är stor allt upp till himmelen och din trofasthet allt upp till skyarna.
Upphöjd vare du, Gud, över himmelen; över hela jorden sträcke sig din ära.
För sångmästaren; »Fördärva icke»; av David; en sång.
Talen I väl i eder stumhet vad rättfärdigt är?
Dömen I såsom rätt är, I människors barn?
Nej, i hjärtat uppgören I onda anslag; I vägen ut i landet edra händers våld.
De ogudaktiga äro avfälliga allt ifrån modersskötet; de lögnaktiga fara vilse ända från sin moders liv.
Gift är i dem, likt ormens gift; en döv huggorm likna de, en som tillstoppar sitt öra,
så att han icke hör tjusarnas röst, icke den förfarne besvärjarens.
Gud, krossa tänderna i deras mun; bryt ut, o HERRE, de unga lejonens kindtänder.
Låt dem bliva till intet, likasom vatten som förrinner.
När någon skjuter sina pilar, blive de såsom utan udd.
Må han vara lik snigeln, som upplöses och förgås, lik en kvinnas foster, som ej fick skåda solen.
Förrän edra grytor hava hunnit märka bränslet, och medan köttet ännu är rått, skall en glödvind rycka bort det.
Den rättfärdige skall glädja sig, när han skådar hämnden, han skall två sina fötter i den ogudaktiges blod.
Och människorna skola säga: »Ja, den rättfärdige får sin lön; ja, det finnes en Gud som dömer på jorden.»
För sångmästaren; »Fördärva icke»; en sång av David, när Saul sände och lät bevaka hans hus för att döda honom.
Rädda mig, min Gud, från mina fiender, beskydda mig för mina motståndare.
Rädda mig från ogärningsmännen, och fräls mig från de blodgiriga.
Ty se, de ligga i försåt för mig; grymma människor rota sig samman mot mig, utan någon min överträdelse eller synd, o HERRE.
Utan någon min missgärning löpa de fram och göra sig redo; vakna upp, kom mig till mötes, och se härtill.
Ja, du HERRE Gud Sebaot, Israels Gud, vakna och hemsök alla hedningar, hemsök utan nåd alla trolösa ogärningsmän.
Sela.
Var afton komma de tillbaka, de tjuta såsom hundar och stryka omkring i staden.
Se, deras mun flödar över, svärd äro på deras läppar, ty »vem skulle höra det?»
Men du, HERRE, ler åt dem; du bespottar alla hedningar.
Mot deras makt vill jag hålla mig till dig, ty Gud är min borg.
Min Gud kommer mig till mötes med sin nåd, Gud låter mig se med lust på mina förföljare.
Dräp dem icke, på det att mitt folk ej må förgäta det; låt dem genom din kraft driva ostadiga omkring, och slå dem ned, du vår sköld, o Herre.
Vart ord på deras läppar är en synd i deras mun.
Må de fångas i sitt högmod, genom den förbannelse och lögn som de tala.
Förgör dem i vrede, förgör dem, så att de ej mer äro till; och må de förnimma att det är Gud som råder i Jakob, allt intill jordens ändar.
Sela.
Ja, var afton komma de tillbaka, de tjuta såsom hundar och stryka omkring i staden.
De driva omkring efter rov; om de icke bliva mätta, så stanna de kvar över natten.
Men jag vill sjunga om din makt och jubla var morgon över din nåd; ty du var för mig en borg och en tillflykt, när jag var i nöd.
Min starkhet, dig vill jag lovsjunga, ty Gud är min borg, min nåderike Gud.
För sångmästaren, efter »Vittnesbördets lilja»; en sång, till att inläras; av David,
när han var i fejd med Aram-Naharaim och Aram-Soba, och Joab kom tillbaka och slog edoméerna i Saltdalen, tolv tusen man.
Gud, du har förkastat och förskingrat oss, du har varit vred; upprätta oss igen.
Du har kommit jorden att bäva och rämna; hela nu dess revor, ty den vacklar.
Du har låtit ditt folk se hårda ting, du har iskänkt åt oss rusande vin.
Men åt dem som frukta dig gav du ett baner, dit de kunde samla sig för att undfly bågen.
Sela.
På det att dina vänner må varda räddade, må du giva seger med din högra hand och bönhöra oss.
Gud har talat i sin helgedom: »Jag skall triumfera, jag skall utskifta Sikem och skall avmäta Suckots dal.
Mitt är Gilead, och mitt är Manasse, Efraim är mitt huvuds värn, Juda min härskarstav;
Moab är mitt tvagningskärl, på Edom kastar jag min sko; höj jubelrop till min ära, du filistéernas land.»
Vem skall föra mig till den fasta staden, vem leder mig till Edom?
Har icke du, o Gud, förkastat oss, så att du ej drager ut med våra härar, o Gud?
Giv oss hjälp mot ovännen; ty människors hjälp är fåfänglighet.
Med Gud kunna vi göra mäktiga ting; han skall förtrampa våra ovänner.
För sångmästaren, till strängaspel; av David.
Hör, o Gud, mitt rop, akta på min bön.
Från jordens ända ropar jag till dig, ty mitt hjärta försmäktar; för mig upp på en klippa, som är mig alltför hög.
Ty du är min tillflykt, ett starkt torn mot fienden.
Låt mig bo i din hydda evinnerligen; under dina vingars beskärm tager jag min tillflykt.
Sela.
Ty du, o Gud, hör mina löften, åt dem som frukta ditt namn giver du en arvedel.
Du förökar konungens dagar; hans år skola vara från släkte till släkte.
Må han sitta på sin tron inför Gud evinnerligen; låt nåd och trofasthet bevara honom.
Då skall jag lovsjunga ditt namn till evig tid, i det jag får infria mina löften dag efter dag.
För sångmästaren, till Jedutun; en psalm av David.
Allenast hos Gud söker min själ sin ro; från honom kommer min frälsning.
Allenast han är min klippa och min frälsning, min borg, jag skall ej mycket vackla.
Huru länge viljen I rasa mot denne man, samfällt slå honom ned, såsom vore han en lutande vägg, en sönderbräckt mur?
De rådslå allenast om att stöta honom ned från hans höjd, de hava behag till lögn; med munnen välsigna de, men i sitt innersta förbanna de.
Sela.
Allenast i Gud må du hava din ro, min själ; ty från honom kommer mitt hopp.
Allenast han är min klippa och min frälsning, min borg, jag skall icke vackla.
Hos Gud är min frälsning och min ära; min starka klippa, min tillflykt har jag i Gud.
Förtrösta på honom alltid, du folk; utgjuten för honom edra hjärtan.
Gud är vår tillflykt.
Sela.
Allenast ett intet äro människors barn, myndiga herrar fåfänglighet; i vågskålen äro de för lätta, mindre än intet äro de allasammans.
Förliten eder icke på orätt vinning, sätten icke ett fåfängligt hopp till rov: om ock eder rikedom växer, så akten icke därpå.
En gång har Gud sagt det, ja, två gånger har jag hört det, att hos Gud är makten;
och hos dig, Herre, är nåd.
Ty du vedergäller var och en efter hans gärningar.
En psalm av David, när han var i Juda öken.
Gud, du är min Gud, bittida söker jag dig; min själ törstar efter dig, min kropp längtar efter dig, i ett torrt land, som försmäktar utan vatten.
Så skådar jag nu efter dig i helgedomen, för att få se din makt och ära.
Ty din nåd är bättre än liv; mina läppar skola prisa dig.
Så skall jag då lova dig, så länge jag lever; i ditt namn skall jag upplyfta mina händer.
Min själ varder mättad såsom av märg och fett; och med jublande läppar lovsjunger min mun,
när jag kommer ihåg dig på mitt läger och under nattens väkter tänker på dig.
Ty du är min hjälp, och under dina vingars skumma jublar jag.
Min själ håller sig intill dig; din högra hand uppehåller mig.
Men dessa som stå efter mitt liv och vilja fördärva det, de skola fara ned i jordens djup.
De skola givas till pris åt svärdet, rovdjurs byte skola de varda.
Men konungen skall glädja sig i Gud; berömma sig skall var och en som svär vid honom, ty de lögnaktigas mun skall varda tillstoppad.
För sångmästaren; en psalm av David.
Hör, o Gud, min röst, när jag klagar, bevara mitt liv, ty fienden förskräcker mig.
Fördölj mig för de ondas hemliga råd, för ogärningsmännens larmande hop;
ty de vässa sina tungor likasom svärd, med bittra ord lägga de an såsom med pilar,
för att i lönndom skjuta den ostrafflige; plötsligt skjuta de på honom, utan försyn.
De befästa sig i sitt onda uppsåt, de orda om huru de skola lägga ut snaror; de säga: »Vem skulle se oss?»
De tänka ut onda anslag: »Nu äro vi redo med det råd vi hava uttänkt!»
Ja, djupa äro männens tankar och hjärtan.
Då skjuter Gud dem; plötsligt sårar dem hans pil.
De bringas på fall och få straff för sina tungors skull; var och en som ser dem rister huvudet.
Och alla människor varda förskräckta; de förkunna vad Gud har gjort och förstå hans verk.
Den rättfärdige skall glädja sig i HERREN och taga sin tillflykt till honom, och alla rättsinniga skola berömma sig.
För sångmästaren; en psalm; en sång av David.
Gud, dig lovar man i stillhet i Sion, och till dig får man infria löfte.
Du som hör bön, till dig kommer allt kött.
Mina missgärningar voro mig övermäktiga; men du förlåter våra överträdelser.
Säll är den som du utväljer och låter komma till dig, så att han får bo i dina gårdar.
Må vi få mätta oss med det goda i ditt hus, det heliga i ditt tempel.
Med underbara gärningar bönhör du oss i rättfärdighet, du vår frälsnings Gud, du som är en tillflykt för alla jordens ändar och för havet i fjärran;
du som gör bergen fasta genom din kraft, ty du är omgjordad med makt;
du som stillar havens brus, deras böljors brus och folkens larm.
De som bo vid jordens ändar häpna för dina tecken; österland och västerland uppfyller du med jubel.
Du låter dig vårda om landet och giver det överflöd, rikedom i ymnigt mått; Guds källa har vatten till fyllest.
Du bereder säd åt människorna, när du så bereder jorden.
Dess fåror vattnar du, du jämnar det som är upplöjt; med regnskurar uppmjukar du den, det som växer därpå välsignar du.
Du kröner året med ditt goda, och dina spår drypa av fetma.
Betesmarkerna i öknen drypa, och höjderna omgjorda sig med fröjd.
Ängarna hölja sig i hjordar, och dalarna betäckas med säd; man höjer jubelrop och sjunger.
För sångmästaren; en sång, en psalm.
Höjen jubel till Gud, alla länder;
lovsjungen hans namns ära, given honom ära och pris.
Sägen till Gud: Huru underbara äro icke dina gärningar!
För din stora makts skull visa dina fiender dig underdånighet.
Alla länder skola tillbedja och lovsjunga dig; de skola lovsjunga ditt namn.
Sela.
Kommen och sen vad Gud har gjort; underbara äro hans gärningar mot människors barn.
Han förvandlade havet till torrt land; till fots gingo de genom floden; då gladdes vi över honom.
Genom sin makt råder han evinnerligen, hans ögon giva akt på hedningarna; de gensträviga må icke förhäva sig.
Sela.
Prisen, I folk, vår Gud, och låten hans lov ljuda högt;
ty han har beskärt liv åt vår själ och har icke låtit vår fot vackla.
Ty väl prövade de oss, o Gud, du luttrade oss, såsom silver luttras;
du förde oss in i fängelse, du lade en tung börda på vår rygg;
du lät människor fara fram över vårt huvud, vi måste gå genom eld och vatten.
Men du har fört oss ut och vederkvickt oss.
Så kommer jag då till ditt hus med brännoffer, jag vill infria mina löften till dig,
dem till vilka mina låppar öppnade sig, och som min mun uttalade i min nöd.
Brännoffer av feta får vill jag frambära åt dig, med offerånga av vädurar; jag vill offra både tjurar och bockar.
Sela.
Kommen och hören, så vill jag förtälja för eder, I alla som frukten Gud, vad han har gjort mot min själ.
Till honom ropade jag med min mun, och lovsång var redan på min tunga.
Om jag hade förehaft något orätt i mitt hjärta, så skulle Herren icke höra mig.
Men Gud har hört mig, han har aktat på mitt bönerop.
Lovad vare Gud, som icke har förkastat min bön eller vänt ifrån mig sin nåd!
För sångmästaren, med strängaspel; en psalm, en sång.
Gud vare oss nådig och välsigne oss, han låte sitt ansikte lysa och ledsaga oss, Sela,
för att man på jorden må känna din väg, bland alla hedningar din frälsning.
Folken tacke dig, o Gud, alla folk tacke dig.
Folkslagen glädje sig och juble, ty du dömer folken rätt, och du leder folkslagen på jorden.
Sela.
Folken tacke dig, o Gud, alla folk tacke dig.
Jorden har givit sin gröda.
Gud, vår Gud, välsigne oss.
Gud välsigne oss, och alla jordens ändar frukte honom.
För sångmästaren; av David; en psalm, en sång.
Gud står upp; hans fiender varda förskingrade, och de som hata honom fly för hans ansikte.
Såsom rök fördrives, så fördrivas de av dig; likasom vaxet smälter för eld, så förgås de ogudaktiga för Guds ansikte.
Men de rättfärdiga äro glada, de fröjda sig inför Gud och jubla i glädje.
Sjungen till Guds ära, lovsägen hans namn.
Gören väg för honom som drager fram genom öknarna.
Hans namn är HERREN, fröjdens inför honom;
de faderlösas fader och änkors försvarare, Gud i sin heliga boning,
en Gud som förhjälper de ensamma till ett hem, och som för de fångna ut till lycka; allenast de gensträviga måste bo i en öken.
Gud, när du drog ut i spetsen för ditt folk, när du gick fram i ödemarken, Sela,
då bävade jorden, då utgöt himmelen sina flöden inför Guds ansikte; ja, Sinai bävade för Guds ansikte; Israels Guds.
Ett nåderikt regn lät du falla, o Gud; ditt arvland, som försmäktade, vederkvickte du.
Din skara fick bo däri; genom din godhet beredde du det åt de betryckta, o Gud.
Herren låter höra sitt ord, stor är skaran av kvinnor som båda glädje:
»Härskarornas konungar fly, de fly, och husmodern därhemma får utskifta byte.
Viljen I då ligga stilla inom edra hägnader?
Duvans vingar äro höljda i silver, och hennes fjädrar skimra av guld.
När den Allsmäktige förströr konungarna i landet, faller snö på Salmon.»
Ett Guds berg är Basans berg, ett högtoppigt berg är Basans berg.
Men varför sen I så avogt, I höga berg, på det berg som Gud har utkorat till sitt säte, det där ock HERREN skall bo för alltid?
Guds vagnar äro tiotusenden, tusen och åter tusen; Herren drog fram med dem, Sinai är nu i helgedomen.
Du for upp i höjden, du tog fångar, du undfick gåvor bland människorna, ja, också de gensträviga skola bo hos HERREN Gud.
Lovad vare Herren!
Dag efter dag bär han oss; Gud är vår frälsning.
Sela.
Gud är för oss en Gud som frälsar, och hos HERREN, Herren finnes räddning från döden.
Men Gud sönderkrossar sina fienders huvuden, krossar hjässan på den som går där med skuld.
Herren säger: »Från Basan skall jag hämta dem, från havets djup skall jag hämta dem upp,
så att du kan stampa med din fot i blod och låta dina hundars tunga få sin del av fienderna.»
Man ser, o Gud, ditt högtidståg, min Guds, min konungs, tåg inne i helgedomen.
Främst gå sångare, harpospelare följa efter, mitt ibland unga kvinnor som slå på pukor.
Lova Gud i församlingarna, loven Herren, I av Israels brunn.
Där går Benjamin, den yngste, han för dem an; där går skaran av Juda furstar, Sebulons furstar, Naftalis furstar.
Din Gud har beskärt dig makt; så håll nu vid makt, o Gud, vad du har gjort för oss.
I ditt tempel i Jerusalem bäre konungar fram sina skänker åt dig.
Näps odjuret i vassen, tjurarnas hop med deras kalvar, folken, må de ödmjukt hylla dig med sina silverstycken.
Ja, han förströr de folk som finna behag i krig.
De mäktige skola komma hit från Egypten, Etiopien skall skynda hit till Gud, med gåvor i händerna.
I riken på jorden, sjungen till Guds ära; lovsägen Herren, Sela,
honom som far fram på urtidshimlarnas himmel.
Ja, där låter han höra sin röst, en mäktig röst.
Given Gud makten; över Israel är hans härlighet, och hans makt är i skyarna.
Fruktansvärd är du, Gud, i din helgedom; Israels Gud, han giver makt och styrka åt sitt folk.
Lovad vare Gud!
För sångmästaren, efter »Liljor»; av David.
Fräls mig, Gud; ty vattnen tränga mig inpå livet.
Jag har sjunkit ned i djup dy, där ingen botten är; jag har kommit i djupa vatten, och svallet vill fördränka mig.
Jag har ropat mig trött, min strupe är förtorkad; mina ögon försmäkta av förbidan efter min Gud.
Flera än håren på mitt huvud äro de som hata mig utan sak; många äro de som vilja förgöra mig, de som äro mina fiender utan skäl; vad jag icke har rövat, det måste jag gälda.
Du, o Gud, känner min dårskap, och mina skulder äro icke förborgade för dig.
Låt icke i mig dem komma på skam, som förbida dig, Herre, HERRE Sebaot; Låt icke i mig dem varda till blygd, som söka dig, du Israels Gud.
Ty för din skull bär jag smälek, för din skull höljer blygsel mitt ansikte;
främmande har jag blivit för mina bröder och en främling för min moders barn.
Ty nitälskan för ditt hus har förtärt mig, och dina smädares smädelser hava fallit över mig.
Jag grät, ja, min själ grät under fasta, men det blev mig till smälek.
Jag klädde mig i sorgdräkt, men jag blev för dem ett ordspråk.
Om mig tassla de, när de sitta i porten; i dryckeslag göra de visor om mig.
Men jag kommer med min bön till dig, HERRE, i behaglig tid, genom din stora nåd, o Gud; svara mig i din frälsande trofasthet.
Rädda mig ur dyn, så att jag icke sjunker ned; låt mig bliva räddad från dem som hata mig och från de djupa vattnen.
Låt icke vattensvallet fördränka mig eller djupet uppsluka mig; och låt ej graven tillsluta sitt gap över mig.
Svara mig, HERRE, ty god är din nåd; vänd dig till mig efter din stora barmhärtighet.
Fördölj icke ditt ansikte för din tjänare, ty jag är i nöd; skynda att svara mig.
Kom till min själ och förlossa henne; befria mig för mina fienders skull.
Du känner min smälek, min skam och blygd; du ser alla mina ovänner.
Smälek har krossat mitt hjärta, så att jag är vanmäktig; jag väntade på medlidande, men där var intet, och på tröstare, men jag fann ingen.
De gåvo mig galla att äta, och ättika att dricka, i min törst.
Må deras bord framför dem bliva till en snara och till ett giller, bäst de gå där säkra;
må deras ögon förmörkas, så att de icke se; gör deras länder vacklande alltid.
Gjut ut över dem din ogunst, och låt din vredes glöd hinna upp dem.
Deras gård blive öde, ingen må finnas, som bor i deras hyddor,
eftersom de förfölja dem som du själv har slagit och orda om huru de plågas, som du har stungit.
Låt dem gå från missgärning till missgärning, och låt dem icke komma till din rättfärdighet.
Må de utplånas ur de levandes bok och icke varda uppskrivna bland de rättfärdiga.
Men mig som är betryckt och plågad, mig skall din frälsning, o Gud, beskydda.
Jag vill lova Guds namn med sång och upphöja honom med tacksägelse.
Det skall behaga HERREN bättre än någon tjur, något offerdjur med horn och klövar.
När de ödmjuka se det, skola de glädja sig; I som söken Gud, edra hjärtan skola leva.
Ty HERREN lyssnar till de fattiga och föraktar icke sina fångna.
Honom love himmelen och jorden, havet och allt vad som rör sig däri.
Ty Gud skall frälsa Sion, han skall bygga upp Juda städer; man skall bo i dem och besitta landet.
Hans tjänares barn skola få det till arvedel, och de som älska hans namn skola bo däri.
För sångmästaren; av David, till åminnelse.
Gud, kom till min räddning; HERRE, skynda till min hjälp.
Må de komma på skam och varda utskämda, som stå efter mitt liv; må de vika tillbaka och blygas, som önska min ofärd.
Må de vända tillbaka i sin skam, som säga: »Rätt så, rätt så!»
Men alla de som söka dig må fröjdas och vara glada i dig; och de som åstunda din frälsning säge alltid: »Lovad vare Gud!»
Jag är betryckt och fattig; Gud, skynda till mig.
Min hjälp och min befriare är du; HERRE, dröj icke.
Till dig, HERRE, tager jag min tillflykt; låt mig aldrig komma på skam.
Rädda mig och befria mig genom din rättfärdighet; böj ditt öra till mig och fräls mig.
Var mig en klippa där jag får bo, och dit jag alltid kan fly, du som beskär mig frälsning.
Ty du är mitt bergfäste och min borg.
Min Gud, befria mig ur den ogudaktiges våld, ur den orättfärdiges och förtryckarens hand.
Ty du är mitt hopp, o Herre, HERRE, du är min förtröstan allt ifrån min ungdom.
Du har varit mitt stöd allt ifrån moderlivet, ja, du har förlöst mig ur min moders liv; dig gäller ständigt mitt lov.
Jag har blivit såsom ett vidunder för många; men du är min starka tillflykt.
Låt min mun vara full av ditt lov, hela dagen av din ära.
Förkasta mig icke i min ålderdoms tid, övergiv mig ej, när min kraft försvinner.
Ty mina fiender säga så om mig, och de som vakta på min själ rådslå så med varandra:
»Gud har övergivit honom; förföljen och gripen honom, ty det finnes ingen som räddar.»
Gud, var icke långt ifrån mig; min Gud, skynda till min hjälp.
Må de komma på skam och förgås, som stå emot min själ; må de höljas med smälek och blygd, som söka min ofärd.
Men jag skall alltid hoppas och än mer föröka allt ditt lov.
Min mun skall förtälja din rättfärdighet, hela dagen din frälsning, ty jag känner intet mått därpå.
Jag skall frambära Herrens, HERRENS väldiga gärningar; jag skall prisa din rättfärdighet, ja, din allenast.
Gud, du har undervisat mig allt ifrån min ungdom; och intill nu förkunnar jag dina under.
Så övergiv mig ej heller, o Gud, i min ålderdom, när jag varder grå, till dess jag får förtälja om din arm för ett annat släkte, om din makt för alla dem som skola komma.
Din rättfärdighet når till himmelen, o Gud.
Du som har gjort så stora ting, o Gud, vem är dig lik?
Du som har låtit oss pröva så mycken nöd och olycka, du skall åter göra oss levande och föra oss upp igen du jordens djup.
Ja, låt mig växa till alltmer; och trösta mig igen.
Så vill ock jag tacka dig med psaltarspel för din trofasthet, min Gud; jag vill lovsjunga dig till harpa, du Israels Helige.
Mina läppar skola jubla, ty jag vill lovsjunga dig; ja, jubla skall min själ, som du har förlossat.
Och min tunga skall hela dagen tala om din rättfärdighet; ty de som sökte min ofärd hava kommit på skam och måst blygas.
Av Salomo.
Gud, giv åt konungen dina rätter och din rättfärdighet åt konungasonen.
Han döme ditt folk med rättfärdighet och dina betryckta med rätt.
Bergen bäre frid åt folket, så ock höjderna, genom rättfärdighet.
Han skaffe rätt åt de betryckta i folket, han frälse de fattiga och krosse förtryckaren.
Dig frukte man, så länge solen varar, och så länge månen skiner, från släkte till släkte.
Han vare lik regnet som faller på ängen, lik en regnskur som vattnar jorden.
I hans dagar blomstre den rättfärdige, och stor frid råde, till dess ingen måne mer finnes.
Må han härska från hav till hav och ifrån floden intill jordens ändar.
För honom buge sig öknens inbyggare, och hans fiender slicke stoftet.
Konungarna från Tarsis och havsländerna hembäre skänker, konungarna av Saba och Seba bäre fram gåvor.
Ja, alla konungar falle ned för honom, alla hedningar tjäne honom.
Ty han skall rädda den fattige som ropar och den betryckte och den som ingen hjälpare har.
Han skall vara mild mot den arme och fattige; de fattigas själar skall han frälsa.
Ifrån förtryck och våld skall han förlossa deras själ, och deras blod skall aktas dyrt i hans ögon.
Må han leva; må man föra till honom guld från Saba.
Ständigt bedje man för honom, alltid välsigne man honom.
Ymnigt växe säden i landet, ända till bergens topp; dess frukt må susa likasom Libanons skog; och folk blomstre upp i städerna såsom örter på marken.
Hans namn förblive evinnerligen; så länge solen skiner, fortplante sig hans namn.
Och i honom välsigne man sig; alla hedningar prise honom säll.
Lovad vare HERREN Gud, Israels Gud, som allena gör under!
Och lovat vare hans härliga namn evinnerligen, och hela jorden vare full av hans ära!
Amen, Amen.
Slut på Davids, Isais sons, böner.
Tredje boken
En psalm av Asaf.
Sannerligen, Gud är god mot Israel, mot dem som hava rena hjärtan.
Men jag hade så när stapplat med mina fötter, mina steg voro nära att slinta;
ty jag upptändes av avund mot de övermodiga, när jag såg att det gick dem väl i deras ogudaktighet.
Ty fria ifrån vedermödor äro de till sin död, och deras hull är frodigt.
De komma icke i olycka såsom andra dödliga och varda icke plågade såsom andra människor.
Därför är högmod deras halsprydnad, våld den klädnad som höljer dem.
Ur fetma skåda deras ögon fram, deras hjärtans inbillningar hava intet mått.
De håna och tala förtryck i sin ondska; med höga åthävor tala de.
Med sin mun stiga de upp i himmelen, och deras tunga far fram på jorden;
därför vänder sig deras folk till dem och super så in vattnet i fulla drag.
Och de säga: »Huru skulle Gud kunna veta det?
Skulle sådan kunskap finnas hos den Högste?»
Ja, så är det med de ogudaktiga; det går dem alltid väl, och de växa i makt.
Sannerligen, förgäves bevarade jag mitt hjärta rent och tvådde mina händer i oskuld;
jag vart dock plågad hela dagen, och var morgon kom tuktan över mig.
Om jag hade sagt: »Så vill jag lära», då hade jag svikit dina barns släkte.
När jag nu tänkte efter för att begripa detta, syntes det mig alltför svårt,
till dess jag trängde in i Guds heliga rådslut och aktade på dess ände.
Sannerligen, på slipprig mark ställer du dem, du störtar dem ned i fördärv.
Huru varda de ej till intet i ett ögonblick!
De förgås och få en ände med förskräckelse.
Såsom det är med en dröm, när man vaknar, o Herre, så aktar du dem för intet, såsom skuggbilder, när du vaknar.
När mitt hjärta förbittrades och jag kände styng i mitt inre,
då var jag oförnuftig och förstod intet; såsom ett oskäligt djur var jag inför dig.
Dock förbliver jag städse hos dig; du håller mig vid min högra hand.
Du skall leda mig efter ditt råd och sedan upptaga mig med ära.
Vem har jag i himmelen utom dig!
Och när jag har dig, då frågar jag efter intet på jorden.
Om än min kropp och min själ försmäkta, så är dock Gud mitt hjärtas klippa och min del evinnerligen.
Ty se, de som hava vikit bort ifrån dig skola förgås; du förgör var och en som trolöst avfaller från dig.
Men jag har min glädje i att hålla mig intill Gud; jag söker min tillflykt hos Herren, HERREN, för att kunna förtälja alla dina gärningar.
En sång av Asaf.
Varför, o Gud, har du så alldeles förkastat oss, varför ryker din vredes eld mot fåren i din hjord?
Tänk på din menighet, som du i fordom tid förvärvade, som du förlossade, till att bliva din arvedels stam; tänk på Sions berg, där du har din boning.
Vänd dina steg till den plats där evig förödelse råder; allt har ju fienden fördärvat i helgedomen.
Dina ovänner hava skränat inne i ditt församlingshus, de hava satt upp sina tecken såsom rätta tecken.
Det var en syn, såsom när man höjer yxor mot en tjock skog.
Och alla dess snidverk hava de nu krossat med yxa och bila.
De hava satt eld på din helgedom och oskärat ända till grunden ditt namns boning.
De hava sagt i sina hjärtan: »Vi vilja alldeles kuva dem.»
Alla Guds församlingshus hava de bränt upp här i landet.
Våra tecken se vi icke; ingen profet finnes mer, och hos oss är ingen som vet för huru länge.
Huru länge, och Gud, skall ovännen få smäda och fienden oavlåtligen få förakta ditt namn?
Varför håller du tillbaka din hand, din högra hand?
Drag den fram ur din barm och förgör dem.
Gud, du är ju min konung av ålder, du är den som skaffar frälsning på jorden.
Det var du som delade havet genom din makt; du krossade drakarnas huvuden mot vattnet.
Det var du som bräckte Leviatans huvuden och gav honom till mat åt öknens skaror.
Det var du som lät källa och bäck bryta fram; du lät ock starka strömmar uttorka.
Din är dagen, din är ock natten, du har berett ljuset och solen.
Det är du som har fastställt alla jordens gränser; sommar och vinter äro skapade av dig.
Så tänk nu på huru fienden smädar HERREN, och huru ett dåraktigt folk föraktar ditt namn.
Lämna ej ut åt vilddjuren din turturduvas själ; förgät icke för alltid dina betrycktas liv.
Tänk på förbundet; ty i landets smygvrår finnes fullt upp av våldsnästen.
Låt icke den förtryckte vika tillbaka med blygd, låt den betryckte och den fattige lova ditt namn.
Stå upp, o Gud; utför din sak.
Betänk huru du varder smädad hela dagen av dåren.
Glöm icke bort dina ovänners rop, dina motståndares larm, som alltjämt höjes.
För sångmästaren; »Fördärva icke»; en psalm, en sång av Asaf.
Vi tacka dig, o Gud, vi tacka dig.
Ditt namn är oss nära; man förtäljer dina under.
»Om jag än bidar min tid, så dömer jag dock rätt.
Om än jorden är i upplösning med alla som bo därpå, så håller dock jag dess pelare stadiga.»
Sela.
Jag säger till de övermodiga: »Varen icke övermodiga», och till de ogudaktiga: »Upphöjen ej hornet.»
Ja, upphöjen icke så högt edert horn, talen ej så hårdnackat vad fräckt är.
Ty icke från öster eller väster, ej heller från bergsöknen kommer hjälpen;
nej, Gud är den som dömer; den ene ödmjukar han, den andre upphöjer han.
Ty en kalk är i HERRENS hand, den skummar av vin och är full av tillblandad dryck, och han skänker i därav; sannerligen, alla ogudaktiga på jorden måste dricka dess drägg i botten.
Men jag skall förkunna det evinnerligen, jag skall lovsjunga Jakobs Gud.
Och de ogudaktigas alla horn skall jag få hugga av; men den rättfärdiges horn skola varda upphöjda.
För sångmästaren, med strängaspel; en psalm, en sång av Asaf.
Gud är känd i Juda, i Israel är hans namn stort;
i Salem vart hans hydda rest och hans boning på Sion.
Där bröt han sönder bågens ljungeldar, sköld och svärd och vad till kriget hör.
Sela.
Full av ljus och härlighet går du fram ifrån segerbytenas berg.
De stormodiga äro avväpnade, de hava slumrat in och sova; alla stridsmännen hava måst låta händerna falla.
För din näpst, du Jakobs Gud, ligga domnade både man och häst.
Du, du är fruktansvärd; vem kan bestå inför dig, när du vredgas?
Från himmelen lät du höra din dom; då förskräcktes jorden och vart stilla,
då när Gud stod upp till dom, till att frälsa alla ödmjuka på jorden.
Sela.
Ty människors vrede varder dig till pris; du har vrede till övers att omgjorda dit med.
Gören löften och infrien dem åt HERREN, eder Gud; alla de som äro omkring honom bäre fram skänker åt den Fruktansvärde.
Ty han stäcker furstarnas övermod; fruktansvärd är han för konungarna på jorden.
För sångmästaren, till Jedutun; av Asaf; en psalm.
Jag vill höja min röst till Gud och ropa; jag vill höja min röst till Gud, för att han må lyssna till mig.
På min nöds dag söker jag Herren; min hand är utsträckt om natten och förtröttas icke; min själ vill icke låta trösta sig.
Jag vill tänka på Gud och klaga; jag vill utgjuta mitt bekymmer, ty min ande försmäktar.
Sela.
Mina ögonlock håller du öppna; jag är full av oro och kan icke tala.
Jag tänker på forntidens dagar, på år som längesedan hava gått.
Jag vill om natten komma ihåg mitt strängaspel; i mitt hjärta vill jag utgjuta mitt bekymmer, och min ande skall eftersinna.
Skall då Herren förkasta evinnerligen och ingen nåd mer bevisa?
Är det då ute med hans godhet för beständigt, har hans ord blivit till intet för alla tider?
Har Gud förgätit att vara nådig eller i vrede tillslutit sin barmhärtighet?
Sela.
Jag svarar: Nej, detta är min plågas tid, den Högstes högra hand är ej såsom förr.
Jag vill prisa HERRENS gärningar, ja, jag vill tänka på dina fordomtima under;
jag vill begrunda alla dina gärningar och eftersinna dina verk.
Gud, i helighet går din väg; vem är en gud så stor som Gud?
Du är Gud, en Gud som gör under; du har uppenbarat din makt bland folken.
Med väldig arm förlossade du ditt folk, Jakobs och Josefs barn.
Sela.
Vattnen sågo dig, och Gud, vattnen sågo dig och våndades, själva djupen darrade.
Molnen göto ut strömmar av vatten, skyarna läto höra sin röst, och dina pilar foro omkring.
Ditt dunder ljöd i stormvirveln, ljungeldar lyste upp jordens krets, jorden darrade och bävade.
Genom havet gick din väg, din stig genom stora vatten, och dina fotspår fann man icke.
Så förde du ditt folk såsom en hjord genom Moses och Arons hand.
En sång av Asaf.
Lyssna, mitt folk, till min undervisning; böjen edra öron till min muns ord.
Jag vill öppna min mun till lärorikt tal, uppenbara förborgade ting ifrån fordom.
Vad vi hava hört och känna, och vad våra fäder hava förtäljt för oss,
det vilja vi icke dölja för deras barn; för ett kommande släkte vilja vi förtälja HERRENS lov och hans makt och de under han har gjort.
Ty han upprättade ett vittnesbörd i Jakob och stiftade en lag i Israel; han påbjöd den för våra fäder, och de skulle kungöra den för sina barn.
Så skulle det bliva kunnigt för ett kommande släkte, för barn som en gång skulle födas, och dessa skulle stå upp och förtälja det för sina barn.
Då skulle de sätta sitt hopp till Gud och icke förgäta Guds verk, utan taga hans bud i akt.
Och de skulle icke bliva, såsom deras fäder, ett gensträvigt och upproriskt släkte, ett släkte som icke höll sitt hjärta ståndaktigt, och vars ande icke var trofast mot Gud.
Efraims barn, välbeväpnade bågskyttar, vände om på stridens dag.
De höllo icke Guds förbund, och efter hans lag ville de ej vandra.
De glömde hans gärningar och de under han hade låtit dem se.
Ja, inför deras fäder hade han gjort under, i Egyptens land, på Soans mark.
Han klöv havet och lät dem gå därigenom och lät vattnet stå såsom en hög.
Han ledde dem om dagen med molnskyn, och hela natten med eldens sken.
Han klöv sönder klippor i öknen och gav dem rikligen att dricka, såsom ur väldiga hav.
Rinnande bäckar lät han framgå ur klippan och vatten flyta ned såsom strömmar.
Likväl syndade de allt framgent mot honom och voro gensträviga mot den Högste, i öknen.
De frestade Gud i sina hjärtan, i det de begärde mat för sin lystnad.
Och de talade mot Gud, de sade: »Kan väl Gud duka ett bord i öknen?
Se, visst slog han klippan, så att vatten flödade och bäckar strömmade fram, men kan han ock giva bröd eller skaffa kött åt sitt folk?»
Så förgrymmades då HERREN, när han hörde det; och eld upptändes i Jakob, jag, vrede kom över Israel,
eftersom de icke trodde på Gud och ej förtröstade på hans frälsning.
Och han gav befallning åt skyarna i höjden och öppnade himmelens dörrar;
han lät manna regna över dem till föda, och korn från himmelen gav han dem.
Änglabröd fingo människor äta; han sände dem mat till fyllest.
Han lät östanvinden fara ut på himmelen, och genom sin makt förde han sunnanvinden fram.
Och han lät kött regna över dem såsom stoft, bevingade fåglar såsom havets sand;
han lät det falla ned i sitt läger, runt omkring sin boning.
Då åto de och blevo övermätta; han lät dem få vad de hade lystnad efter.
Men ännu hade de icke stillat sin lystnad, ännu var maten i deras mun,
då kom Guds vrede över dem; han sände död bland deras ypperste och slog ned Israels unga män.
Likväl syndade de alltjämt och trodde icke på hans under.
Då lät han deras dagar försvinna i förgängelse och deras år i plötslig undergång.
När han dräpte folket, frågade de efter honom och vände om och sökte Gud.
De tänkte då på att Gud var deras klippa, och att Gud den Högste var deras förlossare;
och de talade inställsamt för honom med sin mun och skrymtade för honom med sin tunga.
Men deras hjärtan höllo sig icke ståndaktigt vid honom, och de voro icke trogna i hans förbund.
Dock, han är barmhärtig, han förlåter missgärning, och han vill icke fördärva.
Därför avvände han ofta sin vrede och lät ej hela sin förtörnelse bryta fram.
Ty han tänkte därpå att de voro kött, en vind som far bort och icke kommer åter.
Huru ofta voro de ej gensträviga mot honom i öknen och bedrövade honom i ödemarken!
Ja, de frestade Gud allt framgent och förtörnade Israels Helige.
De betänkte icke vad hans hand hade uträttat på den tid då han förlossade dem från ovännen,
då han gjorde sina tecken i Egypten och sina under på Soans mark.
Där förvandlade han deras strömmar till blod, så att de ej kunde dricka ur sina rinnande vatten;
han sände bland dem flugsvärmar, som åto dem, och paddor, som voro dem till fördärv.
Han gav deras gröda åt gräsmaskar och deras arbetes frukt åt gräshoppor;
han slog deras vinträd med hagel och deras fikonträd med hagelstenar;
han gav deras husdjur till pris åt hagel och deras boskap åt ljungeldar.
Han sände över dem sin vredes glöd, förgrymmelse och ogunst och nöd, en skara av olycksänglar.
Han gav fritt lopp åt sin vrede; han skonade icke deras själ från döden, utan gav deras liv till pris åt pesten.
Och han slog allt förstfött i Egypten, kraftens förstling i Hams hyddor.
Och han lät sitt folk bryta upp såsom en fårhjord och förde dem såsom en boskapshjord genom öknen.
Han ledde dem säkert, så att de icke behövde frukta; men deras fiender övertäcktes av havet.
Och han lät dem komma till sitt heliga land, till det berg som hans högra hand hade förvärvat.
Han förjagade hedningarna för dem och gav dem deras land till arvslott och lät Israels stammar bo i deras hyddor.
Men i sin gensträvighet frestade de Gud den Högste och höllo icke hans vittnesbörd;
de veko trolöst tillbaka, de såsom deras fäder, de vände om, lika en båge som sviker.
De förtörnade honom med sina offerhöjder och retade honom genom sina beläten.
Gud förnam det och vart förgrymmad och förkastade Israel med harm.
Och han försköt sin boning i Silo, det tält han hade slagit upp bland människorna;
han gav sin makt i fångenskap och sin ära i fiendehand.
Ja, han gav sitt folk till pris åt svärdet, och på sin arvedel förgrymmades han.
Deras unga män förtärdes av eld, och deras jungfrur blevo utan brudsång.
Deras präster föllo för svärd, och inga änkor kunde hålla klagogråt.
Då vaknade Herren såsom ur en sömn, han reste sig, lik en hjälte som hade legat dövad av vin.
Och han slog sina ovänner tillbaka, evig smälek lät han komma över dem.
Han förkastade ock Josefs hydda och utvalde icke Efraims stam.
Men han utvalde Juda stam, Sions berg, som han älskade.
Och han byggde sin helgedom hög såsom himmelen, fast såsom jorden, som han har grundat för evigt.
Och han utvalde sin tjänare David och tog honom ifrån fårhjordens fållor.
Ja, ifrån fåren hämtade han honom och satte honom till en herde för Jakob, sitt folk, och för Israel, sin arvedel.
Och han var deras herde med redligt hjärta och ledde dem med förståndig hand.
En psalm av Asaf.
Gud, hedningarna hava fallit in i din arvedel, de hava orenat ditt heliga tempel, de hava gjort Jerusalem till en stenhop.
De hava givit dina tjänares kroppar till mat åt himmelens fåglar, dina frommas kött åt markens djur.
De hava utgjutit deras blod såsom vatten, runt omkring Jerusalem, och ingen fanns, som begrov dem.
Vi hava blivit till smälek för våra grannar, till spott och hån för dem som bo omkring oss.
Huru länge, o HERRE, skall du så oavlåtligen vredgas, huru länge skall din nitälskan brinna såsom eld?
Utgjut din förtörnelse över hedningarna, som ej känna dig, och över de riken som icke åkalla ditt namn.
Ty de hava uppätit Jakob, och hans boning hava de förött.
Tänk ej, oss till men, på förfädernas missgärningar, låt din barmhärtighet snarligen komma oss till mötes, ty vi äro i stort elände.
Hjälp oss, du vår frälsnings Gud, för ditt namns äras skull; rädda oss och förlåt oss våra synder för ditt namns skull.
Varför skulle hedningarna få säga: »Var är nu deras Gud?»
Låt det inför våra ögon bliva kunnigt på hedningarna huru du hämnas dina tjänares utgjutna blod.
Låt de fångnas klagan komma inför ditt ansikte, låt efter din arms väldighet dödens barn bliva vid liv.
Och giv våra grannar sjufalt tillbaka i deras sköte den smädelse varmed de hava smädat dig, Herre.
Men vi som äro ditt folk och får i din hjord, vi vilja tacka dig evinnerligen, vi vilja förtälja ditt lov från släkte till släkte.
För sångmästaren, efter »Liljor»; ett vittnesbörd; av Asaf; en psalm.
Lyssna, du Israels herde, du som leder Josef såsom din hjord; du som tronar på keruberna, träd fram i glans.
Låt din makt vakna upp till att gå framför Efraim och Benjamin och Manasse, och kom till vår frälsning.
Gud, upprätta oss, och låt ditt ansikte lysa, så att vi varda frälsta.
HERRE Gud Sebaot, huru länge skall du vredgas vid ditt folks bön?
Du har låtit dem äta tårebröd och givit dem tårar att dricka i fullt mått.
Du gör oss till ett trätoämne för våra grannar, och våra fiender bespotta oss.
Gud Sebaot, upprätta oss, och låt ditt ansikte lysa, så att vi varda frälsta.
Ett vinträd flyttade du från Egypten, du förjagade hedningarna och planterade det.
Du röjde rum för det, och det slog rötter och uppfyllde landet.
Bergen blevo betäckta av dess skugga och Guds cedrar av dess rankor;
det utbredde sina revor ända till havet och sina telningar intill floden.
Varför har du då brutit ned dess hägnad, så att alla vägfarande riva till sig därav?
Vildsvinet från skogen frossar därpå, och djuren på marken äta därav.
Gud Sebaot, vänd åter, skåda ned från himmelen och se härtill, och låt dig vårda om detta vinträd.
Skydda trädet som din högra hand har planterat, och den son som du har fostrat åt dig.
Det är förbränt av eld och kringhugget; för ditt ansiktes näpst förgås de.
Håll din hand över din högra hands man, över den människoson som du har fostrat åt dig.
Då skola vi icke vika ifrån dig; behåll oss vid liv, så skola vi åkalla ditt namn.
HERRE Gud Sebaot, upprätta oss; låt ditt ansikte lysa, så att vi varda frälsta.
För sångmästaren, till Gittít; av Asaf.
Höjen glädjerop till Gud, vår starkhet, höjen jubel till Jakobs Gud.
Stämmen upp lovsång och låten pukor ljuda, ljuvliga harpor tillsammans med psaltare.
Stöten i basun vid nymånaden, vid fullmånen, på vår högtidsdag.
Ty detta är en stadga för Israel, en Jakobs Guds rätt.
Det bestämde han till ett vittnesbörd i Josef, när han drog ut mot Egyptens land.
Jag hör ett tal som är mig nytt:
»Jag lyfte bördan från hans skuldra, hans händer blevo fria ifrån lastkorgen.
I nöden ropade du, och jag räddade dig; jag svarade dig, höljd i tordön, jag prövade dig vid Meribas vatten.
Sela.
Hör, mitt folk, och låt mig varna dig; Israel, o att du ville höra mig!
Hos dig skall icke finnas någon annan gud, och du skall ej tillbedja någon främmande gud.
Jag är HERREN, din Gud, som har fört dig upp ur Egyptens land; låt din mun vitt upp, så att jag får uppfylla den.
Men mitt folk ville ej höra min röst, och Israel var mig icke till viljes.
Då lät jag dem gå i deras hjärtans hårdhet, det fingo vandra efter sina egna rådslag.
O att mitt folk ville höra mig, och att Israel ville vandra på mina vägar!
Då skulle jag snart kuva deras fiender och vända min hand mot deras ovänner.
De som hata HERREN skulle då visa honom underdånighet, och hans folks tid skulle vara evinnerligen.
Och han skulle bespisa det med bästa vete; ja, med honung ur klippan skulle jag mätta dig.»
En psalm av Asaf.
Gud står i gudaförsamlingen, mitt ibland gudarna håller han dom:
»Huru länge skolen I döma orätt och vara partiska för de ogudaktiga?
Sela.
Skaffen den arme och faderlöse rätt, given den betryckte och torftige rättvisa.
Befrien den arme och fattige, rädden honom från de ogudaktigas hand.
Men de veta intet och hava intet förstånd, de vandra i mörker; jordens alla grundvalar vackla.
Jag har väl sagt att I ären gudar och allasammans den Högstes söner;
men I måsten dock dö, såsom människor dö, och falla, likaväl som var furste faller.»
Ja, stå upp, o Gud; håll dom över jorden, ty med arvsrätt råder du över alla folk.
En sång, en psalm av Asaf.
Gud, var icke så tyst, tig icke och var icke så stilla, o Gud.
Ty se, dina fiender larma, och de som hata dig resa upp huvudet.
Mot ditt folk förehava de listiga anslag och rådslå mot dem som du beskyddar.
De säga: »Kom, låt oss utrota dem, så att de ej mer äro ett folk, och så att ingen mer tänker på Israels namn.»
Ty endräktigt rådslå dem med varandra, de sluta mot dig ett förbund:
Edoms tält och ismaeliterna, Moab och hagariterna,
Gebal och Ammon och Amalek, filistéerna tillika med dem som bo i Tyrus;
Assur har ock slutit sig till dem, han har lånat sin arm åt Lots barn.
Sela.
Gör med dem såsom du gjorde med Midjan, såsom med Sisera och Jabin vid Kisons bäck,
dem som förgjordes vid En-Dor och blevo till gödning åt marken.
Låt det gå deras ädlingar såsom det gick Oreb och Seeb, och alla deras furstar såsom det gick Seba och Salmunna,
eftersom de säga: »Guds ängder vilja vi intaga åt oss.»
Min Gud, låt dem bliva såsom virvlande löv, såsom strå för vinden.
Lik en eld som förbränner skog och lik en låga som avsvedjar berg
förfölje du dem med ditt oväder, och förskräcke du dem med din storm.
Gör deras ansikten fulla med skam, så att de söka ditt namn, o HERRE.
Ja, må de komma på skam och förskräckas till evig tid, må de få blygas och förgås.
Och må de förnimma att du allena bär namnet »HERREN», den Högste över hela jorden.
För sångmästaren, till Gittít; av Koras söner; en psalm.
Huru ljuvliga äro icke dina boningar, HERRE Sebaot!
Min själ längtar och trängtar efter HERRENS gårdar, min själ och min kropp jubla mot levande Gud.
Ty sparven har funnit ett hus och svalan ett bo åt sig, där hon kan lägga sina ungar: dina altaren, HERRE Sebaot, min konung och min Gud.
Saliga äro de som bo i ditt hus; de lova dig beständigt.
Sela.
Saliga äro de människor som i dig hava sin starkhet, de vilkas håg står till dina vägar.
När de vandra genom Tåredalen, göra de den rik på källor, och höstregnet höljer den med välsignelser.
De gå från kraft till kraft; så träda de fram inför Gud på Sion.
HERRE Gud Sebaot, hör min bön, lyssna, du Jakobs Gud.
Sela.
Gud, vår sköld, ser härtill, och akta på din smordes ansikte.
Ty en dag i dina gårdar är bättre än eljest tusen.
Jag vill hellre vakta dörren i min Guds hus än dväljas i de ogudaktigas hyddor.
Ty HERREN Gud är sol och sköld; HERREN giver nåd och ära; han vägrar icke dem något gott, som vandra i ostrafflighet.
HERRE Sebaot, salig är den människa som förtröstar på dig.
För sångmästaren; av Koras söner; en psalm.
HERRE, du var förr ditt land nådig, du upprättade åter Jakobs hus.
Du förlät ditt folks missgärning, du överskylde all dess synd.
Sela.
Du lät all din förgrymmelse fara och vände dig ifrån din vredes glöd.
Så vänd dig nu åter till oss, du vår frälsnings Gud, och upphör med din förtörnelse mot oss.
Vill du då vredgas på oss evinnerligen och låta din vrede vara från släkte till släkte?
Vill du icke åter giva oss liv, så att ditt folk får glädjas i dig?
HERRE, låt oss se din nåd, och giv oss din frälsning.
Jag vill höra vad Gud, HERREN, talar: se, han talar frid till sitt folk och till sina fromma; må de blott icke vända åter till dårskap.
Ja, hans frälsning är nära dem som frukta honom, och så skall ära bo i vårt land.
Godhet och trofasthet skola där mötas, rättfärdighet och frid kyssas;
trofasthet skall växa upp ur jorden och rättfärdighet blicka ned från himmelen.
HERREN skall giva oss vad gott är, och vårt land skall giva sin gröda.
Rättfärdighet skall gå framför honom, den skall ock stadigt följa i hans spår.
En bön av David.
HERRE, böj till mig ditt öra och svara mig, ty jag är betryckt och fattig.
Bevara min själ, ty jag är from; du min Gud, fräls din tjänare, som förtröstar på dig.
Var mig nådig, o Herre, ty hela dagen ropar jag till dig.
Gläd din tjänares själ, ty till dig, Herre, upplyfter jag min själ.
Ty du, o Herre, är god och förlåtande och stor i nåd mot alla som åkalla dig.
Lyssna, HERRE, till mitt bedjande, och akta på mina böners ljud.
På min nöds dag åkallar jag dig, ty du skall svara mig.
Ingen är dig lik bland gudarna, Herre, och intet är såsom dina verk.
Hedningarna, som du har gjort, skola alla komma och tillbedja inför dig, Herre, och skola ära ditt namn.
Ty du är stor, och du gör stora under; du allena är Gud.
Visa mig, HERRE, din väg; jag vill vandra i din sanning.
Behåll mitt hjärta vid det ena att jag fruktar ditt namn.
Då vill jag tacka dig, Herre, min Gud, av allt mitt hjärta och ära ditt namn evinnerligen;
ty din nåd är stor över mig, och du räddar min själ ur dödsrikets djup.
Gud, fräcka människor hava rest sig upp mot mig, och våldsverkarnas hop står efter mitt liv; de hava icke dig för ögonen.
Men du, Herre, är en barmhärtig och nådig Gud, långmodig och stor i mildhet och trofasthet.
Vänd dig till mig och var mig nådig, giv åt din tjänare din makt, och fräls din tjänarinnas son.
Gör ett tecken med mig, så att det går mig väl; och må de som hata mig se med blygd att du, o HERRE, hjälper mig och tröstar mig.
Av Koras söner; en psalm, en sång.
Den stad han har grundat står på de heliga bergen;
HERREN älskar Sions portar mest bland alla Jakobs boningar.
Härliga ting äro talade om dig, du Guds stad.
Sela.
»Rahab och Babel skall jag nämna bland mina bekännare; så ock Filisteen och Tyrus och Kus, dessa äro födda där.»
Ja, om Sion skall det sägas: »Den ene som den andre är född därinne.»
Och han, den Högste, skall hålla det vid makt.
Ja, när HERREN tecknar upp folken, då skall han räkna så: »Dessa äro födda där.»
Sela.
Och under sång och dans skall man säga: »Alla mina källor äro i dig.»
En sång, en psalm av Koras söner; för sångmästaren, till Mahalat-leannót; en sång av esraiten Heman.
HERRE, min frälsnings Gud, dag och natt ropar jag inför dig.
Låt min bön komma inför ditt ansikte, böj ditt öra till mitt rop.
Ty min själ är mättad med lidanden, och mitt liv har kommit nära dödsriket.
Jag är aktad lik dem som hava farit ned i graven, jag är såsom en man utan livskraft.
Jag är övergiven bland de döda, lik de slagna som ligga i graven, dem på vilka du icke mer tänker, och som äro avskilda från din hand.
Ja, du har sänkt mig ned underst i graven, ned i mörkret, ned i djupet.
Den vrede vilar tung på mig, och alla dina böljors svall låter du gå över mig.
Sela.
Du har drivit mina förtrogna långt bort ifrån mig; du har gjort mig till en styggelse för dem; jag ligger fången och kan icke komma ut.
Mitt öga förtvinar av lidande; HERRE, jag åkallar dig dagligen, jag uträcker mina händer till dig.
Gör du väl under för de döda, eller kunna skuggorna stå upp och tacka dig?
Sela.
Förtäljer man i graven om din nåd, i avgrunden om din trofasthet?
Känner man i mörkret dina under, och din rättfärdighet i glömskans land?
Men jag ropar till dig, HERRE, och bittida kommer min bön dig till mötes.
Varför förkastar du, HERRE, min själ, varför döljer du ditt ansikte för mig?
Betryckt är jag och döende allt ifrån min ungdom; jag måste bära dina förskräckelser, så att jag är nära att förtvivla.
Din vredes lågor gå över mig, dina fasor förgöra mig.
De omgiva mig beständigt såsom vatten, de kringränna mig allasammans.
Du har drivit vän och frände långt bort ifrån mig; i mina förtrognas ställe har jag nu mörkret.
En sång av esraiten Etan.
Jag vill sjunga om HERRENS nådegärningar evinnerligen; jag vill låta min mun förkunna din trofasthet, från släkte till släkte.
Ja, jag säger: För evig tid skall nåd byggas upp; i himmelen, där befäster du din trofasthet.
»Jag har slutit ett förbund med min utvalde, med ed har jag lovat min tjänare David:
'Jag skall befästa din säd för evig tid och bygga din tron från släkte till släkte.'»
Sela.
Av himlarna prisas dina under, o HERRE, och i de heligas församling din trofasthet.
Ty vilken i skyn kan liknas vid HERREN, vilken bland Guds söner kan aktas lik HERREN?
Ja, Gud är mycket förskräcklig i de heligas råd och fruktansvärd utöver alla som äro omkring honom.
HERRE, härskarornas Gud, vem är dig lik?
Stark är HERREN; och din trofasthet är runt omkring dig.
Du är den som råder över havets uppror; när dess böljor resa sig, stillar du dem.
Du krossade Rahab, så att han låg lik en slagen; med din mäktiga arm förströdde du dina fiender.
Din är himmelen, din är ock jorden; du har grundat jordens krets med allt vad därpå är.
Norr och söder, dem har du skapat; Tabor och Hermon jubla i ditt namn.
Du har en arm med hjältekraft, mäktig är din hand, hög är din högra hand.
Rättfärdighet och rätt äro din trons fäste, nåd och sanning stå inför ditt ansikte.
Saligt är det folk som vet vad jubel är, de som vandra, o HERRE, i ditt ansiktes ljus.
I ditt namn fröjda de sig alltid, och genom din rättfärdighet upphöjas de.
Ty du är deras starkhet och prydnad, och genom din nåd upphöjer du vårt horn.
Ty han som är vår sköld tillhör HERREN, vår konung tillhör Israels Helige.
På den tiden talade du i en syn till dina fromma och sade: »Jag har lagt hjälp i en hjältes hans, jag har upphöjt en yngling ur folket.
Jag har funnit min tjänare David och smort honom med min helig olja.
Min hand skall stadigt vara med honom, och min arm skall styrka honom.
Ingen fiende skall oförtänkt komma över honom, och ingen orättfärdig skall förtrycka honom;
nej, jag skall krossa hans ovänner framför honom, och jag skall hemsöka dem som hata honom.
Min trofasthet och min nåd skola vara med honom, och i mitt namn skall hans horn varda upphöjt.
Jag skall lägga havet under hans hand och strömmarna under hans högra hand.
Han skall kalla mig så: 'Du min fader, min Gud och min frälsnings klippa.'
Ja, jag skall göra honom till den förstfödde, till den högste bland konungarna på jorden.
Jag skall bevara min nåd åt honom evinnerligen, och mitt förbund med honom skall förbliva fast.
Jag skall låta hans säd bestå till evig tid, och hans tron, så länge himmelen varar.
Om hans barn övergiva min lag och icke vandra efter mina rätter,
om de bryta mot mina stadgar och icke hålla mina bud,
då skall jag väl hemsöka deras överträdelse med ris och deras missgärning med plågor,
men min nåd skall jag ej taga ifrån honom, och jag skall icke svika i trofasthet.
Jag skall icke bryta mitt förbund, och vad mina läppar hava talat skall jag ej förändra.
En gång har jag svurit det vid min helighet, och mitt löfte till David skall jag icke bryta.
Hans säd skall förbliva evinnerligen och hans tron inför mig så länge som solen;
såsom månen skall den bestå evinnerligen.
Och trofast är vittnet i skyn.»
Sela.
Men nu har du förkastat och förskjutit din smorde och handlat i vrede mot honom.
Du har upplöst förbundet med din tjänare, du har oskärat hans krona och kastat den ned till jorden.
Du har brutit ned alla hans murar, du har gjort hans fästen till spillror.
Alla som gå vägen fram plundra honom, han har blivit till smälek för sina grannar.
Du har upphöjt hans ovänners högra hand och berett alla hans fiender glädje.
Ja, du har låtit hans svärdsegg vika tillbaka och icke hållit honom uppe i striden.
Du har gjort slut på hans glans och slagit hans tron till jorden.
Du har förkortat hans ungdoms dagar, du har höljt honom med skam.
Sela.
Huru länge, o HERRE, skall du så alldeles fördölja dig?
Huru länge skall din vrede brinna såsom eld?
Tänk på huru kort mitt liv varar, och huru förgängliga du har skapat alla människors barn.
Ty vilken är den man som får leva och undgår att se döden?
Vem räddar din själ från dödsrikets våld?
Sela.
Herre, var äro din forna nådegärningar, vad du lovade David med ed i din trofasthet.
Tänk, Herre, på dina tjänares smälek, på vad jag måste fördraga av alla de många folken;
tänk på huru dina fiender smäda, o HERRE, huru de smäda din smordes fotspår. ----
Lovad vare HERREN evinnerligen!
Amen, Amen.
Fjärde boken
En bön av gudsmannen Mose.
Herre, du har varit vår tillflykt från släkte till släkte.
Förrän bergen blevo till och du frambragte jorden och världen, ja, från evighet till evighet är du, o Gud.
Du låter människorna vända åter till stoft, du säger: »Vänden åter, I människors barn.»
Ty tusen år äro i dina ögon såsom den dag som förgick i går; ja, de äro såsom en nattväkt.
Du sköljer dem bort; de äro såsom en sömn.
Om morgonen likna de gräset som frodas;
det blomstrar upp och frodas om morgonen, men om aftonen torkar det bort och förvissnar.
Ty vi förgås genom din vrede, och genom din förtörnelse ryckas vi plötsligt bort.
Du ställer våra missgärningar inför dig, våra förborgade synder i ditt ansiktes ljus.
Ja, alla våra dagar försvinna genom din förgrymmelse, vi lykta våra år såsom en suck.
Vårt liv varar sjuttio år eller åttio år, om det bliver långt; och när det är som bäst, är det möda och fåfänglighet, ty det går snart förbi, likasom flöge vi bort.
Vem besinnar din vredes makt och din förgrymmelse, så att han fruktar dig?
Lär oss betänka huru få våra dagar äro, för att vi må undfå visa hjärtan.
HERRE, vänd åter.
Huru länge dröjer du?
Förbarma dig över dina tjänare.
Mätta oss med din nåd, när morgonen gryr, så att vi få jubla och vara glada i alla våra livsdagar.
Giv oss glädje så många dagar som du har plågat oss, så många år som vi hava lidit olycka.
Låt dina gärningar uppenbaras för dina tjänare och din härlighet över deras barn.
Och HERRENS, vår Guds, ljuvlighet komme över oss.
Må du främja för oss våra händers verk; ja, våra händers verk främje du.
Den som sitter under den Högstes beskärm och vilar under den Allsmäktiges skugga,
han säger: »I HERREN har jag min tillflykt och min borg, min Gud, på vilken jag förtröstar.»
Ja, han skall rädda dig ifrån fågelfängarens snara och ifrån pesten, som fördärvar.
Med sina fjädrar skall han betäcka dig, och under hans vingar skall du finna tillflykt; hans trofasthet är sköld och skärm.
Du skall icke behöva frukta nattens fasor, icke pilen, som flyger om dagen,
icke pesten, som går fram i mörkret, eller farsoten, som ödelägger vid middagens ljus.
Om ock tusen falla vid din sida, ja, tio tusen vid din högra sida, så skall det dock icke drabba dig.
Dina ögon skola blott skåda därpå med lust, och du skall se de ogudaktigas lön.
Ty du har sagt: »Du, HERRE, är mitt skygd», och du har gjort den Högste till din tillflykt.
Ingen olycka skall vederfaras dig, och ingen plåga skall nalkas din hydda.
Ty han skall giva sina änglar befallning om dig, att de skola bevara dig på alla dina vägar.
De skola bära dig på händerna, så att du icke stöter din fot mot någon sten.
Över lejon och huggormar skall du gå fram, du skall trampa ned unga lejon och drakar.
»Han håller sig intill mig, därför skall jag befria honom; jag skall beskydda honom, därför att han känner mitt namn.
Han åkallar mig, och jag skall svara honom; jag är med honom i nöden, jag skall rädda honom och låta honom komma till ära.
Jag skall mätta honom med långt liv och låta honom se min frälsning.»
En psalm, en sång för sabbatsdagen.
Det är gott att tacka HERREN och att lovsjunga ditt namn, du den Högste,
att om morgonen förkunna din nåd, och när natten har kommit din trofasthet,
med tiosträngat instrument och psaltare, med spel på harpa.
Ty du gläder mig, HERRE, med dina gärningar; jag vill jubla över dina händers verk.
Huru stora äro icke dina verk, o HERRE!
Ja, övermåttan djupa äro dina tankar.
En oförnuftig man besinnar det ej, och en dåre förstår icke sådant.
Om ock de ogudaktiga grönska såsom gräs och ogärningsmännen blomstra allasammans, så sker det till fördärv för evig tid.
Men du, HERRE, är hög evinnerligen.
Ty se, dina fiender, HERRE, se, dina fiender förgås, alla ogärningsmännen bliva förströdda.
Men mitt horn gör du högt såsom vildoxens; jag varder övergjuten med frisk olja.
Och med lust får mitt öga skåda på mina förföljare och mina öron höra om de onda som resa sig upp mot mig.
Den rättfärdige grönskar såsom ett palmträd, såsom en ceder på Libanon växer han till.
Ja, sådana äro planterade i HERRENS hus; de grönska i vår Guds gårdar.
Ännu när de bliva gamla, skjuta de skott, de frodas och grönska;
så för att de skola förkunna att HERREN är rättfärdig, min klippa, han i vilken orätt icke finnes.
HERREN är min konung!
Han har klätt sig i härlighet.
HERREN har klätt sig, omgjordat sig med makt; därför står jordkretsen fast och vacklar icke.
Din tron står fast ifrån fordom tid, du är från evighet.
HERRE, strömmarna hava upphävt, strömmarna hava upphävt sin röst, ja, strömmarna upphäva sitt dån.
Men väldig är HERREN i höjden, mer än bruset av stora vatten, väldiga vatten, havets bränningar.
Dina vittnesbörd äro fasta alltigenom; helighet höves ditt hus, HERRE, evinnerligen.
Du hämndens Gud, o HERRE, du hämndens Gud, träd fram i glans.
Res dig, du jordens domare, vedergäll de högmodiga vad de hava gjort.
Huru länge skola de ogudaktiga, o HERRE, huru länge skola de ogudaktiga triumfera?
Deras mun flödar över av fräckt tal; de förhäva sig, alla ogärningsmännen.
Ditt folk, o HERRE, krossa de, och din arvedel förtrycka de.
Änkor och främlingar dräpa de, och faderlösa mörda de.
Och de säga: »HERREN ser det icke, Jakobs Gud märker det icke.»
Märken själva, I oförnuftiga bland folket; I dårar, när kommen I till förstånd?
Den som har planterat örat, skulle han icke höra?
Den som har danat ögat, skulle han icke se?
Den som håller hedningarna i tukt, skulle han icke straffa, han som lär människorna förstånd?
HERREN känner människornas tankar, han vet att de själva äro fåfänglighet.
Säll är den man som du, HERRE, undervisar, och som du lär genom din lag,
för att skaffa honom ro för olyckans dagar, till dess de ogudaktigas grav varder grävd.
Ty HERREN förskjuter icke sitt folk, och sin arvedel övergiver han icke.
Nej, rättfärdighet skall åter gälla i rätten, och alla rättsinniga skola hålla sig därtill.
Vem står upp till att försvara mig mot de onda, vem bistår mig mot ogärningsmännen?
Om HERREN icke vore min hjälp, så bodde min själ snart i det tysta.
När jag tänkte: »Min fot vacklar», då stödde mig din når, o HERRE:
När jag hade mycket bekymmer i mitt hjärta, då gladde din tröst min själ.
Kan fördärvets domarsäte hava gemenskap med dig, det säte där man över våld i lagens namn,
där de tränga den rättfärdiges själ och fördöma oskyldigt blod?
Men HERREN bliver för mig en borg, min Gud bliver min tillflykts klippa.
Och han låter deras fördärv vända tillbaka över dem och förgör dem för deras ondskas skull.
Ja, HERREN, vår Gud, förgör dem.
Kommen, låtom oss höja glädjerop till HERREN, jubel till vår frälsnings klippa.
Låtom oss träda fram för hans ansikte med tacksägelse och höja jubel till honom med lovsånger.
Ty HERREN är en stor Gud, en stor konung över alla gudar.
Han har jordens djup i sin hand, och bergens höjder äro hans;
hans är havet, ty han har gjort det, och hans händer hava danat det torra.
Kommen, låtom oss tillbedja och nedfalla, låtom oss knäböja för HERREN, vår skapare.
Ty han är vår Gud, och vi äro det folk som han har till sin hjord, vi äro får som stå under hans vård.
O att I villen i dag höra hans röst!
Förhärden icke edra hjärtan såsom i Meriba, såsom på Massas dag i öknen,
där edra fäder frestade mig, där de prövade mig, fastän de hade sett mina verk.
I fyrtio år var det släktet mig till leda, och jag sade: »De äro ett folk som far vilse med sitt hjärta, och de vilja icke veta av mina vägar.»
Så svor jag då i min vrede: »De skola icke komma in i min vila.»
Sjungen till HERRENS ära en ny sång, sjungen till HERRENS ära, alla länder.
Sjungen till HERRENS ära, loven hans namn.
Båden glädje var dag, förkunnen hans frälsning.
Förtäljen bland hedningarna hans ära, bland alla folk hans under.
Ty stor är HERREN och högt lovad, fruktansvärd är han mer än alla gudar.
Ty folkens alla gudar äro avgudar, men HERREN är den som har gjort himmelen.
Majestät och härlighet äro inför hans ansikte, makt och glans i hans helgedom.
Given åt HERREN, I folkens släkter, given åt HERREN ära och makt;
given åt HERREN hans namns ära, bären fram skänker, och kommen i hans gårdar.
Tillbedjen HERREN i helig skrud, bäven för hans ansikte, alla länder.
Sägen bland hedningarna: »HERREN är nu konung!
Därför står jordkretsen fast och vacklar icke; han dömer folken med rättvisa.»
Himmelen vare glad, och jorden fröjde sig; havet bruse och allt vad däri är.
Marken glädje sig och allt som är därpå, ja, då juble alla skogens träd.
inför HERREN, ty han kommer, ty han kommer för att döma jorden.
Han skall döma jordens krets med rättfärdighet och folken med sin trofasthet.
HERREN är nu konung!
Därför fröjde sig jorden; havsländerna glädje sig, så många som de äro.
Moln och töcken omgiva honom, rättfärdighet och rätt äro hans trons fäste.
Eld går framför honom och förbränner hans ovänner runt omkring.
Hans ljungeldar lysa upp jordens krets; jorden ser det och bävar.
Bergen smälta såsom vax för HERREN, för hela jordens Herre.
Himlarna förkunna hans rättfärdighet, och alla folk se hans ära.
Alla de skola komma på skam, som dyrka beläten, de som berömma sig av avgudar.
Alla gudar skola tillbedja honom.
Sion hör det och gläder sig, och Juda döttrar fröjda sig för dina domars skull, HERRE.
Ty du, HERRE, är den Högste över hela jorden; du är högt upphöjd över alla gudar.
I som älsken HERREN, haten det onda.
Han bevarar sina frommas själar, ur de ogudaktigas hand räddar han dem.
Ljus är utsått för den rättfärdige och glädje för de rättsinniga.
Glädjens, I rättfärdige, i HERREN, och prisen hans heliga namn.
En psalm.
Sjungen till HERREN ära en ny sång, ty han har gjort under.
Han har vunnit seger med sin högra hand och med sin väldiga arm.
HERREN har låtit sin frälsning bliva kunnig, han har uppenbarat sin rättfärdighet för hedningarnas ögon.
Han har tänkt på sin nåd och trofasthet mot Israels hus; alla jordens ändar hava sett huru vår Gud frälsar.
Höjen jubel till HERREN, alla länder; bristen ut i glädjerop och lovsjungen.
Lovsjungen HERREN med harpa, med harpa och med lovsångs ljud.
Höjen jubel med trumpeter och med basuners ljud inför HERREN, konungen.
Havet bruse och allt vad däri är, jordens krets och de som bo därpå.
Strömmarna klappe i händerna, bergen juble med varandra,
inför HERREN, ty han kommer för att döma jorden.
Han skall döma jordens krets med rättfärdighet och folken med rättvisa.
HERREN är nu konung!
Därför darra folken.
Han som tronar på keruberna!
Därför skälver jorden.
HERREN är stor i Sion, och upphöjd är han över alla folk.
Därför prisar man ditt namn, det stora och fruktansvärda.
Helig är han.
Och konungen i sin makt älskar vad rätt är.
Ja, du håller rättvisa vid makt, rätt och rättfärdighet övar du i Jakob.
Upphöjen HERREN, vår Gud, och tillbedjen vid hans fotapall.
Helig är han.
Mose och Aron voro bland hans präster, och Samuel bland dem som åkallade hans namn; de ropade till HERREN, och han svarade dem.
I molnstoden talade han då till dem; de höllo hans vittnesbörd och den lag som han gav dem.
Ja, HERRE, vår Gud, du svarade dem; du var mot dem en förlåtande Gud -- och en hämnare över deras gärningar.
Upphöjen HERREN, vår Gud, och tillbedjen inför hans heliga berg.
Ty helig är HERREN, vår Gud.
En tacksägelsepsalm.
Höjen jubel till HERREN, alla länder.
Tjänen HERREN med glädje, kommen inför hans ansikte med fröjderop.
Förnimmen att HERREN är Gud.
Han har gjort oss, och icke vi själva, till sitt folk och till får i sin hjord.
Gån in i hans portar med tacksägelse, i hans gårdar med lov; tacken honom, loven hans namn.
Ty HERREN är god, hans nåd varar evinnerligen och hans trofasthet från släkte till släkte.
Av David; en psalm.
Om nåd och rätt vill jag sjunga, dig, HERRE, lovsäga.
Jag vill akta på ostrafflighetens väg -- när kommer du till mig?
Jag vill föra en ostrafflig vandel, där jag bor i mitt hus.
Jag vänder mitt öga ej till det som fördärvligt är.
Att öva orättfärdighet hatar jag; sådant skall ej låda vid mig.
Ett vrångt hjärta vare fjärran ifrån mig; vad ont är vill jag ej veta av.
Den som i hemlighet förtalar sin nästa, honom vill jag förgöra; den som har stolta ögon och högmodigt hjärta, honom lider jag icke.
Mina ögon se efter de trogna i landet, för att de må bo hos mig; den som vandrar på ostrafflighetens väg, han får vara min tjänare.
Den får icke bo i mitt hus, som övar svek; den som talar lögn skall ej bestå inför mina ögon.
Morgon efter morgon skall jag förgöra alla ogudaktiga i landet och utrota alla ogärningsmän ur HERRENS stad.
Bön av en betryckt, när han försmäktar och utgjuter sitt bekymmer inför HERREN.
HERRE, hör min bön, och låt mitt rop komma inför dig.
Dölj icke ditt ansikte för mig, när jag är i nöd.
Böj ditt öra till mig; när jag ropar, så skynda att svara mig.
Ty mina dagar hava försvunnit såsom rök, benen i min kropp äro förtorkade såsom av eld.
Mitt hjärta är förbränt såsom gräs och förvissnat; ty jag förgäter att äta mitt bröd.
För min högljudda suckans skull tränga benen i min kropp ut till huden.
Jag är lik en pelikan i öknen, jag är såsom en uggla bland ruiner.
Jag får ingen sömn och har blivit lik en ensam fågel på taket.
Hela dagen smäda mig mina fiender; de som rasa mot mig förbanna med mitt namn.
Ty jag äter aska såsom bröd och blandar min dryck med gråt,
för din vredes och förtörnelses skull, därför att du har gripit mig och kastat mig bort.
Mina dagar äro såsom skuggan, när den förlänges, och jag själv förvissnar såsom gräs.
Men du, o HERRE, tronar evinnerligen, och din åminnelse varar från släkte till släkte.
Du skall stå upp och förbarma dig över Sion; se, det är tid att du bevisar det nåd; ja, stunden har kommit.
Ty dina tjänare hava dess stenar kära och ömka sig över dess grus.
Då skola hedningarna frukta HERRENS namn och alla jordens konungar din härlighet,
när en gång HERREN har byggt upp Sion och uppenbarat sig i sin härlighet;
när han har vänt sig till de utblottades bön och upphört att förakta deras bön.
Det skall tecknas upp för ett kommande släkte, och det folk som varder skapat skall lova HERREN,
att han har blickat ned från sin heliga höjd, att HERREN har skådat från himmelen ned till jorden,
för att höra den fångnes klagan, för att befria dödens barn,
på det att man i Sion må förkunna HERRENS namn och hans lov i Jerusalem,
när alla folk församlas, och alla riken, för att tjäna HERREN.
Han har på vägen nedböjt min kraft, han har förkortat mina dagar.
Jag säger: Min Gud, tag mig icke bort i mina halva dagar, du vilkens år vara från släkte till släkte.
I urtiden lade du jordens grund, och himlarna äro dina händer verk:
de skola förgås, men du förbliver, de skola alla nötas ut såsom en klädnad; du skall förvanda dem såsom man byter om sin dräkt, och de fara hän.
Men du är densamme, och dina år skola icke hava någon ände.
Dina tjänares barn skola få bo i landet, och deras avkomma skall bestå inför dig.
Av David.
Lova HERREN, min själ, och allt det i mig är hans heliga namn.
Lova HERREN, min själ, och förgät icke vad gott han har gjort,
han som förlåter dig alla dina missgärningar och helar alla dina brister,
han som förlossar ditt liv från graven och kröner dig med nåd och barmhärtighet,
han som mättar ditt begär med sitt goda, så att du bliver ung på nytt såsom en örn.
HERREN gör rättfärdighetens verk och skaffar rätt åt alla förtryckta.
Han lät Mose se sina vägar, Israels barn sina gärningar.
Barmhärtig och nådig är HERREN, långmodig och stor i mildhet.
Han går icke ständigt till rätta och behåller ej vrede evinnerligen.
Han handlar icke med oss efter våra synder och vedergäller oss icke efter våra missgärningar.
Ty så hög som himmelen är över jorden, så väldig är hans nåd över dem som frukta honom.
Så långt som öster är från väster låter han våra överträdelser vara från oss.
Såsom en fader förbarmar sig över barnen, så förbarmar sig HERREN över dem som frukta honom.
Ty han vet vad för ett verk vi äro, han tänker därpå att vi äro stoft.
En människas dagar äro såsom gräset, hon blomstrar såsom ett blomster på marken.
När vinden går däröver, då är det icke mer, och dess plats vet icke mer därav.
Men HERRENS nåd varar från evighet till evighet över dem som frukta honom, och hans rättfärdighet intill barnbarn,
när man håller hans förbund och tänker på hans befallningar och gör efter dem.
HERREN har ställt sin tron i himmelen, och hans konungavälde omfattar allt.
Loven HERREN, I hans änglar, I starke hjältar, som uträtten hans befallning, så snart I hören ljudet av hans befallning.
Loven HERREN, I alla hans härskaror, I hans tjänare, som uträtten hans vilja.
Loven HERREN, I alla hans verk, varhelst hans herradöme är.
Min själ, lova HERREN.
Lova HERREN, min själ.
HERRE, min Gud, du är hög och stor, i majestät och härlighet är du klädd.
Du höljer dig i ljus såsom i en mantel, du spänner ut himmelen såsom ett tält;
du timrar på vattnen dina salar, molnen gör du till din vagn, och du far fram på vindens vingar.
Du gör vindar till dina sändebud, eldslågor till dina tjänare.
Du grundade jorden på hennes fästen, så att hon icke vacklar till evig tid.
Med djupet betäckte du henne såsom med en klädnad; uppöver bergen stodo vattnen.
Men för din näpst flydde de; för ljudet av ditt dunder hastade de undan.
Berg höjde sig, och dalar sänkte sig, på den plats som du hade bestämt för dem.
En gräns satte du, som vattnen ej fingo överskrida, så att de icke åter skulle betäcka jorden.
Du lät källor flyta fram i dalarna, mellan bergen togo de sin väg.
De vattna alla markens djur, vildåsnorna släcka i dem sin törst.
Vid dem bo himmelens fåglar, från trädens grenar höja de sin röst.
Du vattnar bergen från dina salar, jorden mättas av den frukt du skapar.
Du låter gräs skjuta upp för djuren och örter till människans tjänst.
Så framalstrar du bröd ur jorden
och vin, som gläder människans hjärta; så gör du hennes ansikte glänsande av olja, och brödet styrker människans hjärta.
HERRENS träd varda ock mättade, Libanons cedrar, som han har planterat;
fåglarna bygga där sina nästen, hägern gör sitt bo i cypresserna.
Stenbockarna hava fått de höga bergen, klyftorna är klippdassarnas tillflykt.
Du gjorde månen till att bestämma tiderna; solen vet stunden då den skall gå ned.
Du sänder mörker, och det bliver natt; då komma alla skogens djur i rörelse,
de unga lejonen ryta efter rov och begära sin föda av Gud.
Solen går upp; då draga de sig tillbaka och lägga sig ned i sina kulor.
Människan går då ut till sin gärning och till sitt arbete intill aftonen.
Huru mångfaldiga äro icke dina verk, o HERRE!
Med vishet har du gjort dem alla.
Jorden är full av vad du har skapat.
Se ock havet, det stora ock vida: ett tallöst vimmel rör sig däri, djur både stora och små.
Där gå skeppen sin väg fram, Leviatan, som du har skapat att leka däri.
Alla vänta de efter dig, att du skall giva dem deras mat i rätt tid.
Du giver dem, då samla de in; du upplåter din hand, då varda de mättade med goda håvor.
Du fördöljer ditt ansikte, då förskräckas de; du tager bort deras ande, då förgås de och vända åter till sitt stoft igen.
Du sänder ut din ande, då varda de skapade, och du förnyar jordens anlete.
HERRENS ära förblive evinnerligen; må HERREN glädja sig över sina verk,
han som skådar på jorden, och hon bävar, han som rör vid bergen, och de ryka.
Jag vill sjunga till HERRENS ära, så länge jag lever; jag vill lovsjunga min Gud, så länge jag är till.
Mitt tal behage honom väl; må jag själv få glädja mig i HERREN.
Men må syndare försvinna ifrån jorden och inga ogudaktiga mer vara till.
Lova HERREN, min själ Halleluja!
Tacken HERREN, åkallen hans namn, gören hans gärningar kunniga bland folken.
Sjungen till hans ära, lovsägen honom, talen om alla hans under.
Berömmen eder av hans heliga namn; glädje sig av hjärtat de som söka HERREN.
Frågen efter HERREN och hans makt, söken hans ansikte beständigt.
Tänken på de underbara verk som han har gjort, på hans under och hans muns domar,
I Abrahams, hans tjänares, säd, I Jakobs barn, hans utvalda.
Han är HERREN, vår Gud; över hela jorden gå hans domar.
Han tänker evinnerligen på sitt förbund, intill tusen släkten på vad han har stadgat,
på det förbund han slöt med Abraham och på sin ed till Isak.
Han fastställde det för Jakob till en stadga, för Israel till ett evigt förbund;
han sade: »Åt dig vill jag giva Kanaans land, det skall bliva eder arvedels lott.»
Då voro de ännu en liten hop, de voro ringa och främlingar därinne.
Och de vandrade åstad ifrån folk till folk, ifrån ett rike bort till ett annat.
Han tillstadde ingen att göra dem skada, han straffade konungar för deras skull:
»Kommen icke vid mina smorda, och gören ej mina profeter något ont.»
Och när han bjöd hungersnöd komma över landet och fördärvade allt deras livsuppehälle,
då sände han åstad en man framför dem: Josef blev såld till träl.
Man slog hans fötter i bojor, i järn fick han ligga fjättrad,
till den tid då hans ord uppfylldes, då HERRENS tal bevisade hans oskuld.
Då sände konungen och lät släppa honom lös, folkens behärskare gav honom fri.
Han satte honom till herre över sitt hus, till att råda över all hans egendom;
han skulle binda hans furstar efter sin vilja och lära hans äldste vishet.
Och Israel kom till Egypten, Jakob blev en gäst i Hams land.
Och HERREN gjorde sitt folk mycket fruktsamt och mäktigare än dess ovänner voro,
de vilkas hjärtan han vände till att hata hans folk, till att lägga onda råd mot hans tjänare.
Han sände Mose, sin tjänare, och Aron, som han hade utvalt.
De gjorde hans tecken ibland dem och under i Hams land.
Han sände mörker och lät allt bliva mörkt; och de stodo icke emot hans ord.
Han förvandlade deras vatten till blod och lät så deras fiskar dö.
Deras land kom att vimla av paddor, ända in i deras konungars kamrar.
Han bjöd, och flugsvärmar kommo, mygg i hela deras land.
Han gav dem hagel för regn, eldslågor sände han i deras land.
Och han slog deras vinträd och fikonträd och bröt sönder träden i deras land.
Han bjöd, och gräshoppor kommo, och gräsmaskar i tallös mängd.
De åto upp alla örter i deras land, de åto upp frukten på deras mark.
Och han slog allt förstfött i deras land, förstlingen av all deras kraft.
Så förde han dem ut, med silver och guld, och i hans stammar var ingen som stapplade.
Egyptierna gladde sig, när de drogo ut; ty förskräckelse för Israel hade fallit över dem.
Han bredde ut ett moln till skygd, och en eld för att lysa om natten.
De begärde, då lät han vaktlar komma, och med bröd från himmelen mättade han dem.
Han öppnade klippan, och vatten flödade; det gick genom öknen såsom en ström.
Ty han tänkte på sitt heliga ord, på sin tjänare Abraham.
Så förde han ut sitt folk med fröjd, med jubel dem som han hade utvalt.
Han gav åt dem hedningarnas länder, och folkens förvärv fingo de till besittning,
för att de skulle hålla hans stadgar och taga hans lagar i akt.
Halleluja!
Halleluja!
Tacken HERREN, ty han är god, ty hans nåd varar evinnerligen.
Vem kan uttala HERRENS väldiga gärningar och förkunna allt hans lov?
Saliga äro de som akta på vad rätt är, de som alltid öva rättfärdighet.
Tänk på mig, HERRE, efter din nåd mot ditt folk, besök mig med din frälsning,
så att jag med lust får se dina utvaldas lycka, glädja mig med ditt folks glädje, berömma mig med din arvedel.
Vi hava syndat likasom våra fäder, vi hava gjort illa, vi hava varit ogudaktiga.
Våra fäder i Egypten aktade icke på dina under; de tänkte icke på dina många nådegärningar, utan voro gensträviga vid havet, invid Röda havet.
Men han frälste dem för sitt namns skull, för att göra sin makt kunnig.
Han näpste Röda havet, så att det blev torrt, och förde dem genom djupen såsom genom en öken.
Han frälste dem från deras motståndares hand och förlossade dem ifrån fiendens hand.
Vattnet övertäckte deras ovänner; icke en enda av dem blev kvar.
Då trodde de på hans ord, då sjöngo de hans lov.
Men snart glömde de hans gärningar, de förbidade icke hans råd.
De grepos av lystnad i öknen och frestade Gud i ödemarken.
Då gav han dem vad de begärde, men sände tärande sjukdom över dem.
Och de upptändes av avund mot Mose i lägret, mot Aron, HERRENS helige.
Men jorden öppnade sig och uppslukade Datan och övertäckte Abirams hop.
Och eld begynte brinna i deras hop, en låga brände upp de ogudaktiga.
De gjorde en kalv vid Horeb och tillbådo ett gjutet beläte;
sin ära bytte de bort mot bilden av en oxe, som äter gräs.
De glömde Gud, sin frälsare, som hade gjort så stora ting i Egypten,
så underbara verk i Hams land, så fruktansvärda gärningar vid Röda havet.
Då hotade han att förgöra dem; men Mose, den man som han hade utvalt, trädde fram såsom medlare inför honom till att avvända hans vrede, så att den icke skulle fördärva.
De föraktade det ljuvliga landet och trodde icke på hans ord.
De knorrade i sina tält och lyssnade icke till HERRENS röst.
Då lyfte han upp sin hand mot dem och svor att slå ned dem i öknen,
att slå ned deras barn ibland hedningarna och förströ dem i länderna.
Och de slöto sig till Baal-Peor och åto det som var offrat åt döda.
De förtörnade Gud med sina gärningar, och en hemsökelse bröt in över dem.
Men Pinehas trädde fram och skipade rätt, och så upphörde hemsökelsen;
det vart honom räknat till rättfärdighet från släkte till släkte, för evig tid.
De förtörnade honom ock vid Meribas vatten, och det gick Mose illa för deras skull.
Ty de voro gensträviga mot hans Ande, och han talade obetänksamt med sina läppar.
De förgjorde icke de folk om vilka HERREN hade givit dem befallning,
utan beblandade sig med hedningarna och lärde sig deras gärningar.
De tjänade deras avgudar, och dessa blevo dem till en snara.
Och de offrade sina söner och döttrar till offer åt onda andar.
Ja, de utgöto oskyldigt blod, sina söners och döttrars blod och offrade dessa åt Kanaans avgudar; och landet vart ohelgat genom blodskulder.
Så blevo de orena genom sina gärningar och betedde sig trolöst i sina verk.
Då upptändes HERRENS vrede mot hans folk, och hans arvedel blev honom en styggelse.
Och han gav dem i hedningars hand, så att de som hatade dem fingo råda över dem.
Deras fiender trängde dem, och de blevo kuvade under deras hand.
Många gånger räddade han dem, men de voro gensträviga i sin egenvilja och förgingos så genom sin missgärning.
Men han såg till dem i deras nöd, när han hörde deras rop.
Och han tänkte, dem till fromma, på sitt förbund och ömkade sig efter sin stora nåd.
Och han lät dem finna barmhärtighet inför alla dem som hade fört dem i fångenskap.
Fräls oss, HERRE, vår Gud, och församla oss från hedningarna, så att vi få prisa ditt heliga namn och berömma oss av ditt lov. ----
Lovad vare HERREN, Israels Gud, från evighet till evighet!
Och allt folket säge: »Amen, Halleluja!»
Femte boken
Tacken HERREN, ty han är god, ty hans nåd varar evinnerligen.
Så säge HERRENS förlossade, de som han har förlossat ur nöden,
de som han har församlat ifrån länderna, från öster och från väster, från norr och från havssidan.
De irrade omkring i öknen på öde stigar, de funno ingen stad där de kunde bo;
de hungrade och törstade, deras själ försmäktade i dem.
Men de ropade till HERREN i sin nöd, och han räddade dem ur deras trångmål.
Och han ledde dem på en rätt väg, så att de kommo till en stad där de kunde bo.
De må tacka HERREN för hans nåd och för hans under med människors barn,
att han mättade den försmäktande själen och uppfyllde den hungrande själen med sitt goda.
De sutto i mörker och dödsskugga, fångna i elände och järnbojor,
därför att de hade varit gensträviga mot Guds ord och hade föraktat den Högstes råd.
Han kuvade deras hjärtan med olycka; de kommo på fall och hade ingen hjälpare.
Men de ropade till HERREN i sin nöd, och han frälste dem ur deras trångmål;
han förde dem ut ur mörkret och dödsskuggan, och deras bojor slet han sönder.
De må tacka HERREN för hans nåd och för hans under med människors barn,
att han krossade kopparportarna och bröt sönder järnbommarna.
De voro oförnuftiga, ty de vandrade i överträdelse, och blevo nu plågade för sina missgärningars skull;
deras själ vämjdes vid all mat, och de voro nära dödens portar.
Men de ropade till HERREN i sin nöd, och han frälste dem ur deras trångmål.
Han sände sitt ord och botade dem och räddade dem från graven.
De må tacka HERREN för hans nåd och för hans under med människors barn;
de må offra lovets offer och förtälja hans verk med jubel.
De foro på havet med skepp och drevo sin handel på stora vatten;
där fingo de se HERRENS gärningar och hans under på havsdjupet.
Med sitt ord uppväckte han stormvinden, så att den hävde upp dess böljor.
De foro upp mot himmelen, ned i djupen; deras själ upplöstes av ångest.
De raglade och stapplade såsom druckna, och all deras vishet blev till intet.
Men de ropade till HERREN i sin nöd, och han förde dem ut ur deras trångmål.
Han förbytte stormen i lugn, så att böljorna omkring dem tystnade.
Och de blevo glada att det vart stilla, och han förde dem till den hamn dit de ville.
De må tacka HERREN för hans nåd och för hans under med människors barn;
de må upphöja honom i folkets församling och lova honom där de äldste sitta.
Han gjorde strömmar till öken, källsprång till torr mark,
bördigt land till salthed, för dess inbyggares ondskas skull.
Han gjorde öknen till en vattenrik sjö och torrt land till källsprång.
Och han lät de hungrande bo där, och de byggde en stad där de kunde bo.
De besådde åkrar och planterade vingårdar, som gåvo dem sin frukt i avkastning.
Han välsignade dem, och de förökades storligen, och deras boskapshjordar lät han icke förminskas.
Väl blevo de sedan ringa och nedböjda, i det olycka och bedrövelse tryckte dem,
men han som utgjuter förakt över furstar och låter dem irra omkring i väglösa ödemarker,
han upphöjde då den fattige ur eländet och lät släkterna växa till såsom fårhjordar.
De redliga se det och glädja sig, och all orättfärdighet måste tillsluta sin mun.
Den som är vis, han akte härpå och besinne HERRENS nådegärningar.
En sång, en psalm av David.
Mitt hjärta är frimodigt, o Gud, jag vill sjunga och lova; ja, så vill min ära.
Vakna upp, psaltare och harpa; jag vill väcka morgonrodnaden.
Jag vill tacka dig bland folken, HERREN, och lovsjunga dig bland folkslagen.
Ty din nåd är stor ända uppöver himmelen, och din trofasthet allt upp till skyarna.
Upphöjd vare du, Gud, över himmelen, och över hela jorden sträcke sig din ära.
På det att dina vänner må varda räddade, må du giva seger med din högra hand och bönhöra mig.
Gud har talat i sin helgedom: »Jag skall triumfera, jag skall utskifta Sikem och skall avmäta Suckots dal.
Mitt är Gilead, mitt är Manasse, Efraim är mitt huvuds värn,
Juda min härskarstav; Moab är mitt tvagningskärl, på Edom kastar jag min sko; över filistéernas land höjer jag jubelrop.»
Vem skall föra mig till den fasta staden, vem leder mig till Edom?
Har icke du, o Gud, förkastat oss, så att du ej drager ut med våra härar, o Gud?
Giv oss hjälp mot ovännen; ty människors hjälp är fåfänglighet.
Med Gud kunna vi göra mäktiga ting; han skall förtrampa våra ovänner.
För sångmästaren; av David; en psalm.
Min lovsångs Gud, tig icke.
Ty sin ogudaktiga mun, sin falska mun hava de upplåtit mot mig, de hava talat mot mig med lögnaktig tunga.
Med hätska ord hava de omgivit mig, de hava begynt strid mot mig utan sak.
Till lön för min kärlek stå de mig emot, men jag beder allenast.
De hava bevisat mig ont för gott och hat för min kärlek.
Låt en ogudaktig man träda upp emot honom, och låt en åklagare stå på hans högra sida.
När han kommer inför rätta, må han dömas skyldig, och hans bön vare synd.
Blive hans dagar få, hans ämbete tage en annan.
Varde hans barn faderlösa och hans hustru änka.
Må hans barn alltid gå husvilla och tigga och söka sitt bröd fjärran ifrån ödelagda hem.
Må ockraren få i sin snara allt vad han äger, och må främmande plundra hans gods.
Må ingen finnas, som hyser misskund med honom, och ingen, som förbarmar sig över hans faderlösa.
Hans framtid varde avskuren, i nästa led vare sådanas namn utplånat.
Hans fäders missgärning varde ihågkommen inför HERREN, och hans moders synd varde icke utplånad.
Må den alltid stå inför HERRENS ögon; ja, sådana mäns åminnelse må utrotas från jorden.
Ty han tänkte ju icke på att öva misskund, utan förföljde den som var betryckt och fattig och den vilkens hjärta var bedrövat, för att döda dem.
Han älskade förbannelse, och den kom över honom; han hade icke behag till välsignelse, och den blev fjärran ifrån honom.
Han klädde sig i förbannelse såsom i en klädnad, och såsom vatten trängde den in i hans liv och såsom olja in i hans ben.
Den varde honom såsom en mantel att hölja sig i, och såsom en gördel att alltid omgjorda sig med.
Detta vare mina motståndares lön från HERREN, och deras som tala ont mot min själ.
Men du, HERRE, Herre, stå mig bi för ditt namn skull; god är ju din nåd, så må du då rädda mig.
Ty jag är betryckt och fattig, och mitt hjärta är genomborrat i mitt bröst.
Såsom skuggan, när den förlänges, går jag bort; jag ryckes bort såsom en gräshoppssvärm.
Mina knän äro vacklande av fasta, och min kropp förlorar sitt hull.
Till smälek har jag blivit inför dem; när de se mig, skaka de huvudet.
Hjälp mig, HERRE, min Gud; fräls mig efter din nåd;
och må de förnimma att det är din hand, att du, HERRE, har gjort det.
Om de förbanna, så välsigna du; om de resa sig upp, så komme de på skam, men må din tjänare få glädja sig.
Mina motståndare varde klädda i blygd och höljda i skam såsom i en mantel.
Min mun skall storligen tacka HERREN; mitt ibland många vill jag lova honom.
Ty han står på den fattiges högra sida för att frälsa honom från dem som fördöma hans själ.
Av David; en psalm.
HERREN sade till min herre: »Sätt dig på min högra sida, till dess jag har lagt dina fiender dig till en fotapall.»
Din makts spira skall HERREN utsträcka från Sion; du skall härska mitt ibland dina fiender.
Villigt kommer ditt folk, när du samlar din här; i helig skrud kommer din unga skara inför dig, såsom daggen kommer ur morgonrodnadens sköte.
HERREN har svurit och skall icke ångra sig: »Du är en präst till evig tid efter Melki-Sedeks sätt.»
Herren är på din högra sida, han skall krossa konungar på sin vredes dag.
Han skall hålla dom bland hedningarna, överallt skola döda ligga; han skall sönderkrossa huvuden vida omkring på jorden.
Ur bäcken skall han dricka på vägen; därför skall han upplyfta huvudet.
Halleluja!
Jag vill tacka HERREN av allt hjärta i de rättsinnigas råd och församling.
Stora äro HERRENS verk, de begrundas av alla som hava sin lust i dem.
Majestät och härlighet är vad han gör, och hans rättfärdighet förbliver evinnerligen.
Han har så gjort, att hans under äro i åminnelse; nådig och barmhärtig är HERREN.
Han giver mat åt dem som frukta honom, han tänker evinnerligen på sitt förbund.
Sina gärningars kraft har han gjort kunnig för sitt folk, i det han gav dem hedningarnas arvedel.
Hans händers verk äro trofasthet och rätt, oryggliga äro alla hans ordningar.
De stå fasta för alltid och för evigt, de fullbordas med trofasthet och rättvisa.
Han har sänt sitt folk förlossning, han har stadgat sitt förbund för evig tid; heligt och fruktansvärt är hans namn.
HERRENS fruktan är vishetens begynnelse, ett gott förstånd få alla de som göra därefter.
Hans lov förbliver evinnerligen.
Halleluja!
Säll är den man som fruktar HERREN och har sin stora lust i hans bud.
Hans efterkommande skola bliva väldiga på jorden; de redligas släkte skall varda välsignat.
Gods och rikedom skall finnas i hans hus, och hans rättfärdighet består evinnerligen.
För de redliga går han upp såsom ett ljus i mörkret, nådig och barmhärtig och rättfärdig.
Väl den som är barmhärtig och giver lån, den som stöder all sin sak på rätt!
Ty han skall icke vackla till evig tid; den rättfärdige skall vara i evig åminnelse.
För ont budskap fruktar han icke; hans hjärta är frimodigt, det förtröstar på HERREN.
Hans hjärta är fast, det fruktar icke, till dess han får se med lust på sina ovänner.
Han utströr, han giver åt de fattiga, hans rättfärdighet förbliver evinnerligen; hans horn skall varda upphöjt med ära.
Den ogudaktige skall se det och harmas; han skall bita sina tänder samman och täras bort.
Vad de ogudaktiga önska bliver till intet.
Halleluja!
Loven, I HERRENS tjänare, loven HERRENS namn.
Välsignat vare HERRENS namn från nu och till evig tid.
Från solens uppgång ända till dess nedgång vare HERRENS namn högtlovat.
HERREN är hög över alla folk, hans ära når över himmelen.
Ja, vem är såsom HERREN, vår Gud, han som sitter så högt,
han som ser ned så djupt -- ja, vem i himmelen och på jorden?
Han som upprättar den ringe ur stoftet, han som lyfter den fattige ur dyn,
för att sätta honom bredvid furstar, bredvid sitt folks furstar;
han som låter den ofruktsamma hustrun sitta med glädje såsom moder, omgiven av barn!
Halleluja!
När Israel drog ut ur Egypten, Jakobs hus ut ifrån folket med främmande tunga,
då vart Juda hans helgedom, Israel hans herradöme.
Havet såg det och flydde, Jordan vände tillbaka.
Bergen hoppade såsom vädurar, höjderna såsom lamm.
Varför flyr du undan, du hav?
Du Jordan, varför vänder du tillbaka?
I berg, varför hoppen I såsom vädurar, I höjder, såsom lamm?
För Herren må du väl bäva, du jord, för Jakobs Guds ansikte,
för honom som förvandlar klippan till en vattenrik sjö, hårda stenen till en vattenkälla.
Icke åt oss, HERRE, icke åt oss, utan åt ditt namn giv äran, för din nåds, för din sannings skull.
Varför skulle hedningarna få säga: »Var är nu deras Gud?»
Vår Gud är ju i himmelen; han kan göra allt vad han vill.
Men deras avgudar äro silver och guld, verk av människohänder.
De hava mun och tala icke, de hava ögon och se icke,
de hava öron och höra icke, de hava näsa och lukta icke.
Med sina händer taga de icke, med sina fötter gå de icke; de hava intet ljud i sin strupe.
De som hava gjort dem skola bliva dem lika, ja, alla som förtrösta på dem.
I av Israel, förtrösten på HERREN.
Ja, han är deras hjälp och sköld.
I av Arons hus, förtrösten på HERREN.
Ja, han är deras hjälp och sköld.
I som frukten HERREN, förtrösten på HERREN.
Ja, han är deras hjälp och sköld.
HERREN har tänkt på oss, han skall välsigna, han skall välsigna Israels hus, han skall välsigna Arons hus,
han skall välsigna dem som frukta HERREN, de små såväl som de stora.
Ja, HERREN föröke eder, seder själva och edra barn.
Varen välsignade av HERREN, av honom som har gjort himmel och jord.
Himmelen är HERRENS himmel, och jorden har han givit åt människors barn.
De döda prisa icke HERREN, ingen som har farit ned i det tysta.
Men vi, vi skola lova HERREN från nu och till evig tid.
Halleluja!
Jag har HERREN kär, ty han hör min röst och mina böner.
Ja, han har böjt sitt öra till mig; i hela mitt liv skall jag åkalla honom.
Dödens band omvärvde mig, och dödsrikets ångest grep mig; jag kom i nöd och bedrövelse.
Men jag åkallade HERRENS namn: »Ack HERRE, rädda min själ.»
HERREN är nådig och rättfärdig, vår Gud är barmhärtig.
HERREN bevarar de enfaldiga; jag var i elände, och han frälste mig.
Vänd nu åter till din ro, min själ, ty HERREN har gjort väl mot dig.
Ja, du har räddat min själ från döden, mitt öga från tårar, min fot ifrån fall;
jag skall få vandra inför HERREN i de levandes land.
Jag tror, ty därför talar jag, jag som var storligen plågad,
jag som måste säga i min ångest: »Alla människor äro lögnaktiga.»
Huru skall jag vedergälla HERREN alla hans välgärningar mot mig?
Jag vill taga frälsningens bägare och åkalla HERRENS namn.
Jag vill infria åt HERREN mina löften, ja, i hela hans folks åsyn.
Dyrt aktad i HERRENS ögon är hans frommas död.
Ack HERRE, jag är ju din tjänare, jag är din tjänare, din tjänarinnas son; du har lossat mina band.
Dig vill jag offra lovets offer, och HERRENS namn vill jag åkalla.
Jag vill infria åt HERREN mina löften, ja, i hela hans folks åsyn,
i gårdarna till HERRENS hus, mitt i dig, Jerusalem.
Halleluja!
Loven HERREN, alla hedningar, prisen honom, alla folk.
Ty hans nåd är väldig över oss, och HERRENS sanning varar i evighet.
Halleluja!
Tacken HERREN, ty han är god, ty hans nåd varar evinnerligen.
Så säge Israel, ty hans nåd varar evinnerligen.
Så säge Arons hus, ty hans nåd varar evinnerligen.
Så säge de som frukta HERREN, ty hans nåd varar evinnerligen.
I mitt trångmål åkallade jag HERREN, och HERREN svarade mig och ställde mig på rymlig plats.
HERREN står mig bi, jag skall icke frukta; vad kunna människor göra mig?
HERREN står mig bi, han är min hjälpare, och jag skall få se med lust på dem som hata mig.
Bättre är att taga sin tillflykt till HERREN än att förlita sig på människor.
Bättre är att taga sin tillflykt till HERREN än att förlita sig på furstar.
Alla hedningar omringa mig, men i HERRENS namn skall jag förgöra dem.
De omringa mig, ja, de omringa mig, men i HERRENS namn skall jag förgöra dem.
De omringa mig såsom bin, men de slockna såsom eld i törne; i HERRENS namn skall jag förgöra dem.
Man stöter mig hårdeligen, för att jag skall falla, men HERREN hjälper mig.
HERREN är min starkhet och min lovsång, och han blev mig till frälsning.
Man sjunger med jubel om frälsning i de rättfärdigas hyddor: »HERRENS högra hand gör mäktiga ting.
HERRENS högra han upphöjer, HERRENS högra hand gör mäktiga ting.»
Jag skall icke dö, utan leva och förtälja HERRENS gärningar.
Väl tuktade mig HERREN, men han gav mig icke åt döden.
Öppnen för mig rättfärdighetens portar; jag vill gå in genom dem och tacka HERREN.
Detta är HERRENS port, de rättfärdiga skola gå in genom den.
Jag tackar dig för att du svarade mig och blev mig till frälsning.
Den sten som byggningsmännen förkastade har blivit en hörnsten.
Av HERREN har den blivit detta; underbart är det i våra ögon.
Detta är den dag som HERREN har gjort; låtom oss på den fröjdas och vara glada.
Ack HERRE, fräls!
Ack HERRE, låt väl gå!
Välsignad vare han som kommer, i HERRENS namn.
Vi välsigna eder från HERRENS hus.
HERREN är Gud, och han gav oss ljus.
Ordnen eder i högtidsled, med lövrika kvistar i händerna, fram till altarets horn.
Du är min Gud, och jag vill tacka dig; min Gud, jag vill upphöja dig.
Tacka HERREN, ty han är god, ty hans nåd varar evinnerligen.
Saliga äro de vilkas väg är ostrafflig, de som vandra efter HERRENS lag.
Saliga äro de som taga hans vittnesbörd i akt, de som av allt hjärta söka honom,
de som icke göra vad orätt är, utan vandra på hans vägar.
Du har givit befallningar, för att de skola hållas med all flit.
O att mina vägar vore rätta, så att jag hölle dina stadgar!
Då skulle jag icke komma på skam, när jag skådade på alla dina bud.
Jag vill tacka dig av uppriktigt hjärta, när jag får lära din rättfärdighets rätter.
Dina stadgar vill jag hålla; övergiv mig icke så helt och hållet.
Huru skall en yngling bevara sin väg obesmittad?
När han håller sig efter ditt ord.
Jag söker dig av allt mitt hjärta; låt mig icke fara vilse från dina bud.
Jag gömmer ditt tal i mitt hjärta, för att jag icke skall synda mot dig.
Lovad vare du, HERRE!
Lär mig dina stadgar.
Med mina läppar förtäljer jag alla din muns rätter.
Jag fröjdar mig över dina vittnesbörds väg såsom över alla skatter.
Jag vill begrunda dina befallningar och skåda på dina stigar.
Jag har min lust i dina stadgar, jag förgäter icke ditt ord.
Gör väl mot din tjänare, så att jag får leva, då vill jag hålla ditt ord.
Öppna mina ögon, så att jag kan skåda undren i din lag.
Jag är en främling på jorden; fördölj icke dina bud för mig.
Min själ är sönderkrossad av ständig trängtan efter dina rätter.
Du näpser de fräcka, de förbannade, dem som fara vilse från dina bud.
Tag bort ifrån mig smälek och förakt, ty jag tager i akt dina vittnesbörd.
Ja, furstar sitta och lägga råd mot mig, men din tjänare begrundar dina stadgar;
ja, dina vittnesbörd äro min lust, de äro mina rådgivare.
Min själ ligger nedtryckt i stoftet; behåll mig vid liv efter ditt ord.
Jag förtäljde om mina vägar, och du svarade mig; lär mig dina stadgar.
Lär mig att förstå dina befallningars väg, så vill jag begrunda dina under.
Min själ gråter av bedrövelse; upprätta mig efter ditt ord.
Låt lögnens väg vara fjärran ifrån mig, och förunna mig din undervisning.
Jag har utvalt sanningens väg, dina rätter har jag ställt framför mig.
Jag håller mig till dina vittnesbörd; HERRE, låt mig icke komma på skam.
Jag vill löpa dina buds väg, ty du tröstar mitt hjärta.
Visa mig, HERRE, dina stadgars väg, så vill jag taga den i akt intill änden.
Giv mig förstånd, så vill jag taga din lag i akt och hålla den av allt hjärta.
Led mig på dina buds stig, ty till den har jag behag.
Böj mitt hjärta till dina vittnesbörd, och låt det icke vika av till orätt vinning.
Vänd bort mina ögon, så att de icke se efter fåfänglighet; behåll mig vid liv på dina vägar.
Uppfyll på din tjänare ditt tal, ty det leder till din fruktan.
Vänd bort ifrån mig den smälek som jag fruktar; ty dina rätter äro goda.
Se, jag längtar efter dina befallningar; behåll mig vid liv genom din rättfärdighet.
Din nåd komme över mig, HERRE, din frälsning efter ditt tal;
Så kan jag giva den svar, som smädar mig; ty jag förtröstar på ditt ord.
Ryck icke sanningens ord så helt och hållet bort ifrån min mun, ty jag hoppas på dina domar.
Så vill jag hålla din lag beständigt, ja, alltid och evinnerligen.
Låt mig gå fram på rymlig plats, ty jag begrundar dina befallningar.
Jag vill tala om dina vittnesbörd inför konungar, och jag skall icke komma på skam.
Jag vill hava min lust i dina bud, ty de äro mig kära;
jag vill lyfta mina händer upp till dina bud, ty de äro mig kära, och jag vill begrunda dina stadgar.
Tänk på ordet till din tjänare, eftersom du har givit mig hopp.
Det är min tröst i mitt lidande att ditt tal behåller mig vid liv.
De fräcka bespotta mig övermåttan; likväl viker jag icke ifrån din lag.
Jag tänker på dina domar i forna tider, HERRE, och jag varder tröstar.
Glödande harm griper mig för de ogudaktigas skull, därför att de övergiva din lag.
Dina stadgar äro lovsånger för mig i det hus där jag dväljes.
Jag tänker om natten på ditt namn, HERRE, och jag håller din lag.
Detta har blivit mig beskärt: att jag får taga dina befallningar i akt.
Min del är HERREN; jag har beslutit att hålla dina ord.
Jag bönfaller inför dig av allt hjärta; var mig nådig efter ditt tal.
Jag betänker mina vägar och vänder mina fötter till dina vittnesbörd.
Jag skyndar mig och dröjer icke att hålla dina bud.
De ogudaktigas snaror omgiva mig, men jag förgäter icke din lag.
Mitt i natten står jag upp för att tacka dig för din rättfärdighets rätter.
Jag sluter mig till alla dem som frukta dig och till dem som hålla dina befallningar.
Jorden är full av din nåd, o HERRE; lär mig dina stadgar.
Du gör din tjänare gott, HERRE, efter ditt ord.
Lär mig gott förstånd och kunskap, ty jag tror på dina bud.
Förrän jag fick lida, for jag vilse, men nu håller jag mig vid ditt tal.
Du är god och gör vad gott är; lär mig dina stadgar.
De fräcka hopspinna lögn mot mig, men jag vill av allt hjärta taga dina befallningar i akt.
Deras hjärtan äro okänsliga såsom fett, men jag har min lust i din lag.
Det var mig gott att jag vart tuktad, så att jag fick lära mig dina stadgar.
Din muns lag är mig bättre än tusentals stycken guld och silver.
Dina händer hava gjort och berett mig; giv mig förstånd, så att jag kan lära dina bud.
De som frukta dig skola se mig och glädjas, ty jag hoppas på ditt ord.
HERRE, jag vet att dina domar äro rättfärdiga, och att du har tuktat mig i trofasthet.
Din nåd vare min tröst, såsom du har lovat din tjänare.
Din barmhärtighet komme över mig, så att jag får leva; ty din lag är min lust.
På skam komme de fräcka, ty de hava gjort mig orätt utan sak; men jag vill begrunda dina befallningar.
Till mig må de vända sig, som frukta dig, och de om känna dina vittnesbörd.
Mitt hjärta vare ostraffligt i dina stadgar, så att jag icke kommer på skam.
Min själ trängtar efter din frälsning, jag hoppas på ditt ord.
Mina ögon trängta efter ditt tal, och jag säger: »När vill du trösta mig?»
Ty jag är såsom en vinlägel i rök, men jag förgäter icke dina stadgar.
Huru få äro icke din tjänares dagar!
När vill du hålla dom över mina förföljare?
De fräcka gräva gropar för mig, de som icke leva efter din lag.
Alla dina bud äro sanning; utan sak förföljer man mig; hjälp mig.
De hava så när fördärvat mig på jorden, fastän jag icke har övergivit dina befallningar.
Behåll mig vid liv efter din nåd, så vill jag hålla din muns vittnesbörd.
Evinnerligen, HERRE, står ditt ord fast i himmelen.
Från släkte till släkte varar din trofasthet; du har grundat jorden, och den består.
Till att utföra dina rätter består allt än i dag, ty allting måste tjäna dig.
Om din lag icke hade varit min lust, så hade jag förgåtts i mitt elände.
Aldrig skall jag förgäta dina befallningar, ty genom dem har du behållit mig vid liv.
Jag är din, fräls mig; ty jag begrundar dina befallningar.
På mig vakta de ogudaktiga för att förgöra mig; men jag aktar på dina vittnesbörd.
På all annan fullkomlighet har jag sett en ände, men ditt bud är omätligt i vidd.
Huru kär har jag icke din lag!
Hela dagen begrundar jag den.
Visare än mina fiender äro, göra mig dina bud, ty de tillhöra mig för evig tid.
Jag är klokare än alla mina lärare, ty jag begrundar dina vittnesbörd.
Jag är förståndigare än de gamle, ty jag tager dina befallningar i akt.
Jag avhåller mina fötter ifrån alla onda vägar, för att jag må hålla ditt ord.
Jag viker icke ifrån dina rätter, ty du undervisar mig.
Huru ljuvt för min tunga är icke ditt tal!
Det är ljuvare än honung för min mun.
Av dina befallningar får jag förstånd; därför hatar jag alla lögnens vägar.
Ditt ord är mina fötters lykta och ett ljus på min stig.
Jag har svurit och hållit det: att taga din rättfärdighets rätter i akt.
Jag är storligen plågad; HERRE, behåll mig vid liv efter ditt ord.
Låt min muns frivilliga offer behaga dig, HERRE, och lär mig dina rätter.
Jag bär min själ alltid i min hand, men jag förgäter icke din lag.
De ogudaktiga lägga ut snaror för mig, men jag far icke vilse från dina befallningar.
Jag har dina vittnesbörd till min eviga arvedel, ty de äro mitt hjärtas fröjd.
Jag har böjt mitt hjärta till att göra efter dina stadgar, alltid och intill änden.
Jag hatar dem som halta på båda sidor, men din lag har jag kär.
Du är mitt beskärm och min sköld; jag hoppas på ditt ord.
Viken bort ifrån mig, I onde; jag vill taga min Guds bud i akt.
Uppehåll mig efter ditt tal, så att jag får leva, och låt mig icke komma på skam med mitt hopp.
Stöd mig, så att jag varder frälst, så vill jag alltid se med lust på dina stadgar.
Du aktar för intet alla som fara vilse från dina stadgar, ty förgäves är deras svek.
Du förkastar såsom slagg alla ogudaktiga på jorden; därför har jag dina vittnesbörd kära.
Av fruktan för dig ryser mitt kött, och jag rädes för dina domar.
Jag övar rätt och rättfärdighet; du skall icke överlämna mig åt mina förtryckare.
Tag dig an din tjänares sak, och låt det gå honom väl; låt icke de fräcka förtrycka mig.
Mina ögon trängta efter din frälsning och efter din rättfärdighets tal.
Gör med din tjänare efter din nåd, och lär mig dina stadgar.
Jag är din tjänare; giv mig förstånd, så att jag kan känna dina vittnesbörd.
Det är tid för HERREN att handla, ty de hava gjort din lag om intet.
Därför har jag dina bud kära mer än guld, jag, mer än fint guld.
Därför håller jag alla dina befallningar i allo för rätta, men alla lögnens vägar hatar jag.
Underbara äro dina vittnesbörd, därför tager min själ dem i akt.
När dina ord upplåtas, giva de ljus och skänka förstånd åt de enfaldiga.
Jag spärrar upp min mun och flämtar, ty jag längtar ivrigt efter dina bud.
Vänd dig till mig och var mig nådig, såsom rätt är mot dem som hava ditt namn kärt.
Gör mina steg fasta genom ditt tal, och låt ingen orätt varda mig övermäktig.
Förlossa mig från människors förtryck, så vill jag hålla dina befallningar.