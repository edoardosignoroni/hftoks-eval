Och alla som kommo till honom tog han emot;
och han predikade om Guds rike och undervisade om Herren Jesus Kristus med all frimodighet, utan att någon hindrade honom däri.
Paulus, Jesu Kristi tjänare, kallad till apostel, avskild till att förkunna Guds evangelium,
vilket Gud redan förut genom sina profeter hade i heliga skrifter utlovat,
evangelium om hans Son, vilken såsom människa i köttet är född av Davids säd
och såsom helig andevarelse är med kraft bevisad vara Guds Son, allt ifrån uppståndelsen från de döda, ja, evangelium om Jesus Kristus, vår Herre,
genom vilken vi hava fått nåd och apostlaämbete för att, hans namn till ära, upprätta trons lydnad bland alla hednafolk,
bland vilka jämväl I ären, I som ären kallade och Jesu Kristi egna --
jag, Paulus, hälsar alla Guds älskade som bo i Rom, dem som äro kallade och heliga.
Nåd vare med eder och frid ifrån Gud, vår Fader, och Herren Jesus Kristus.
Först och främst tackar jag min Gud genom Jesus Kristus för eder alla, därför att man i hela världen talar om eder tro.
Ty Gud, som jag i min ande tjänar såsom förkunnare av evangelium om hans Son, han är mitt vittne, han vet huru oavlåtligt jag tänker på eder
och i mina böner alltid beder att jag dock nu omsider må få ett gynnsamt tillfälle att komma till eder, om Gud så vill.
Ty jag längtar efter att se eder, för att jag må kunna meddela eder någon andlig nådegåva till att styrka eder;
jag menar: för att jag i eder krets må tillsammans med eder få hämta hugnad ur vår gemensamma tro, eder och min.
Jag vill säga eder, mina bröder, att jag ofta har haft i sinnet att komma till eder, för att också bland eder få skörda någon frukt, såsom bland övriga hednafolk; dock har jag allt hittills blivit hindrad.
Både mot greker och mot andra folk, både mot visa och mot ovisa har jag förpliktelser.
Därför är jag villig att förkunna evangelium också för eder som bon i Rom.
Ty jag blyges icke för evangelium; ty det är en Guds kraft till frälsning för var och en som tror, först och främst för juden, så ock för greken.
Rättfärdighet från Gud uppenbaras nämligen däri, av tro till tro; så är ock skrivet: »Den rättfärdige skall leva av tro.»
Ty Guds vrede uppenbarar sig från himmelen över all ogudaktighet och orättfärdighet hos människor som i orättfärdighet undertrycka sanningen.
Vad man kan känna om Gud är nämligen uppenbart bland dem; Gud har ju uppenbarat det för dem.
Ty hans osynliga väsen, hans eviga makt och gudomshärlighet hava ända ifrån världens skapelse varit synliga, i det att de kunna förstås genom hans verk.
Så äro de då utan ursäkt.
Ty fastän de hade lärt känna Gud, prisade och tackade de honom dock icke såsom Gud, utan förföllo till fåfängliga tankar; och så blevo deras oförståndiga hjärtan förmörkade.
När de berömde sig av att vara visa, blevo de dårar
och bytte bort den oförgänglige Gudens härlighet mot beläten, som voro avbilder av förgängliga människor, ja ock av fåglar och fyrfotadjur och krälande djur.
Därför prisgav Gud dem i deras hjärtans begärelser åt orenhet, så att de med varandra skändade sina kroppar.
De hade ju bytt bort Guds sanning mot lögn och tagit sig för att dyrka och tjäna det skapade framför Skaparen, honom som är högtlovad i evighet, amen.
Fördenskull gav Gud dem till pris åt skamliga lustar: deras kvinnor utbytte det naturliga umgänget mot ett onaturligt;
sammalunda övergåvo ock männen det naturliga umgänget med kvinnan och upptändes i lusta till varandra och bedrevo styggelse, man med man.
Så fingo de på sig själva uppbära sin villas tillbörliga lön.
Och eftersom de icke hade aktat det något värt att taga vara på sin kunskap om Gud, gav Gud dem till pris åt ett ovärdigt sinnelag, till att bedriva otillbörliga ting.
Så hava de blivit uppfyllda av allt slags orättfärdighet, ondska, girighet, elakhet; de äro fulla av avund, mordlust, trätlystnad, svek, vrångsinthet;
de äro örontasslare, förtalare, styggelser för Gud, våldsverkare, övermodiga, stortaliga, illfundiga, olydiga mot sina föräldrar,
oförståndiga, trolösa, utan kärlek till sina egna, utan barmhärtighet mot andra.
Och fastän de väl veta vad Gud har stadgat såsom rätt, att nämligen de som handla så förtjäna döden, är det dem icke nog att själva så göra, de giva ock sitt bifall åt andra som handla likaså.
Därför är du utan ursäkt, du människa, vem du än är, som dömer.
Ty därmed att du dömer en annan fördömer du dig själv, eftersom du, som dömer den andre, själv handlar på samma sätt.
Och vi veta att Guds dom verkligen kommer över dem som handla så.
Men du menar väl detta, att du skall kunna undfly Guds dom, du människa, som dömer dem som handla så, och dock gör detsamma som de?
Eller föraktar du hans godhets, skonsamhets och långmodighets rikedom, utan att förstå att denna Guds godhet vill föra dig till bättring?
Genom din hårdhet och ditt hjärtas obotfärdighet samlar du ju över dig vrede, som skall drabba dig på vredens dag, då när det bliver uppenbart att Gud är en rättvis domare.
Ty »han skall vedergälla var och en efter hans gärningar».
Evigt liv skall han giva åt dem som med uthållighet i att göra det goda söka härlighet och ära och oförgänglighet.
Men över dem som äro genstridiga och icke lyda sanningen, utan lyda orättfärdigheten, över dem kommer vrede och förtörnelse.
Ja, bedrövelse och ångest skall komma över den människas själ, som gör det onda, först och främst över judens, så ock över grekens.
Men härlighet och ära och frid skall tillfalla var och en som gör det goda, först och främst juden, så ock greken.
Ty hos Gud finnes intet anseende till personen;
alla de som utan lag hava syndat skola ock utan lag förgås, och alla de som med lag hava syndat skola genom lag bliva dömda.
Ty icke lagens hörare äro rättfärdiga inför Gud, men lagens görare skola förklaras rättfärdiga.
Ty då hedningarna, som icke hava lag, av naturen göra vad lagen innehåller, så äro dessa, utan att hava lag, sig själv en lag,
då de ju sålunda visa att lagens verk äro skrivna i deras hjärtan.
Därom utgöra också deras egna samveten ett vittnesbörd, så ock, i den inbördes umgängelsen, deras tankar, när dessa anklaga eller ock försvara dem.
Ja, så skall det befinnas vara på den dag då Gud, enligt det evangelium jag förkunnar, genom Kristus Jesus dömer över vad som är fördolt hos människorna.
Du kallar dig jude och förlitar dig på lagen och berömmer dig av Gud.
Du känner ock hans vilja, och eftersom du har fått din undervisning ur lagen, kan du döma om vad rättast är;
och du tilltror dig att vara en ledare för blinda, ett ljus för människor som vandra i mörker,
en uppfostrare för oförståndiga, en lärare för enfaldiga, eftersom du i lagen har uttrycket för kunskapen och sanningen.
Du som vill lära andra, du lär icke dig själv!
Du som predikar att man icke skall stjäla, du begår själv stöld!
Du som säger att man icke skall begå äktenskapsbrott, du begår själv sådant brott!
Du som håller avgudarna för styggelser, du gör dig själv skyldig till tempelrån!
Du som berömmer dig av lagen, du vanärar Gud genom att överträda lagen,
ty, såsom det är skrivet, »för eder skull varder Guds namn smädat bland hedningarna».
Ty väl är omskärelse till gagn, om du håller lagen; men om du är en lagöverträdare, så är du med din omskärelse dock oomskuren.
Om nu den oomskurne håller lagens stadgar, skall han då icke, fastän han är oomskuren, räknas såsom omskuren?
Jo, och han som i följd av sin härkomst är oomskuren, men ändå fullgör lagen, skall bliva dig till dom, dig som äger lagens bokstav och omskärelsen, men likväl är en lagöverträdare.
Ty den är icke jude, som är det i utvärtes måtto, ej heller är det omskärelse, som sker utvärtes på köttet.
Nej, den är jude, som är det i invärtes måtto, och omskärelse är hjärtats omskärelse, en som sker i Anden, och icke i kraft av bokstaven; och han har sin berömmelse, icke från människor, utan från Gud.
Vilket företräde hava då judarna, eller vad gagn hava de av omskärelsen?
Jo, ett stort företräde, på allt sätt; först och främst det, att de hava blivit betrodda med Guds löftesord.
Ty vad betyder det, om några av dem blevo trolösa?
Kan då deras trolöshet göra Guds trofasthet om intet?
Bort det!
Må Gud stå såsom sannfärdig, om ock »var människa är en lögnare».
Så är ju skrivet: »På det att du må finnas rättfärdig i dina ord och få rätt, när man sätter sig till doms över dig.»
Men är det nu så, att vår orättfärdighet tjänar till att bevisa Guds rättfärdighet, vad skola vi då säga?
Kan väl Gud, han som låter vredesdomen drabba, vara orättfärdig?
(Jag talar såsom vore det fråga om en människa.)
Bort det!
Huru skulle Gud då kunna döma världen?
Och å andra sidan, om Guds sannfärdighet genom min lögnaktighet ännu mer har trätt i dagen, honom till ära, varför skall då jag likväl dömas såsom syndare?
Och varför skulle vi icke »göra vad ont är, för att gott måtte komma därav», såsom man, för att smäda oss, påstår att vi göra, och såsom några föregiva att vi lära? -- Sådana få med rätta sin dom.
Huru är det alltså?
Äro vi då något förmer än de andra?
Ingalunda.
Redan härförut har jag ju måst anklaga både judar och greker för att allasammans vara under synd.
Så är ock skrivet: »Ingen rättfärdig finnes, icke en enda.
Ingen förståndig finnes, ingen finnes som söker Gud.
Nej, alla hava de avvikit, allasammans hava de blivit odugliga, ingen finnes som gör vad gott är, det finnes ingen enda.
En öppen grav är deras strupe, sina tungor bruka de till svek.
Huggormsgift är inom deras läppar.
Deras mun är full av förbannelse och bitterhet.
Deras fötter äro snara, när det gäller att utgjuta blod.
Förödelse och elände är på deras vägar,
och fridens väg känna de icke.
Guds fruktan är icke för deras ögon.»
Nu veta vi att allt vad lagen säger, det talar den till dem som hava lagen, för att var mun skall bliva tillstoppad och hela världen stå med skuld inför Gud;
ty av laggärningar bliver intet kött rättfärdigt inför honom.
Vad som kommer genom lagen är kännedom om synden.
Men nu har, utan lag, en rättfärdighet från Gud blivit uppenbarad, en som lagen och profeterna vittna om,
en rättfärdighet från Gud genom tro på Jesus Kristus, för alla dem som tro.
Ty här är ingen åtskillnad.
Alla hava ju syndat och äro i saknad av härligheten från Gud;
och de bliva rättfärdiggjorda utan förskyllan, av hans nåd, genom förlossningen i Kristus Jesus,
honom som Gud har ställt fram såsom ett försoningsmedel genom tro, i hans blod.
Så ville Gud -- då han i sin skonsamhet hade haft fördrag med de synder som förut hade blivit begångna -- nu visa att han dock var rättfärdig.
Ja, så ville han i den tid som nu är lämna beviset för att han är rättfärdig.
Härigenom skulle han både själv befinnas vara rättfärdig och göra den rättfärdig, som låter det bero på tro på Jesus.
Huru bliver det då med vår berömmelse?
Den är utestängd.
Genom vilken lag?
Månne genom en gärningarnas lag?
Nej, genom en trons lag.
Vi hålla nämligen före att människan bliver rättfärdig genom tro, utan laggärningar.
Eller är Gud allenast judarnas Gud?
Är han icke ock hedningarnas?
Jo, förvisso också hedningarnas,
så visst som Gud är en, han som skall göra de omskurna rättfärdiga av tro, så ock de oomskurna genom tron.
Göra vi då vad lag är om intet genom tron?
Bort det!
Vi göra tvärtom lag gällande.
Vad skola vi då säga om Abraham, vår stamfader efter köttet?
Om Abraham blev rättfärdig av gärningar, så har han ju något att berömma sig av.
Dock icke inför Gud.
Ty vad säger skriften? »Abraham trodde Gud, och det räknades honom till rättfärdighet.»
Den som håller sig till gärningar, honom bliver lönen tillräknad icke på grund av nåd, utan på grund av förtjänst.
Men den som icke håller sig till gärningar, utan tror på honom som gör den ogudaktige rättfärdig, honom räknas hans tro till rättfärdighet.
Så prisar ock David den människa salig, som Gud tillräknar rättfärdighet, utan gärningar:
»Saliga äro de vilkas överträdelser äro förlåtna, och vilkas synder äro överskylda.
Salig är den man som Herren icke tillräknar synd.»
Gäller nu detta ordet »salig» de omskurna allenast eller ock de oomskurna?
Vi säga ju att »tron räknades Abraham till rättfärdighet».
Huru blev den honom då tillräknad?
Skedde det sedan han hade blivit omskuren, eller medan han ännu var oomskuren?
Det skedde icke sedan han hade blivit omskuren, utan medan han ännu var oomskuren.
Och han undfick omskärelsens tecken såsom ett insegel på den rättfärdighet genom tron, som han hade, medan han ännu var oomskuren.
Ty så skulle han bliva en fader för alla oomskurna som tro, och så skulle rättfärdighet tillräknas dem.
Han skulle ock bliva en fader för omskurna, nämligen för sådana som icke allenast äro omskurna, utan ock vandra i spåren av den tro som vår fader Abraham hade, medan han ännu var oomskuren.
Det var nämligen icke genom lag som Abraham och hans säd undfick det löftet att han skulle få världen till arvedel; det var genom rättfärdighet av tro.
Ty om de som låta det bero på lag skola få arvedelen, så är tron till intet nyttig, och löftet är gjort om intet.
Vad lagen kommer åstad är ju vredesdom; men där ingen lag finnes, där finnes icke heller någon överträdelse.
Därför måste det bero på tro, för att det skulle vara av nåd, så att löftet kunde bliva beståndande för all hans säd, icke blott för dem som hörde till lagens folk, utan ock för dem som allenast hade Abrahams tro.
Han är ju allas vår fader,
enligt detta skriftens ord: »Jag har bestämt dig till att bliva en fader till många folk»; han är detta inför den Gud som han trodde, inför honom som gör de döda levande och kallar på de ting som icke äro till, likasom voro de till.
Och där ingen förhoppning fanns, där hoppades han ändå och trodde; och han kunde så bliva »en fader till många folk», efter vad som var förutsagt: »Så skall din säd bliva.»
Och han försvagades icke i sin tro, när han betänkte huru hans egen kropp var såsom död -- han var ju omkring hundra år gammal -- och huru jämväl Saras moderliv var såsom dött.
Han tvivlade icke på Guds löfte i otro, utan blev fastmer starkare i sin tro; ty han ärade Gud
och var fullt viss om att vad Gud hade lovat, det var han också mäktig att hålla.
Därför räknades det honom ock till rättfärdighet.
Men att det så tillräknades honom, det är skrivet icke såsom gällde det allenast honom,
utan det skulle gälla också oss; ty det skall tillräknas jämväl oss, oss som tro på honom som från de döda uppväckte Jesus, vår Herre,
vilken utgavs för våra synders skull och uppväcktes för vår rättfärdiggörelses skull.
Då vi nu hava blivit rättfärdiggjorda av tro, hava vi frid med Gud genom vår Herre Jesus Kristus
-- genom vilken vi ock hava fått tillträde till den nåd vari vi nu stå -- och vi berömma oss i hoppet om Guds härlighet.
Och icke det allenast, vi till och med berömma oss av våra lidanden, eftersom vi veta att lidandet verkar ståndaktighet,
och ståndaktigheten beprövad fasthet, och fastheten hopp,
och hoppet låter oss icke komma på skam; ty Guds kärlek är utgjuten i våra hjärtan genom den helige Ande, vilken har blivit oss given.
Ty medan vi ännu voro svaga, led Kristus, när tiden var inne, döden för oss ogudaktiga.
Näppeligen vill ju eljest någon dö ens för en rättfärdig man -- om nu ock till äventyrs någon kan hava mod att dö för den som har gjort honom gott --
men Gud bevisar sin kärlek till oss däri att Kristus dog för oss, medan vi ännu voro syndare.
Så mycket mer skola vi därför, sedan vi nu hava blivit rättfärdiggjorda i och genom hans blod, också genom honom bliva frälsta undan vredesdomen.
Ty om vi, medan vi voro Guds ovänner, blevo försonade med honom genom hans Sons död, så skola vi, sedan vi hava blivit försonade, ännu mycket mer bliva frälsta i och genom hans liv.
Och icke det allenast; vi berömma oss ock av Gud genom vår Herre Jesus Kristus, genom vilken vi nu hava undfått försoningen.
Därför är det så: Genom en enda människa har synden kommit in i världen och genom synden döden; och så har döden kommit över alla människor, eftersom de alla hava syndat.
Ty synd fanns i världen redan innan lagen fanns.
Men synd tillräknas icke där ingen lag finnes;
och dock har under tiden från Adam till Moses döden haft väldet också över dem som icke hade syndat genom en överträdelse, i likhet med vad Adam gjorde, han som är en förebild till den som skulle komma.
Likväl är det icke så med nådegåvan, som det var med syndafallet.
Ty om genom en endas fall de många hava blivit döden underlagda, så har ännu mycket mer Guds nåd och gåvan i och genom nåd -- vilken, också den, är kommen genom en enda människa, Jesus Kristus -- blivit på ett överflödande sätt de många beskärd.
Och med gåvan är det icke såsom det var med det som kom genom denne ene som syndade: domen kom genom en enda, och ledde till en fördömelsedom, men nådegåvan kom i följd av mångas fall, och ledde till en rättfärdiggörelsedom.
Och om döden på grund av en endas fall kom till konungavälde genom denne ene, så skola ännu mycket mer de som undfå den överflödande nåden och rättfärdighetsgåvan få konungsligt välde i liv, också det genom en enda, Jesus Kristus. --
Alltså, likasom det, som kom genom en endas fall, för alla människor ledde till en fördömelsedom, så leder det, som kom genom rättfärdiggörelsedomen förmedelst en enda, för alla människor till en rättfärdiggörelse som medför liv.
Ty såsom genom en enda människas olydnad de många fingo stå såsom syndare, så skola ock genom en endas lydnad de många stå såsom rättfärdiga.
Men lagen har därjämte kommit in, för att fallet skulle bliva så mycket större; dock, där synden blev större, där överflödade nåden mycket mer.
Ty såsom synden hade utövat sitt välde i och genom döden, så skulle nu ock nåden genom rättfärdighet utöva sitt välde till evigt liv, och det genom Jesus Kristus, vår Herre.
Vad skola vi då säga?
Skola vi förbliva i synden, för att nåden skall bliva så mycket större?
Bort det!
Vi som hava dött från synden, huru skulle vi ännu kunna leva i den?
Veten I då icke att vi alla som hava blivit döpta till Kristus Jesus, vi hava blivit döpta till hans död?
Och vi hava så, genom detta dop till döden, blivit begravna med honom, för att, såsom Kristus uppväcktes från de döda genom Faderns härlighet, också vi skola vandra i ett nytt väsende, i liv.
Ty om vi hava vuxit samman med honom genom en lika död, så skola vi ock vara sammanvuxna med honom genom en lika uppståndelse.
Vi veta ju detta, att vår gamla människa har blivit korsfäst med honom, för att syndakroppen skall göras om intet, så att vi icke mer tjäna synden.
Ty den som är död, han är friad ifrån synden.
Hava vi nu dött med Kristus, så tro vi att vi ock skola leva med honom,
eftersom vi veta att Kristus, sedan han har uppstått från de döda, icke mer dör; döden råder icke mer över honom.
Ty hans död var en död från synden en gång för alla, men hans liv är ett liv för Gud.
Så mån ock I hålla före att I ären döda från synden och leven för Gud, i Kristus Jesus.
Låten därför icke synden hava väldet i edra dödliga kroppar, så att I lyden deras begärelser.
Och ställen icke edra lemmar i syndens tjänst, att vara orättfärdighetsvapen, utan ställen eder själva i Guds tjänst, såsom de där från döden hava kommit till livet, och edra lemmar i Guds tjänst, att vara rättfärdighetsvapen.
Ty synden skall icke råda över eder, eftersom I icke stån under lagen, utan under nåden.
Huru är det alltså?
Skola vi synda, eftersom vi icke stå under lagen, utan under nåden?
Bort det!
I veten ju, att när I ställen eder i någons tjänst för att lyda honom, så ären I tjänare under denne, som I sålunda lyden, vare sig det är under synden, vilket leder till död, eller under lydnaden, vilket leder till rättfärdighet.
Men Gud vare tack för att den tid är förbi, då I voren syndens tjänare, och för att I haven blivit av hjärtat lydiga, så att I följen den lära som har givits eder till mönsterbild,
och för att I, när I nu haven gjorts fria ifrån synden, haven blivit tjänare under rättfärdigheten --
om jag nu får tala på människosätt, för eder köttsliga svaghets skull.
Ja, likasom I förr ställden edra lemmar i orenhetens och orättfärdighetens tjänst, till orättfärdighet, så mån I nu ställa edra lemmar i rättfärdighetens tjänst, till helgelse.
Medan I voren syndens tjänare, voren I ju fria ifrån rättfärdighetens tjänst;
men vilken frukt skördaden I då därav?
Jo, det som I nu blygens för; änden på sådant är ju döden.
Men nu, då I haven gjorts fria ifrån synden och blivit Guds tjänare, nu skörden I frukten av detta: I varden helgade; och änden bliver att I undfån evigt liv.
Ty den lön som synden giver är döden, men den gåva som Gud av nåd giver är evigt liv, i Kristus Jesus, vår Herre.
Eller veten I icke, mina bröder -- jag talar ju till sådana som känna lagen -- att lagen råder över en människa för så lång tid som hon lever?
Så är ju en gift kvinna genom lag bunden vid sin man, så länge denne lever; men om mannen dör, då är hon löst från den lag som band henne vid mannen.
Alltså, om hon giver sig åt en annan man, medan hennes man lever, så kallas hon äktenskapsbryterska; men om mannen dör, då är hon fri ifrån lagen, så att hon icke är äktenskapsbryterska, om hon giver sig åt en annan man.
Så haven ock I, mina bröder, genom Kristi kropp blivit dödade från lagen för att tillhöra en annan, nämligen honom som har uppstått från de döda, på det att vi må bära frukt åt Gud.
Ty medan vi ännu voro i ett köttsligt väsende, voro de syndiga lustar, som uppväcktes genom lagen, verksamma i våra lemmar till att bära frukt åt döden.
Men nu äro vi lösta från lagen, i det att vi hava dött från det varunder vi förr höllos fångna; och så tjäna vi nu i Andens nya väsende, och icke i bokstavens gamla väsende.
Vad skola vi då säga?
Är lagen synd?
Bort det!
Men synden skulle jag icke hava lärt känna, om icke genom lagen; ty jag hade icke vetat av begärelsen, om icke lagen hade sagt: »Du skall icke hava begärelse.»
Men då nu synden fick tillfälle, uppväckte den genom budordet allt slags begärelse i mig.
Ty utan lag är synden död.
Jag levde en gång utan lag; men när budordet kom, fick synden liv,
och jag hemföll åt döden.
Så befanns det att budordet, som var givet till liv, det blev mig till död;
ty då synden fick tillfälle, förledde den mig genom budordet och dödade mig genom det.
Alltså är visserligen lagen helig, och budordet heligt och rättfärdigt och gott.
Har då verkligen det som är gott blivit mig till död?
Bort det!
Men synden har blivit det, för att så skulle varda uppenbart att den var synd, i det att den genom något som självt var gott drog över mig död; och så skulle synden bliva till övermått syndig, genom budordet.
Vi veta ju att lagen är andlig, men jag är av köttslig natur, såld till träl under synden.
Ty jag kan icke fatta att jag handlar såsom jag gör; jag gör ju icke vad jag vill, men vad jag hatar, det gör jag.
Om jag nu gör det som jag icke vill, så giver jag mitt bifall åt lagen och vidgår att den är god.
Så är det nu icke mer jag som gör sådant, utan synden, som bor i mig.
Ty jag vet att i mig, det är i mitt kött, bor icke något gott; viljan är väl tillstädes hos mig, men att göra det goda förmår jag icke.
Ja, det goda som jag vill gör jag icke; men det onda som jag icke vill, det gör jag.
Om jag alltså gör vad jag icke vill, så är det icke mer jag som gör det, utan synden, som bor i mig.
Så finner jag nu hos mig, som har viljan att göra det goda, den lagen, att det onda fastmer är tillstädes hos mig.
Ty efter min invärtes människa har jag min lust i Guds lag;
men i mina lemmar ser jag en annan lag, en som ligger i strid med den lag som är i min håg, en som gör mig till fånge under syndens lag, som är i mina lemmar.
Jag arma människa!
Vem skall frälsa mig från denna dödens kropp? --
Gud vare tack, genom Jesus Kristus, vår Herre!
Alltså tjänar jag, sådan jag är i mig själv, visserligen med min håg Guds lag, men med köttet tjänar jag syndens lag.
Så finnes nu ingen fördömelse för dem som äro i Kristus Jesus.
Ty livets Andes lag har i Kristus Jesus gjort mig fri ifrån syndens och dödens lag.
Ty det som lagen icke kunde åstadkomma, i det den var försvagad genom köttet, det gjorde Gud, då han, för att borttaga synden, sände sin Son i syndigt kötts gestalt och fördömde synden i köttet.
Så skulle lagens krav uppfyllas i oss, som vandra icke efter köttet, utan efter Anden.
Ty de som äro köttsliga, de hava sitt sinne vänt till vad köttet tillhör; men de som äro andliga, de hava sitt sinne vänt till vad Anden tillhör.
Och köttets sinne är död, medan Andens sinne är liv och frid.
Köttets sinne är nämligen fiendskap mot Gud, eftersom det icke är Guds lag underdånigt, ej heller kan vara det.
Men de som äro i ett köttsligt väsende kunna icke behaga Gud.
I åter ären icke i ett köttsligt väsende, utan i ett andligt, om eljest Guds Ande bor i eder; men den som icke har Kristi Ande, han hör icke honom till.
Om nu Kristus är i eder, så är väl kroppen hemfallen åt döden, för syndens skull, men Anden är liv, för rättfärdighetens skull.
Och om dens Ande, som uppväckte Jesus från de döda, bor i eder, så skall han som uppväckte Kristus Jesus från de döda göra också edra dödliga kroppar levande, genom sin Ande, som bor i eder.
Alltså, mina bröder, hava vi icke någon förpliktelse mot köttet, så att vi skola leva efter köttet.
Ty om i leven efter köttet, så skolen I dö; men om I genom ande döden kroppens gärningar, så skolen I leva.
Ty alla de som drivas av Guds Ande, de äro Guds barn.
I haven ju icke fått en träldomens ande, så att I åter skullen känna fruktan; I haven fått en barnaskapets ande, i vilken vi ropa: »Abba!
Fader!»
Anden själv vittnar med vår ande att vi äro Guds barn.
Men äro vi barn, så äro vi ock arvingar, nämligen Guds arvingar och Kristi medarvingar, om vi eljest lida med honom, för att också med honom bliva förhärligade.
Ty jag håller före att denna tidens lidanden intet betyda, i jämförelse med den härlighet som kommer att uppenbaras på oss.
Ty skapelsens trängtan sträcker sig efter Guds barns uppenbarelse.
Skapelsen har ju blivit lagd under förgängligheten, icke av eget val, utan för dens skull, som lade den därunder; dock så, att en förhoppning skulle finnas,
att också skapelsen en gång skall bliva frigjord ifrån sin träldom under förgängelsen och komma till den frihet som tillhör Guds barns härlighet.
Vi veta ju att ännu i denna stund hela skapelsen samfällt suckar och våndas.
Och icke den allenast; också vi själva, som hava fått Anden såsom förstlingsgåva, också vi sucka inom oss och bida efter barnaskapet, vår kropps förlossning.
Ty i hoppet äro vi frälsta.
Men ett hopp som man ser fullbordat är icke mer ett hopp; huru kan någon hoppas det som han redan ser?
Om vi nu hoppas på det som vi icke se, så bida vi därefter med ståndaktighet.
Så kommer ock Anden vår svaghet till hjälp; ty vad vi rätteligen böra bedja om, det veta vi icke, men Anden själv manar gott för oss med outsägliga suckar.
Och han som rannsakar hjärtan, han vet vad Anden menar, ty det är efter Guds behag som han manar gott för de heliga.
Men vi veta att för dem som älska Gud samverkar allt till det bästa, för dem som äro kallade efter hans rådslut.
Ty dem som förut hava blivit kända av honom, dem har han ock förut bestämt till att bliva hans Sons avbilder, honom lika, så att denne skulle bliva den förstfödde bland många bröder.
Och dem som han har förut bestämt, dem kallar han ock, och dem som han har kallat, dem rättfärdiggör han ock, och dem som han har rättfärdiggjort, dem förhärligar han ock.
Vad skola vi nu säga härom?
Är Gud för oss, vem kan då vara emot oss?
Han som icke har skonat sin egen Son, utan utgivit honom för oss alla, huru skulle han kunna annat än också skänka oss allt med honom?
Vem vill anklaga Guds utvalda?
Gud är den som rättfärdiggör.
Vem är den som vill fördöma?
Kristus Jesus är den som har dött, ja, än mer, den som har uppstått; och han sitter på Guds högra sida, han manar ock gott för oss.
Vem skulle kunna skilja oss från Kristi kärlek?
Månne bedrövelse eller ångest eller förföljelse eller hunger eller nakenhet eller fara eller svärd?
Så är ju skrivet: »För din skull varda vi dödade hela dagen; vi hava blivit aktade såsom slaktfår.»
Nej, i allt detta vinna vi en härlig seger genom honom som har älskat oss.
Ty jag är viss om att varken död eller liv, varken änglar eller andefurstar, varken något som nu är eller något som skall komma,
varken någon makt i höjden eller någon makt i djupet, ej heller något annat skapat skall kunna skilja oss från Guds kärlek i Kristus Jesus, vår Herre.
Jag talar sanning i Kristus, jag ljuger icke -- därom bär mitt samvete mig vittnesbörd i den helige Ande --
när jag säger att jag har stor bedrövelse och oavlåtligt kval i mitt hjärta.
Ja, jag skulle önska att jag själv vore förbannad och bortkastad från Kristus, om detta kunde gagna mina bröder, mina fränder efter köttet.
De äro ju israeliter, dem tillhöra barnaskapet och härligheten och förbunden och lagstiftningen och tempeltjänsten och löftena.
Dem tillhöra ock fäderna, och från dem är Kristus kommen efter köttet, han som är över allting, Gud, högtlovad i evighet, amen.
Detta säger jag icke som om Guds löftesord skulle hava blivit om intet.
Ty »Israel», det är icke detsamma som alla de som härstamma från Israel.
Ej heller äro de alla »barn», därför att de äro Abrahams säd.
Nej, det heter: »Genom Isak är det som säd skall uppkallas efter dig.»
Detta vill säga: Icke de äro Guds barn, som äro barn efter köttet, men de som äro barn efter löftet, de räknas för säd.
Ty ett löftesord var det ordet: »Vid denna tid skall jag komma tillbaka, och då skall Sara hava en son.»
Än mer: så skedde ock, när Rebecka genom en och samme man, nämligen vår fader Isak, blev moder till sina barn.
Ty förrän dessa voro födda, och innan de ännu hade gjort vare sig gott eller ont, blev det ordet henne sagt -- för att Guds utkorelse-rådslut skulle bliva beståndande, varvid det icke skulle bero på någons gärningar, utan på honom som kallar --
det ordet: »Den äldre skall tjäna den yngre.»
Så är ock skrivet: »Jakob älskade jag, men Esau hatade jag.»
Vad skola vi då säga?
Kan väl orättfärdighet finnas hos Gud?
Bort det!
Han säger ju till Moses: »Jag skall vara barmhärtig mot den jag vill vara barmhärtig emot, och jag skall förbarma mig över den jag vill förbarma mig över.»
Alltså beror det icke på någon människas vilja eller strävan, utan på Guds barmhärtighet.
Ty skriften säger till Farao: »Just därtill har jag låtit dig uppstå, att jag skall visa min makt på dig, och att mitt namn skall varda förkunnat på hela jorden.»
Alltså är han barmhärtig mot vem han vill, och vem han vill förhärdar han.
Nu torde du säga till mig: »Vad har han då att förebrå oss?
Kan väl någon stå emot hans vilja?»
O människa, vem är då du, som vill träta med Gud?
Icke skall verket säga till sin mästare: »Varför gjorde du mig så?»
Har icke krukmakaren den makten över leret, att han av samma lerklump kan göra ett kärl till hedersamt bruk, ett annat till mindre hedersamt?
Men om nu Gud, när han ville visa sin vrede och uppenbara sin makt, likväl i stor långmodighet hade fördrag med »vredens kärl», som voro färdiga till fördärv, vad har du då att säga?
Och om han gjorde detta för att tillika få uppenbara sin härlighets rikedom på »barmhärtighetens kärl», som han förut hade berett till härlighet?
Och till att vara sådana har han ock kallat oss, icke allenast dem som äro av judisk börd, utan jämväl dem som äro av hednisk.
Så säger han ock hos Oseas: »Det folk som icke var mitt folk, det skall jag kalla 'mitt folk', och henne som jag icke älskade skall jag kalla 'min älskade'.
Och det skall ske att på den ort där det sades till dem: 'I ären icke mitt folk', där skola de kallas 'den levande Gudens barn'.»
Men Esaias utropar om Israel: »Om än Israels barn vore till antalet såsom sanden i havet, så skall dock allenast en kvarleva bliva frälst.
Ty dom skall Herren hålla på jorden, en slutdom, som avgör saken med hast.»
Och det är såsom redan Esaias har sagt: »Om Herren Sebaot icke hade lämnat en avkomma kvar åt oss, då vore vi såsom Sodom, vi vore Gomorra lika.»
Vad skola vi då säga?
Jo, att hedningarna, som icke foro efter rättfärdighet, hava vunnit rättfärdighet, nämligen den rättfärdighet som kommer av tro,
under det att Israel, som for efter en rättfärdighetslag, icke har kommit till någon sådan lag.
Varför?
Därför att de icke sökte den på trons väg, utan såsom något som skulle vinnas på gärningarnas väg.
De stötte sig mot stötestenen,
såsom det är skrivet: »Se, jag lägger i Sion en stötesten och en klippa som skall bliva dem till fall; men den som tror på den skall icke komma på skam.»
Mina bröder, mitt hjärtas åstundan och min bön till Gud för dem är att de må bliva frälsta.
Ty det vittnesbördet giver jag dem, att de nitälska för Gud.
Dock göra de detta icke med rätt insikt.
De förstå nämligen icke rättfärdigheten från Gud, utan söka att komma åstad en sin egen rättfärdighet och hava icke givit sig under rättfärdigheten från Gud.
Ty lagen har fått sin ände i Kristus, till rättfärdighet för var och en som tror.
Moses skriver ju om den rättfärdighet som kommer av lagen, att den människa som övar sådan rättfärdighet skall leva genom den.
Men den rättfärdighet som kommer av tro säger så: »Du behöver icke fråga i ditt hjärta: 'Vem vill fara upp till himmelen (nämligen för att hämta Kristus ned)?'
ej heller: 'Vem vill fara ned till avgrunden (nämligen för att hämta Kristus upp ifrån de döda?'»
Vad säger den då? »Ordet är dig nära, i din mun och i ditt hjärta (nämligen ordet om tron, det som vi predika).»
Ty om du med din mun bekänner Jesus vara Herre och i ditt hjärta tror att Gud har uppväckt honom från de döda, då bliver du frälst.
Ty genom hjärtats tro bliver man rättfärdig, och genom munnens bekännelse bliver man frälst.
Skriften säger ju: »Ingen som tror på honom skall komma på skam.»
Det är ingen åtskillnad mellan jude och grek; alla hava ju en och samme Herre, och han har rikedomar att giva åt alla som åkalla honom.
Ty »var och en som åkallar Herrens namn, han skall varda frälst».
Men huru skulle de kunna åkalla den som de icke hava kommit till tro på?
Och huru skulle de kunna tro den som de icke hava hört?
Och huru skulle de kunna höra, om ingen predikade?
Och huru skulle predikare kunna komma, om de icke bleve sända?
Så är och skrivet: »Huru ljuvliga äro icke fotstegen av de män som frambära gott budskap!»
Dock, icke alla hava blivit evangelium lydiga.
Esaias säger ju: »Herre, vem trodde vad som predikades för oss?»
Alltså kommer tron av predikan, men predikan i kraft av Kristi ord.
Jag frågar då: Hava de kanhända icke hört predikas?
Jo, visserligen; det heter ju: »Deras tal har gått ut över hela jorden, och deras ord till världens ändar.»
Jag frågar då vidare: Har Israel kanhända icke förstått det?
Redan Moses säger: »Jag skall uppväcka eder avund mot ett folk som icke är ett folk; mot ett hednafolk utan förstånd skall jag reta eder till vrede.»
Och Esaias går så långt, att han säger: »Jag har låtit mig finnas av dem som icke sökte mig, jag har låtit mig bliva uppenbar för dem som icke frågade efter mig.»
Men om Israel säger han: »Hela dagen har jag uträckt mina händer till ett ohörsamt och gensträvigt folk.»
Så frågar jag nu: Har då Gud förskjutit sitt folk?
Bort det!
Jag är ju själv en israelit, av Abrahams säd och av Benjamins stam.
Gud har icke förskjutit sitt folk, som redan förut hade blivit känt av honom.
Eller veten I icke vad skriften säger, där den talar om Elias, huru denne inför Gud träder upp mot Israel med dessa ord:
»Herre, de hava dräpt dina profeter och rivit ned dina altaren; jag allena är kvar, och de stå efter mitt liv»?
Och vad får han då för svar av Gud? »Jag har låtit bliva kvar åt mig sju tusen män, som icke hava böjt knä för Baal.»
Likaså finnes ock, i den tid som nu är, en kvarleva, i kraft av en utkorelse som har skett av nåd.
Men har den skett av nåd, så har den icke skett på grund av gärningar; annars vore nåd icke mer nåd.
Huru är det alltså?
Vad Israel står efter, det har det icke fått; allenast de utvalda hava fått det, medan de andra hava blivit förstockade.
Så är ju skrivet: »Gud har givit dem en sömnaktighetens ande, ögon som de icke kunna se med och öron som de icke kunna höra med; så är det ännu i dag.»
Och David säger: »Må deras bord bliva dem till en snara, så att de bliva fångade; må det bliva dem till ett giller, så att de få sin vedergällning.
Må deras ögon förmörkas, så att de icke se; böj deras rygg alltid.»
Så frågar jag nu: Var det då för att de skulle komma på fall som de stapplade?
Bort det!
Men genom deras fall har frälsningen kommit till hedningarna, för att de själva skola »uppväckas till avund».
Och har nu redan deras fall varit till rikedom för världen, och har deras fåtalighet varit till rikedom för hedningarna, huru mycket mer skall icke deras fulltalighet så bliva!
Men till eder, I som ären av hednisk börd, säger jag: Eftersom jag nu är en hedningarnas apostel, håller jag mitt ämbete högt --
om jag till äventyrs så skulle kunna »uppväcka avund» hos dem som äro mitt kött och blod och frälsa några bland dem.
Ty om redan deras förkastelse hade med sig världens försoning, vad skall då deras upptagande hava med sig, om icke liv från de döda?
Om förstlingsbrödet är heligt, så är ock hela degen helig; och om roten är helig, så äro ock grenarna heliga.
Men om nu några av grenarna hava brutits bort, och du, som är av ett vilt olivträd, har blivit inympad bland grenarna och med dem har fått delaktighet i det äkta olivträdets saftrika rot,
så må du icke därför förhäva dig över grenarna.
Nej, om du skulle vilja förhäva dig, så besinna att det icke är du som bär roten, utan att roten bär dig.
Nu säger du kanhända: »Det var för att jag skulle bliva inympad som en del grenar brötos bort.»
Visserligen.
För sin otros skull blevo de bortbrutna, och du får vara kvar genom din tro.
Hav då inga högmodiga tankar, utan lev i fruktan.
Ty har Gud icke skonat de naturliga grenarna, så skall han icke heller skona dig.
Se alltså här Guds godhet och stränghet: Guds stränghet mot dem som föllo och hans godhet mot dig, om du nämligen håller dig fast vid hans godhet; annars bliver också du borthuggen.
Men jämväl de andra skola bliva inympade, om de icke hålla fast vid sin otro; Gud är ju mäktig att åter inympa dem.
Ty om du har blivit borthuggen från ditt av naturen vilda olivträd och mot naturen inympats i ett ädelt olivträd, huru mycket snarare skola då icke dessa kunna inympas i sitt eget äkta olivträd, det som de efter naturen tillhöra!
Ty för att I, mina bröder, icke skolen hålla eder själva för kloka, vill jag yppa för eder denna hemlighet: Förstockelse har drabbat en del av Israel och skall fortfara intill dess hedningarna i fulltalig skara hava kommit in;
och så skall hela Israel bliva frälst, såsom det är skrivet: »Från Sion skall förlossaren komma, han skall skaffa bort all ogudaktighet från Jakob.
Och när jag borttager deras synder, då skall detta vara det förbund, som jag gör med dem.»
Se vi nu på evangelium, så äro de hans ovänner, för eder skull; men se vi på utkorelsen, så äro de hans älskade, för fädernas skull.
Ty sina nådegåvor och sin kallelse kan Gud icke ångra.
Såsom I förut voren ohörsamma mot Gud, men nu genom dessas ohörsamhet haven fått barmhärtighet,
så hava nu ock dessa varit ohörsamma, för att de, genom den barmhärtighet som har vederfarits eder, också själva skola få barmhärtighet.
Ty Gud har givit dem alla till pris åt ohörsamhet, för att sedan förbarma sig över dem alla.
O, vilket djup av rikedom och vishet och kunskap hos Gud!
Huru outgrundliga äro icke hans domar, och huru outrannsakliga hans vägar!
Ty »vem har lärt känna Herrens sinne, eller vem har varit hans rådgivare?
Eller vem har först givit honom något, som han alltså bör betala igen?»
Av honom och genom honom och till honom är ju allting.
Honom tillhör äran i evighet, amen.
Så förmanar jag nu eder, mina bröder, vid Guds barmhärtighet, att frambära edra kroppar till ett levande, heligt och Gud välbehagligt offer -- eder andliga tempeltjänst.
Och skicken eder icke efter denna tidsålders väsende, utan förvandlen eder genom edert sinnes förnyelse, så att I kunnen pröva vad som är Guds vilja, vad som är gott och välbehagligt och fullkomligt.
Ty i kraft av den nåd som har blivit mig given, tillsäger jag var och en av eder att icke hava högre tankar om sig än tillbörligt är, utan tänka blygsamt, i överensstämmelse med det mått av tro som Gud har tilldelat var och en.
Ty såsom vi i en och samma kropp hava många lemmar, men alla lemmarna icke hava samma förrättning,
så utgöra ock vi, fastän många, en enda kropp i Kristus, men var för sig äro vi lemmar, varandra till tjänst.
Och vi hava olika gåvor, alltefter den nåd som har blivit oss given.
Har någon profetians gåva, så bruke han den efter måttet av sin tro;
har någon fått en tjänst, så akte han på tjänsten; är någon satt till lärare, så akte han på sitt lärarkall;
är någon satt till att förmana, så akte han på sin plikt att förmana.
Den som delar ut gåvor, han göre det med gott hjärta; den som är satt till föreståndare, han vare det med nit; den som övar barmhärtighet, han göre det med glädje.
Eder kärlek vare utan skrymtan; avskyn det onda, hållen fast vid det goda.
Älsken varandra av hjärtat i broderlig kärlek; söken överträffa varandra i inbördes hedersbevisning.
Varen icke tröga, där det gäller nit; varen brinnande i anden, tjänen Herren.
Varen glada i hoppet, tåliga i bedrövelsen, uthålliga i bönen.
Tagen del i de heligas behov.
Varen angelägna om att bevisa gästvänlighet.
Välsignen dem som förfölja eder; välsignen, och förbannen icke.
Glädjens med dem som äro glada, gråten med dem som gråta.
Varen ens till sinnes med varandra.
Haven icke edert sinne vänt till vad högt är, utan hållen eder till det som är ringa.
Hållen icke eder själva för kloka.
Vedergällen ingen med ont för ont.
Vinnläggen eder om vad gott är inför var man.
Hållen frid med alla människor, om möjligt är, och så mycket som på eder beror.
Hämnens icke eder själva, mina älskade, utan lämnen rum för vredesdomen; ty det är skrivet: »Min är hämnden, jag skall vedergälla det, säger Herren.»
Fastmer, »om din ovän är hungrig, så giv honom att äta, om han är törstig, så giv honom att dricka; ty om du så gör, samlar du glödande kol på hans huvud.»
Låt dig icke övervinnas av det onda, utan övervinn det onda med det goda.
Var och en vare underdånig den överhet som han har över sig.
Ty ingen överhet finnes, som icke är av Gud; all överhet som finnes är förordnad av Gud.
Därför, den som sätter sig upp mot överheten, han står emot vad Gud har förordnat; men de som stå emot detta, de skola få sin dom.
Ty de som hava väldet äro till skräck, icke för dem som göra vad gott är, utan för dem som göra vad ont är.
Vill du vara utan fruktan för överheten, så gör vad gott är; du skall då bliva prisad av den,
ty överheten är en Guds tjänare, dig till fromma.
Men gör du vad ont är, då må du frukta; ty överheten bär icke svärdet förgäves, utan är en Guds tjänare, en hämnare, till att utföra vredesdomen över den som gör vad ont är.
Därför måste man vara den underdånig, icke allenast för vredesdomens skull, utan ock för samvetets skull.
Fördenskull betalen I ju ock skatt; ty överheten förrättar Guds tjänst och är just för detta ändamål ständigt verksam.
Så given åt alla vad I ären dem skyldiga; skatt åt den som skatt tillkommer, tull åt den som tull tillkommer, fruktan åt den som fruktan tillkommer, heder åt den som heder tillkommer.
Varen ingen något skyldiga -- utom när det gäller kärlek till varandra; ty den som älskar sin nästa, han har uppfyllt lagen.
De buden: »Du skall icke begå äktenskapsbrott», »Du skall icke dräpa», »Du skall icke stjäla», »Du skall icke hava begärelse» och vilka andra bud som helst, de sammanfattas ju alla i det ordet: »Du skall älska din nästa såsom dig själv.»
Kärleken gör intet ont mot nästan; alltså är kärleken lagens uppfyllelse.
Akten på allt detta, så mycket mer som I veten vad tiden lider, att stunden nu är inne för eder att vakna upp ur sömnen.
Ty frälsningen är oss nu närmare, än då vi kommo till tro.
Natten är framskriden, och dagen är nära.
Låtom oss därför avlägga mörkrets gärningar och ikläda oss ljusets vapenrustning.
Låtom oss föra en hövisk vandel, såsom om dagen, icke med vilt leverne och dryckenskap, icke i otukt och lösaktighet, icke i kiv och avund.
Ikläden eder fastmer Herren Jesus Kristus, och haven icke sådan omsorg om köttet, att onda begärelser därav uppväckas.
Om någon är svag i tron, så upptagen honom dock vänligt, utan att döma över andras betänkligheter.
Den ene har tro till att äta vad som helst, under det att den som är svag allenast äter vad som växer på jorden.
Den som äter må icke förakta den som icke äter.
Ej heller må den som icke äter döma den som äter; ty Gud har upptagit honom,
och vem är du som dömer en annans tjänare?
Om han står eller faller, det kommer allenast hans egen herre vid; men han skall väl bliva stående, ty Herren är mäktig att hålla honom stående.
Den ene gör skillnad mellan dag och dag, den andre håller alla dagar för lika; var och en vare fullt viss i sitt sinne.
Om någon särskilt aktar på någon dag, så gör han detta för Herren, och om någon äter, så gör han detta för Herren; han tackar ju Gud.
Så ock, om någon avhåller sig från att äta, gör han detta för Herren, och han tackar Gud.
Ty ingen av oss lever för sig själv, och ingen dör för sig själv.
Leva vi, så leva vi för Herren; dö vi, så dö vi för Herren.
Evad vi leva eller dö, höra vi alltså Herren till.
Ty därför har Kristus dött och åter blivit levande, att han skall vara herre över både döda och levande.
Men du, varför dömer du din broder?
Och du åter, varför föraktar du din broder?
Vi skola ju alla en gång stå inför Guds domstol.
Ty det är skrivet: »Så sant jag lever, säger Herren, för mig skola alla knän böja sig, och alla tungor skola prisa Gud.»
Alltså skall var och en av oss inför Gud göra räkenskap för sig själv.
Låtom oss därför icke mer döma varandra.
Dömen hellre så, att ingen må för sin broder lägga en stötesten eller något som bliver honom till fall.
Jag vet väl och är i Herren Jesus viss om att intet i sig självt är orent; allenast om någon håller något för orent, så är det för honom orent.
Om nu genom din mat bekymmer vållas din broder, så vandrar du icke mer i kärleken.
Bliv icke genom din mat till fördärv för den som Kristus har lidit döden för.
Låten alltså icke det goda som I haven fått bliva utsatt för smädelse.
Ty Guds rike består icke i mat och dryck, utan i rättfärdighet och frid och glädje i den helige Ande.
Den som häri tjänar Kristus, han är välbehaglig för Gud och håller provet inför människor.
Vi vilja alltså fara efter det som länder till frid och till inbördes uppbyggelse.
Bryt icke för mats skull ned Guds verk.
Väl är allting rent, men om ätandet för någon är en stötesten, så bliver det för den människan till ondo;
du gör väl i att avhålla dig från att äta kött och dricka vin och från annat som för din broder bliver en stötesten.
Den tro du har må du hava för dig själv inför Gud.
Salig är den som icke måste döma sig själv, när det gäller något som han har prövat vara rätt.
Men om någon hyser betänkligheter och likväl äter, då är han dömd, eftersom det icke sker av tro.
Ty allt som icke sker av tro, det är synd.
Vi som äro starka äro pliktiga att bära de svagas skröpligheter och att icke leva oss själva till behag.
Var och en av oss må leva sin nästa till behag, honom till fromma och honom till uppbyggelse.
Kristus levde ju icke sig själv till behag, utan med honom skedde såsom det är skrivet: »Dina smädares smädelser hava fallit över mig.»
Ty allt vad som fordom har blivit skrivet, det är skrivet oss till undervisning, för att vi, genom ståndaktighet och genom den tröst som skrifterna giva, skola bevara vårt hopp.
Och ståndaktighetens och tröstens Gud give eder att vara ens till sinnes med varandra i Kristi Jesu efterföljelse,
så att I endräktigt och med en mun prisen vår Herres, Jesu Kristi, Gud och Fader.
Därför må den ene av eder vänligt upptaga den andre, såsom Kristus, Gud till ära, har upptagit eder.
Vad jag vill säga är detta: För de omskurna har Kristus blivit en tjänare, till ett vittnesbörd om Guds sannfärdighet, för att bekräfta de löften som hade givits åt fäderna;
hedningarna åter hava fått prisa Gud för hans barmhärtighets skull.
Så är ock skrivet: »Fördenskull vill jag prisa dig bland hedningarna och lovsjunga ditt namn.»
Och åter heter det: »Jublen, I hedningar, med hans folk»;
så ock: »Loven Herren, alla hedningar, ja, honom prise alla folk.»
Så säger ock Esaias: »Telningen från Jessais rot skall komma, ja, han som skall stå upp för att råda över hedningarna; på honom skola hedningarna hoppas.»
Men hoppets Gud uppfylle eder med all glädje och frid i tron, så att I haven ett överflödande hopp i den helige Andes kraft.
Jag är väl redan nu viss om att I, mina bröder, av eder själva ären fulla av godhet, uppfyllda med all kunskap, i stånd jämväl att förmana varandra.
Dock har jag, på ett delvis något dristigt sätt, skrivit till eder med ytterligare påminnelser, detta i kraft av den nåd som har blivit mig given av Gud:
att jag nämligen skall förrätta Kristi Jesu tjänst bland hedningarna och vara en prästerlig förvaltare av Guds evangelium, så att hedningarna bliva ett honom välbehagligt offer, helgat i den helige Ande.
Alltså är det i Kristus Jesus som jag har något att berömma mig av i fråga om min tjänst inför Gud.
Ty jag skall icke drista mig att orda om något annat än vad Kristus, för att göra hedningarna lydaktiga, har verkat genom mig, med ord och med gärning,
genom kraften i tecken och under, genom Andens kraft.
Så har jag, från Jerusalem och runt omkring ända till Illyrien, överallt förkunnat evangelium om Kristus.
Och jag har härvid satt min ära i att icke förkunna evangelium, där Kristi namn redan var känt, ty jag ville icke bygga på en annans grundval;
utan så har skett, som skrivet är: »De för vilka intet har varit förkunnat om honom skola få se, och de som intet hava hört skola förstå.»
Det är också härigenom som jag så många gånger har blivit förhindrad att komma till eder.
Men då jag nu icke mer har något att uträtta i dessa trakter och under ganska många år har längtat efter att komma till eder,
vill jag besöka eder, när jag begiver mig till Spanien.
Jag hoppas nämligen att på genomresan få se eder och att därefter av eder bliva utrustad för färden dit, sedan jag först i någon mån har fått min längtan efter eder stillad.
Men nu far jag till Jerusalem med understöd åt de heliga.
Macedonien och Akaja hava nämligen känt sig manade att göra ett sammanskott åt dem bland de heliga i Jerusalem, som leva i fattigdom.
Ja, därtill hava de känt sig manade; de stå också i skuld hos dem.
Ty om hedningarna hava fått del i deras andliga goda, så äro de å sin sida skyldiga att vara dem till tjänst med sitt lekamliga goda. --
När jag så har fullgjort detta och lämnat i deras händer vad som har blivit insamlat, ämnar jag därifrån begiva mig till Spanien och taga vägen genom eder stad.
Och jag vet, att när jag kommer till eder, kommer jag med Kristi välsignelse i fullt mått.
Och nu uppmanar jag eder, mina bröder, vid vår Herre Jesus Kristus och vid vår kärlek i Anden, att bistå mig i min kamp, genom att bedja för mig till Gud,
att jag må bliva frälst undan de ohörsamma i Judeen, och att det understöd som jag för med mig till Jerusalem må bliva väl mottaget av de heliga.
Så skall jag, om Gud vill, med glädje komma till eder och vederkvicka mig tillsammans med eder.
Fridens Gud vare med eder alla.
Amen.
Jag anbefaller åt eder vår syster Febe, som är församlingstjänarinna i Kenkrea.
Så mottagen då henne i Herren, såsom det höves de heliga, och bistån henne i allt vari hon kan behöva eder; ty hon har själv varit ett stöd för många och jämväl för mig.
Hälsen Priska och Akvila, mina medarbetare i Kristus Jesus.
De hava ju vågat sitt liv för mig; och icke allenast jag tackar dem därför, utan också alla hednaförsamlingar.
Hälsen ock den församling som kommer tillhopa i deras hus.
Hälsen Epenetus, min älskade broder, som är förstlingen av dem som i provinsen Asien hava kommit till Kristus.
Hälsen Maria, som har arbetat så mycket för eder.
Hälsen Andronikus och Junias, mina landsmän och medfångar, som hava ett så gott anseende bland apostlarna, och som längre än jag hava varit i Kristus.
Hälsen Ampliatus, min älskade broder i Herren.
Hälsen Urbanus, vår medarbetare i Kristus, och Stakys, min älskade broder.
Hälsen Apelles, den i Kristus beprövade.
Hälsen dem som höra till Aristobulus' hus.
Hälsen Herodion, min landsman.
Hälsen dem av Narcissus' hus, som äro i Herren.
Hälsen Tryfena och Tryfosa, som arbeta i Herren.
Hälsen Persis, den älskade systern, som har så mycket arbetat i Herren.
Hälsen Rufus, den i Herren utvalde, och hans moder, som också för mig har varit en moder.
Hälsen Asynkritus, Flegon, Hermes, Patrobas, Hermas och de bröder som äro tillsammans med dem.
Hälsen Filologus och Julia, Nereus och hans syster och Olympas och alla de heliga som äro tillsammans med dem.
Hälsen varandra med en helig kyss.
Alla Kristi församlingar hälsa eder.
Men jag förmanar eder, mina bröder, att hava akt på dem som vålla tvedräkt och kunna bliva eder till fall, i strid med den lära som I haven inhämtat; dragen eder ifrån dem.
Ty sådana tjäna icke vår Herre Kristus, utan sin egen buk; och genom sina milda ord och sitt fagra tal bedraga de oskyldiga människors hjärtan.
Eder lydnad är ju känd av alla.
Över eder gläder jag mig därför; men jag skulle önska att I voren visa i fråga om det goda, och menlösa i fråga om det onda.
Och fridens Gud skall snart låta Satan bliva krossad under edra fötter.
Vår Herres, Jesu Kristi, nåd vare med eder.
Timoteus, min medarbetare, hälsar eder: så göra ock Lucius och Jason och Sosipater, mina landsmän.
Jag, Tertius, som har nedskrivit detta brev, hälsar eder i Herren.
Gajus, min och hela församlingens värd, hälsar eder.
Erastus, stadens kamrerare, och brodern Kvartus hälsar eder.
284260
Men honom som förmår styrka eder, enligt det evangelium jag förkunnar och min predikan om Jesus Kristus, ja, enligt den nu avslöjade hemlighet som förut under evärdliga tider har varit outtalad,
men som nu har blivit uppenbarad och, enligt den eviga Gudens befallning, blivit, med stöd av profetiska skrifter, kungjord bland alla hedningar, för att bland dem upprätta trons lydnad --
honom, den ende vise Guden, tillhör äran, genom Jesus Kristus, i evigheternas evigheter.
Amen.
Paulus, genom Guds vilja kallad till Kristi Jesu apostel, så ock brodern Sostenes,
hälsar den Guds församling som finnes i Korint, de i Kristus Jesus helgade, dem som äro kallade och heliga, jämte alla andra som åkalla vår Herres, Jesu Kristi, namn, på alla orter där de eller vi bo.
Nåd vare med eder och frid ifrån Gud, vår Fader, och Herren Jesus Kristus.
Jag tackar Gud alltid för eder skull, för den Guds nåd som har blivit eder given i Kristus Jesus,
att I haven i honom blivit rikligen begåvade i alla stycken, i fråga om allt vad tal och kunskap heter.
Så har ju ock vittnesbördet om Kristus blivit befäst hos eder,
så att I icke stån tillbaka i fråga om någon nådegåva, medan I vänten på vår Herres, Jesu Kristi, uppenbarelse.
Han skall ock göra eder ståndaktiga intill änden, så att I ären ostraffliga på vår Herres, Jesu Kristi, dag.
Gud är trofast, han genom vilken I haven blivit kallade till gemenskap med hans Son, Jesus Kristus, vår Herre.
Men jag förmanar eder, mina bröder, vid vår Herres, Jesu Kristi, namn, att alla vara eniga i edert tal och att icke låta söndringar finnas bland eder, utan hålla fast tillhopa i samma sinnelag och samma tänkesätt.
Det har nämligen av Kloes husfolk blivit mig berättat om eder, mina bröder, att tvister hava uppstått bland eder.
Härmed menar jag att bland eder den ene säger: »Jag håller mig till Paulus», den andre: »Jag håller mig till Apollos», en annan: »Jag håller mig till Cefas», åter en annan: »Jag håller mig till Kristus.» --
Är då Kristus delad?
Icke blev väl Paulus korsfäst för eder?
Och icke bleven I väl döpta i Paulus' namn?
Jag tackar Gud för att jag icke har döpt någon bland eder utom Krispus och Gajus,
så att ingen kan säga att I haven blivit döpta i mitt namn.
Dock, jag har döpt också Stefanas' husfolk; om jag eljest har döpt någon vet jag icke.
Ty Kristus har icke sänt mig till att döpa, utan till att förkunna evangelium, och detta icke med en visdom som består i ord, för att Kristi kors icke skall berövas sin kraft.
Ty talet om korset är visserligen en dårskap för dem som gå förlorade, men för oss som bliva frälsta är det en Guds kraft.
Det är ju skrivet: »Jag skall göra de visas vishet om intet, och de förståndigas förstånd skall jag slå ned.»
Ja, var äro de visa?
Var äro de skriftlärda?
Var äro denna tidsålders klyftiga män?
Har icke Gud gjort denna världens visdom till dårskap?
Jo, eftersom världen icke genom sin visdom lärde känna Gud i hans visdom, behagade det Gud att genom den dårskap han lät predikas frälsa dem som tro.
Ty judarna begära tecken, och grekerna åstunda visdom,
vi åter predika en korsfäst Kristus, en som för judarna är en stötesten och för hedningarna en dårskap,
men som för de kallade, vare sig judar eller greker, är en Kristus som är Guds kraft och Guds visdom.
Ty Guds dårskap är visare än människor, och Guds svaghet är starkare än människor.
Ty betänken, mina bröder, huru det var vid eder kallelse: icke många som voro visa efter köttet blevo kallade, icke många mäktiga, icke många av förnämlig släkt.
Men det som för världen var dåraktigt, det utvalde Gud, för att han skulle låta de visa komma på skam.
Och det som i världen var svagt, det utvalde Gud, för att han skulle låta det starka komma på skam.
Och det som i världen var ringa och föraktat, det utvalde Gud -- ja, det som ingenting var -- för att han skulle göra det till intet, som någonting var.
Ty han ville icke att något kött skulle kunna berömma sig inför Gud.
Men hans verk är det, att I ären i Kristus Jesus, som för oss har blivit till visdom från Gud, till rättfärdighet och helgelse och till förlossning,
för att så skall ske, som det är skrivet: »Den som vill berömma sig, han berömme sig av Herren.»
När jag kom till eder, mina bröder, var det också icke med höga ord eller hög visdom som jag kom och frambar för eder Guds vittnesbörd.
Ty jag hade beslutit mig för, att medan jag var bland eder icke veta om något annat än Jesus Kristus, och honom såsom korsfäst.
Och jag uppträdde hos eder i svaghet och med fruktan och mycken bävan.
Och mitt tal och min predikan framställdes icke med övertalande visdomsord, utan med en bevisning i ande och kraft;
ty eder tro skulle icke vara grundad på människors visdom, utan på Guds kraft.
Visdom tala vi dock bland dem som äro fullmogna, men en visdom som icke tillhör denna tidsålder eller denna tidsålders mäktige, vilkas makt bliver till intet.
Nej, vi tala Guds hemliga visdom, den fördolda, om vilken Gud, redan före tidsåldrarnas begynnelse, har bestämt att den skall bliva oss till härlighet,
och som ingen av denna tidsålders mäktige har känt; ty om de hade känt den, så hade de icke korsfäst härlighetens Herre.
Vi tala -- såsom det heter i skriften -- »vad intet öga har sett och intet öra har hört, och vad ingen människas hjärta har kunnat tänka, vad Gud har berett åt dem som älska honom».
Ty för oss har Gud uppenbarat det genom sin Ande.
Anden utrannsakar ju allt, ja ock Guds djuphet.
Ty vilken människa vet vad som är i en människa, utom den människans egen ande?
Likaså känner ingen vad som är i Gud, utom Guds Ande.
Men vi hava icke fått världens ande, utan den Ande som är av Gud, för att vi skola veta vad som har blivit oss skänkt av Gud.
Om detta tala vi ock, icke med sådana ord som mänsklig visdom lär oss, utan med sådana ord som Anden lär oss; vi hava ju att tyda andliga ting för andliga människor.
Men en »själisk» människa tager icke emot vad som hör Guds Ande till.
Det är henne en dårskap, och hon kan icke förstå det, ty det måste utgrundas på ett andligt sätt.
Den andliga människan åter kan utgrunda allt, men själv kan hon icke utgrundas av någon.
Ty »vem har lärt känna Herrens sinne, så att han skulle kunna undervisa honom?»
Men vi hava Kristi sinne.
Och jag kunde icke tala till eder, mina bröder, såsom till andliga människor, utan måste tala såsom till människor av köttslig natur, såsom till dem som ännu äro barn i Kristus.
Mjölk gav jag eder att dricka; fast föda gav jag eder icke, ty det fördrogen I då ännu icke.
Ja, icke ens nu fördragen I det,
eftersom I ännu haven ett köttsligt sinne.
Ty om avund och kiv finnes bland eder, haven I icke då ett köttsligt sinne, och vandren I icke då på vanligt människosätt?
När den ene säger: »Jag håller mig till Paulus» och den andre: »Jag håller mig till Apollos», ären I icke då lika hopen av människor?
Vad är då Apollos?
Vad är Paulus?
Allenast tjänare, genom vilka I haven kommit till tro; och de äro det i mån av vad Herren har beskärt åt var och en av dem.
Jag planterade, Apollos vattnade, men Gud gav växten.
Alltså kommer det icke an på den som planterar, ej heller på den som vattnar, utan på Gud, som giver växten.
Den som planterar och den som vattnar -- den ene är såsom den andre, dock så, att var och en skall få sin särskilda lön efter sitt särskilda arbete.
Ty vi äro Guds medarbetare; I ären ett Guds åkerfält, en Guds byggnad.
Efter den Guds nåd som blev mig given lade jag grunden såsom en förfaren byggmästare, och en annan bygger nu vidare därpå.
Men var och en må se till, huru han bygger därpå.
Ty en annan grund kan ingen lägga, än den som är lagd, nämligen Jesus Kristus;
men om någon bygger på den grunden med guld, silver och dyrbara stenar eller med trä, hö och strå,
så skall det en gång visa sig huru det är med vars och ens verk. »Den dagen» skall göra det kunnigt; ty den skall uppenbaras i eld, och hurudant vars och ens verk är, det skall elden pröva.
Om det byggnadsverk, som någon har uppfört på den grunden, bliver beståndande, så skall han undfå lön;
men om hans verk brännes upp, så skall han gå miste om lönen.
Själv skall han dock bliva frälst, men såsom igenom eld.
Veten I icke att I ären ett Guds tempel och att Guds Ande bor i eder?
Om nu någon fördärvar Guds tempel, så skall Gud fördärva honom; ty Guds tempel är heligt, och det templet ären I.
Ingen bedrage sig själv.
Om någon bland eder menar sig vara vis genom denna tidsålders visdom, så blive han en dåre, för att han skall kunna bliva vis.
Ty denna världens visdom är dårskap inför Gud.
Det är ju skrivet: »Han fångar de visa i deras klokskap»;
så ock: »Herren känner de visas tankar, han vet att de äro fåfängliga.»
Så berömme sig då ingen av människor.
Allt hör ju eder till;
det må vara Paulus eller Apollos eller Cefas eller hela världen, det må vara liv eller död, vad som nu är, eller vad som skall komma, alltsammans hör eder till.
Men I hören Kristus till, och Kristus hör Gud till.
Såsom Kristi tjänare och såsom förvaltare av Guds hemligheter, så må man anse oss.
Vad man nu därutöver söker hos förvaltare är att en sådan må befinnas vara trogen.
För mig betyder det likväl föga att I -- eller överhuvud någon mänsklig domstol -- sätten eder till doms över mig.
Ja, jag vill icke ens sätta mig till doms över mig själv.
Ty väl vet jag intet med mig, men därigenom är jag icke rättfärdigad; det är Herren som sitter till doms över mig.
Dömen därför icke förrän tid är, icke förrän Herren kommer, han som skall draga fram i ljuset vad som är fördolt i mörker och uppenbara alla hjärtans rådslag.
Och då skall var och en undfå av Gud den berömmelse som honom tillkommer.
Detta, mina bröder, har jag nu för eder skull så framställt, som gällde det mig och Apollos; ty jag vill att I skolen i fråga om oss lära eder detta: »Icke utöver vad skrivet är.»
Jag vill icke att I skolen stå emot varandra, uppblåsta var och en över sin lärare.
Vem säger då att du har något företräde?
Och vad äger du, som du icke har fått dig givet?
Men har du nu fått dig givet vad du har, huru kan du då berömma dig, såsom om du icke hade fått det dig givet?
I ären kantänka redan mätta, I haven redan blivit rika; oss förutan haven I blivit sannskyldiga konungar!
Ja, jag skulle önska att I verkligen haden blivit konungar, så att vi kunde få bliva edra medkonungar.
Mig tyckes nämligen att Gud har ställt oss apostlar här såsom de ringaste bland alla, såsom livdömda män; ett skådespel hava vi ju blivit för världen, för både änglar och människor.
Vi äro dårar för Kristi skull, men I ären kloka i Kristus; vi äro svaga, men I ären starka; I ären ärade, men vi äro föraktade.
Ännu i denna stund lida vi både hunger och törst, vi måste gå nakna, vi få uppbära hugg och slag, vi hava intet stadigt hemvist,
vi måste möda oss och arbeta med våra händer.
Vi bliva smädade och välsigna likväl; vi lida förföljelse och härda dock ut;
man talar illa om oss, men vi tala goda ord.
Vi hava blivit såsom världens avskum, såsom var mans avskrap, och vi äro så ännu alltjämt.
Detta skriver jag, icke för att komma eder att blygas, utan såsom en förmaning till mina älskade barn.
Ty om I än haden tio tusen uppfostrare i Kristus, så haven I dock icke många fäder; det var ju jag som i Kristus Jesus genom evangelium födde eder till liv.
Därför förmanar jag eder: Bliven mina efterföljare.
Just för denna saks skull sänder jag nu till eder Timoteus, min älskade och trogne son i Herren; han skall påminna eder om huru jag går till väga i Kristus, i enlighet med den lära jag förkunnar allestädes, i alla församlingar.
Nu är det väl så, att somliga hava blivit uppblåsta, under förmenande att jag icke skulle komma till eder.
Men om Herren så vill, skall jag snart komma till eder; och då skall jag lära känna, icke dessa uppblåsta människors ord, utan deras kraft.
Ty Guds rike består icke i ord, utan i kraft.
Vilketdera viljen I nu: skall jag komma till eder med ris eller i kärlek och saktmods ande?
Det förljudes såväl att överhuvud otukt bedrives bland eder, som ock att sådan otukt förekommer, som man icke ens finner bland hedningarna, nämligen att en son har sin faders hustru.
Och ändå ären I uppblåsta och haven icke fastmer blivit uppfyllda av sådan sorg, att I haven drivit ut ur eder krets den som har gjort detta.
Jag, som väl till kroppen är frånvarande, men till anden närvarande, har för min del redan, såsom vore jag närvarande, fällt domen över den som har förövat en sådan ogärning:
i Herren Jesu namn skola vi komma tillsammans, I och min ande, med vår Herre Jesu kraft,
och överlämna den mannen åt Satan till köttets fördärv, för att anden skall bliva frälst på Herren Jesu dag.
Det är icke väl beställt med eder berömmelse.
Veten I icke att litet surdeg syrar hela degen?
Rensen bort den gamla surdegen, så att I bliven en ny deg.
I ären ju osyrade; ty vi hava ock ett påskalamm, som är slaktat, nämligen Kristus.
Låtom oss därför hålla högtid, icke med gammal surdeg, icke med elakhetens och ondskans surdeg, utan med renhetens och sanningens osyrade bröd.
Jag skrev till eder i mitt brev att I icke skullen hava något umgänge med otuktiga människor --
detta icke sagt i allmänhet, om alla denna världens otuktiga människor eller om giriga och roffare eller om avgudadyrkare; annars måsten I ju rymma ur världen.
Nej, då jag skrev så till eder, menade jag, att om någon som kallades broder vore en otuktig människa eller en girig eller en avgudadyrkare eller en smädare eller en drinkare eller en roffare, så skullen I icke hava något umgänge med en sådan eller äta tillsammans med honom.
Ty icke tillkommer det väl mig att döma dem som äro utanför?
Dem som äro innanför haven I ju att döma;
dem som äro utanför skall Gud döma. »I skolen driva ut ifrån eder den som är ond.»
Huru kan någon av eder taga sig för, att när han har sak med en annan, gå till rätta icke inför de heliga, utan inför de orättfärdiga?
Veten I då icke att de heliga skola döma världen?
Men om nu I skolen sitta till doms över världen, ären I då icke goda nog att döma i helt ringa mål?
I veten ju att vi skola döma änglar; huru mycket mer böra vi icke då kunna döma i timliga ting?
Och likväl, när I nu haven före något mål som gäller sådana ting, sätten I till domare just dem som äro ringa aktade i församlingen!
Eder till blygd säger jag detta.
Är det då så omöjligt att bland eder finna någon vis man, som kan bliva skiljedomare mellan sina bröder?
Måste i stället den ene brodern gå till rätta med den andre, och det inför de otrogna?
Överhuvud är redan det en brist hos eder, att I gån till rätta med varandra.
Varför liden I icke hellre orätt?
Varför låten I icke hellre andra göra eder skada?
I stället gören I nu själva orätt och skada, och detta mot bröder.
Veten I då icke att de orättfärdiga icke skola få Guds rike till arvedel?
Faren icke vilse.
Varken otuktiga människor eller avgudadyrkare eller äktenskapsbrytare, varken de som låta bruka sig till synd mot naturen eller de som själva öva sådan synd,
varken tjuvar eller giriga eller drinkare eller smädare eller roffare skola få Guds rike till arvedel.
Sådana voro ock somliga bland eder, men I haven låtit två eder rena, I haven blivit helgade, I haven blivit rättfärdiggjorda i Herrens, Jesu Kristi, namn och i vår Guds Ande.
»Allt är mig lovligt»; ja, men icke allt är nyttigt. »Allt är mig lovligt»; ja, men jag bör icke låta något få makt över mig.
Maten är för buken och buken för maten, men bådadera skall Gud göra till intet.
Däremot är kroppen icke för otukt, utan för Herren, och Herren för kroppen;
och Gud, som har uppväckt Herren, skall ock genom sin kraft uppväcka oss.
Veten I icke att edra kroppar äro Kristi lemmar?
Skall jag nu taga Kristi lemmar och göra dem till en skökas lemmar?
Bort det!
Veten I då icke att den som håller sig till en sköka, han bliver en kropp med henne?
Det heter ju: »De tu skola varda ett kött.»
Men den som håller sig till Herren, han är en ande med honom.
Flyn otukten.
All annan synd som en människa kan begå är utom kroppen; men den som bedriver otukt, han syndar på sin egen kropp.
Veten I då icke att eder kropp är ett tempel åt den helige Ande, som bor i eder, och som I haven undfått av Gud, och att I icke ären edra egna?
I ären ju köpta, och betalning är given.
Så förhärligen då Gud i eder kropp.
Vad nu angår det I haven skrivit om, så svarar jag detta: En man gör visserligen väl i att icke komma vid någon kvinna;
men för att undgå otuktssynder må var man hava sin egen hustru, och var kvinna sin egen man.
Mannen give sin hustru vad han är henne pliktig, sammalunda ock hustrun sin man.
Hustrun råder icke själv över sin kropp, utan mannen; sammalunda råder ej heller mannen över sin kropp, utan hustrun.
Dragen eder icke undan från varandra, om icke möjligen, med bådas samtycke, till en tid, för att I skolen hava ledighet till bönen.
Kommen sedan åter tillsammans, så att Satan icke frestar eder, då I nu icke kunnen leva återhållsamt.
Detta säger jag likväl såsom en tillstädjelse, icke såsom en befallning.
Jag skulle dock vilja att alla människor vore såsom jag.
Men var och en har fått sin särskilda nådegåva från Gud, den ene så, den andre så.
Till de ogifta åter och till änkorna säger jag att de göra väl, om de förbliva i samma ställning som jag.
Men kunna de icke leva återhållsamt, så må de gifta sig; ty det är bättre att gifta sig än att vara upptänd av begär.
Men dem som äro gifta bjuder jag -- dock icke jag, utan Herren; En hustru må icke skilja sig från sin man
(om hon likväl skulle skilja sig, så förblive hon ogift eller förlike sig åter med mannen), ej heller må en man förskjuta sin hustru.
Till de andra åter säger jag själv, icke Herren: Om någon som hör till bröderna har en hustru som icke är troende, och denna är villig att leva tillsammans med honom, så må han icke förskjuta henne.
Likaså, om en hustru har en man som icke är troende, och denne är villig att leva tillsammans med henne, så må hon icke förskjuta mannen.
Ty den icke troende mannen är helgad i och genom sin hustru, och den icke troende hustrun är helgad i och genom sin man, då han är en broder; annars vore ju edra barn orena, men nu äro de heliga. --
Om däremot den icke troende vill skiljas, så må han få skiljas.
En broder eller syster är i sådana fall intet tvång underkastad, och Gud har kallat oss till att leva i frid.
Ty huru kan du veta, du hustru, om du skall frälsa din man?
Eller du man, huru vet du om du skall frälsa din hustru?
Må allenast var och en vandra den väg fram, som Herren har bestämt åt honom, var och en i den ställning vari Gud har kallat honom.
Den ordningen stadgar jag för alla församlingar.
Har någon blivit kallad såsom omskuren, så göre han sig icke åter lik de oomskurna; har någon blivit kallad såsom oomskuren, så låte han icke omskära sig.
Det kommer icke an på om någon är omskuren eller oomskuren; allt beror på huruvida han håller Guds bud.
Var och en förblive i den kallelse vari han var, när han blev kallad.
Har du blivit kallad såsom träl, så låt detta icke gå dig till sinnes; dock, om du kan bliva fri, så begagna dig hellre därav.
Ty den träl som har blivit kallad till att vara i Herren, han är en Herrens frigivne; sammalunda är ock den frie, som har blivit kallad, en Kristi livegne.
I ären köpta, och betalningen är given; bliven icke människors trälar.
Ja, mina bröder, var och en förblive inför Gud i den ställning vari han har blivit kallad.
Vad vidare angår dem som äro jungfrur, så har jag icke att åberopa någon befallning av Herren, utan giver allenast ett råd, såsom en som genom Herrens barmhärtighet har blivit förtroende värd.
Jag menar alltså, med tanke på den nöd som står för dörren, att den människa gör väl, som förbliver såsom hon är.
Är du bunden vid hustru, så sök icke att bliva lös.
Är du utan hustru, så sök icke att få hustru.
Om du likväl skulle gifta dig, så syndar du icke därmed; ej heller syndar en jungfru, om hon gifter sig.
Dock komma de som så göra att draga över sig lekamliga vedermödor; och jag skulle gärna vilja skona eder.
Men det säger jag, mina bröder: Tiden är kort; därför må härefter de som hava hustrur vara såsom hade de inga,
och de som gråta såsom gräte de icke, och de som glädja sig såsom gladde de sig icke, och de som köpa något såsom finge de icke behålla det,
och de som bruka denna världen såsom gjorde de icke något bruk av den.
Ty den nuvarande världsordningen går mot sitt slut;
och jag skulle gärna vilja att I voren fria ifrån omsorger.
Den man som icke är gift ägnar nämligen sin omsorg åt vad som hör Herren till, huru han skall behaga Herren;
men den gifte mannen ägnar sin omsorg åt vad som hör världen till, huru han skall behaga sin hustru,
och så är hans hjärta delat.
Likaså ägnar den kvinna, som icke längre är gift eller som är jungfru, sin omsorg åt vad som hör Herren till, att hon må vara helig till både kropp och ande; men den gifta kvinnan ägnar sin omsorg åt vad som hör världen till, huru hon skall behaga sin man.
Detta säger jag till eder egen nytta, och icke för att lägga något band på eder, utan för att I skolen föra en hövisk vandel och stadigt förbliva vid Herren.
Men om någon menar sig handla otillbörligt mot sin ogifta dotter därmed att hon får bliva överårig, då må han göra såsom han vill, om det nu måste så vara; han begår därmed ingen synd.
Må hon få gifta sig.
Om däremot någon är fast i sitt sinne och icke bindes av något nödtvång, utan kan följa sin egen vilja, och så i sitt sinne är besluten att låta sin ogifta dotter förbliva såsom hon är, då gör denne väl.
Alltså: den som gifter bort sin dotter, han gör väl; och den som icke gifter bort henne, han gör ännu bättre.
En hustru är bunden så länge hennes man lever; men när hennes man är avsomnad, står det henne fritt att gifta sig med vem hon vill, blott det sker i Herren.
Men lyckligare är hon, om hon förbliver såsom hon är.
Så är min mening, och jag tror att också jag har Guds Ande.
Vad åter angår kött från avgudaoffer, så känna vi nog det talet: »Alla hava vi 'kunskap'.» »Kunskapen» uppblåser, men kärleken uppbygger.
Om någon menar sig hava fått någon »kunskap», så har han ännu icke fått kunskap på sådant sätt som han borde hava.
Men den som älskar Gud, han är känd av honom.
Vad alltså angår ätandet av kött från avgudaoffer, så säger jag detta: Vi veta visserligen att ingen avgud finnes till i världen, och att det icke finnes mer än en enda Gud.
Ty om ock några så kallade gudar skulle finnas, vare sig i himmelen eller på jorden -- och det finnes ju många »gudar» och många »herrar» --
så finnes dock för oss allenast en enda Gud: Fadern, av vilken allt är, och till vilken vi själva äro, och en enda Herre: Jesus Kristus, genom vilken allt är, och genom vilken vi själva äro.
Dock, icke alla hava denna kunskap, utan somliga, som äro vana att ännu alltjämt tänka på avguden, äta köttet såsom avgudaofferskött.
Och eftersom deras samvete är svagt, bliver det härigenom befläckat.
Men maten skall icke avgöra vår ställning till Gud.
Avhålla vi oss från att äta, så bliva vi icke därigenom sämre; äta vi, så bliva vi icke därigenom bättre.
Sen likväl till, att denna eder frihet icke till äventyrs bliver en stötesten för de svaga.
Ty om någon får se dig, som har undfått »kunskap», ligga till bords i ett avgudahus, skall då icke hans samvete, om han är svag, därav »bliva uppbyggt» på det sätt att han äter köttet från avgudaoffer?
Genom din »kunskap» går ju då den svage förlorad -- han, din broder, som Kristus har lidit döden för.
Om I på sådant sätt synden mot bröderna och såren deras svaga samveten, då synden I mot Kristus själv.
Därför, om maten kan bliva min broder till fall, så vill jag sannerligen hellre för alltid avstå från att äta kött, på det att jag icke må bliva min broder till fall.
Är jag icke fri?
Är jag icke en apostel?
Har jag icke sett Jesus, vår Herre?
Ären icke I mitt verk i Herren?
Om jag icke för andra är en apostel, så är jag det åtminstone för eder, ty I själva ären i Herren inseglet på mitt apostlaämbete.
Detta är mitt försvar mot dem som sätta sig till doms över mig.
Skulle vi kanhända icke hava rätt att få mat och dryck?
Skulle vi icke hava rätt att få såsom hustru föra med oss på våra resor någon som är en syster, vi likaväl som de andra apostlarna och Herrens bröder och särskilt Cefas?
Eller äro jag och Barnabas de enda som icke hava rätt att vara fritagna ifrån kroppsarbete?
Vem tjänar någonsin i krig på egen sold?
Vem planterar en vingård och äter icke dess frukt?
Eller vem vaktar en hjord och förtär icke mjölk från hjorden?
Icke talar jag väl detta därför att människor pläga så tala?
Säger icke själva lagen detsamma?
I Moses' lag är ju skrivet: »Du skall icke binda munnen till på oxen som tröskar.»
Månne det är om oxarna som Gud har sådan omsorg?
Eller säger han det icke i alla händelser med tanke på oss?
Jo, för vår skull blev det skrivet, att den som plöjer bör plöja med en förhoppning, och att den som tröskar bör göra det i förhoppning om att få sin del.
Om vi hava sått åt eder ett utsäde av andligt gott, är det då för mycket, om vi få inbärga från eder en skörd av lekamligt gott?
Om andra hava en viss rättighet över eder, skulle då icke vi än mer hava det?
Och likväl hava vi icke gjort bruk av den rättigheten, utan vi fördraga allt, för att icke lägga något hinder i vägen för Kristi evangelium.
I veten ju att de som förrätta tjänsten i helgedomen få sin föda ifrån helgedomen, och att de som äro anställda vid altaret få sin del, när altaret får sin.
Så har ock Herren förordnat att de som förkunna evangelium skola hava sitt uppehälle av evangelium.
Men jag för min del har icke gjort bruk av någon sådan förmån.
Detta skriver jag nu icke, för att jag själv skall få någon sådan; långt hellre ville jag dö.
Nej, ingen skall göra min berömmelse om intet.
Ty om jag förkunnar evangelium, så är detta ingen berömmelse för mig.
Jag måste ju så göra; och ve mig, om jag icke förkunnade evangelium!
Gör jag det av egen drift, så har jag rätt till lön; men då jag nu icke gör det av egen drift, så är den syssla som jag är betrodd med allenast en livegen förvaltares. --
Vilken är alltså min lön?
Jo, just den, att när jag förkunnar evangelium, så gör jag detta utan kostnad för någon, i det att jag avstår från att göra bruk av den rättighet jag har såsom förkunnare av evangelium.
Ty fastän jag är fri och oberoende av alla, har jag dock gjort mig till allas tjänare, för att jag skall vinna dess flera.
För judarna har jag blivit såsom en jude, för att kunna vinna judar; för dom som stå under lagen har jag, som själv icke står under lagen, blivit såsom stode jag under lagen, för att kunna vinna dem som stå under lagen.
För dem som äro utan lag har jag, som icke är utan Guds lag, men är i Kristi lag, blivit såsom vore jag utan lag, för att jag skall vinna dem som äro utan lag.
För de svaga har jag blivit svag, för att kunna vinna de svaga; för alla har jag blivit allt, för att jag i alla händelser skall frälsa några.
Men allt gör jag för evangelii skull, för att också jag skall bliva delaktig av dess goda.
I veten ju, att fastän de som löpa på tävlingsbanan allasammans löpa, så vinner allenast en segerlönen.
Löpen såsom denne, för att I mån vinna lönen.
Men alla som vilja deltaga i en sådan tävlan pålägga sig återhållsamhet i alla stycken: dessa för att vinna en förgänglig segerkrans, men vi för att vinna en oförgänglig.
Jag för min del löper alltså icke såsom gällde det ett ovisst mål; jag kämpar icke likasom en man som hugger i vädret.
Fastmer tuktar jag min kropp och kuvar den, för att jag icke, när jag predikar för andra, själv skall komma till korta vid provet.
Ty jag vill säga eder detta, mina bröder: Våra fäder voro alla under molnskyn och gingo alla genom havet;
alla blevo de i molnskyn och i havet döpta till Moses;
alla åto de samma andliga mat,
och alla drucko de samma andliga dryck -- de drucko nämligen ur en andlig klippa, som åtföljde dem, och den klippan var Kristus.
Men de flesta av dem hade Gud icke behag till; de blevo ju nedgjorda i öknen.
Detta skedde oss till en varnagel, för att vi icke skulle hava begärelse till det onda, såsom de hade begärelse därtill.
Ej heller skolen I bliva avgudadyrkare, såsom somliga av dem blevo; så är ju skrivet: »Folket satte sig ned till att äta och dricka, och därpå stodo de upp till all leka.»
Låtom oss icke heller bedriva otukt, såsom somliga av dem gjorde, varför ock tjugutre tusen föllo på en enda dag.
Låtom oss icke heller fresta Kristus, såsom somliga av dem gjorde, varför de ock blevo dödade av ormarna.
Knorren icke heller, såsom somliga av dem gjorde, varför de ock blevo dödade av »Fördärvaren».
Men detta vederfors dem för att tjäna till en varnagel, och det blev upptecknat till lärdom för oss, som hava tidernas ände inpå oss.
Därför, den som menar sig stå, han må se till, att han icke faller.
Inga andra frestelser hava mött eder än sådana som vanligen möta människor.
Och Gud är trofast; han skall icke tillstädja att I bliven frestade över eder förmåga, utan när han låter frestelsen komma, skall han ock bereda en utväg därur, så att I kunnen härda ut i den.
Alltså, mina älskade, undflyn avgudadyrkan.
Jag säger detta till eder såsom till förståndiga människor; själva mån I döma om det som jag säger.
Välsignelsens kalk, över vilken vi uttala välsignelsen, är icke den en delaktighet av Kristi blod?
Brödet, som vi bryta, är icke det en delaktighet av Kristi kropp?
Eftersom det är ett enda bröd, så äro vi, fastän många, en enda kropp, ty alla få vi vår del av detta ena bröd.
Sen på det lekamliga Israel: äro icke de som äta av offren delaktiga i altaret?
Vad vill jag då säga härmed?
Månne att avgudaofferskött är någonting, eller att en avgud är någonting?
Nej, det vill jag säga, att vad hedningarna offra, det offra de åt onda andar och icke åt Gud; och jag vill icke att I skolen hava någon gemenskap med de onda andarna.
I kunnen icke dricka Herrens kalk och tillika onda andars kalk; I kunnen icke hava del i Herrens bord och tillika i onda andars bord.
Eller vilja vi reta Herren?
Äro då vi starkare än han?
»Allt är lovligt»; ja, men icke allt är nyttigt. »Allt är lovligt»; ja, men icke allt uppbygger.
Ingen söke sitt eget bästa, utan envar den andres.
Allt som säljes i köttboden mån I äta; I behöven icke för samvetets skull göra någon undersökning därom.
Ty »jorden är Herrens, och allt vad därpå är».
Om någon av dem som icke äro troende bjuder eder till sig och I viljen gå till honom, så mån I äta av allt som sättes fram åt eder; I behöven icke för samvetets skull göra någon undersökning därom.
Men om någon då säger till eder: »Detta är offerkött», så skolen I avhålla eder från att äta, för den mans skull, som gav saken till känna, och för samvetets skull --
jag menar icke ditt eget samvete, utan den andres; ty varför skulle jag låta min frihet dömas av en annans samvete?
Om jag äter därav med tacksägelse, varför skulle jag då bliva smädad för det som jag tackar Gud för?
Alltså, vare sig I äten eller dricken, eller vadhelst annat I gören, så gören allt till Guds ära.
Bliven icke för någon till en stötesten, varken för judar eller för greker eller för Guds församling;
varen såsom jag, som i alla stycken fogar mig efter alla och icke söker min egen nytta, utan de mångas, för att de skola bliva frälsta.
Varen I mina efterföljare, såsom jag är Kristi.
Jag prisar eder för det att I i alla stycken haven mig i minne och hållen fast vid mina lärdomar, såsom de äro eder givna av mig.
Men jag vill att I skolen inse detta, att Kristus är envar mans huvud, och att mannen är kvinnans huvud, och att Gud är Kristi huvud.
Var och en man som har sitt huvud betäckt, när han beder eller profeterar, han vanärar sitt huvud.
Men var kvinna som beder eller profeterar med ohöljt huvud, hon vanärar sitt huvud, ty det är då alldeles som om hon hade sitt hår avrakat.
Om en kvinna icke vill hölja sig, så kan hon lika väl låta skära av sitt hår; men eftersom det är en skam för en kvinna att låta skära av sitt hår eller att låta raka av det, så må hon hölja sig.
En man är icke pliktig att hölja sitt huvud, eftersom han är Guds avbild och återspeglar hans härlighet, då kvinnan däremot återspeglar mannens härlighet.
Ty mannen är icke av kvinnan, utan kvinnan av mannen.
Icke heller skapades mannen för kvinnans skull, utan kvinnan för mannens skull.
Därför bör kvinnan på sitt huvud hava en »makt», för änglarnas skull.
Dock är det i Herren så, att varken kvinnan är till utan mannen, eller mannen utan kvinnan.
Ty såsom kvinnan är av mannen, så är ock mannen genom kvinnan; men alltsammans är av Gud. --
Dömen själva: höves det en kvinnan att ohöljd bedja till Gud?
Lär icke själva naturen eder att det länder en man till vanheder, om han har långt hår,
men att det länder en kvinna till ära, om hon har långt hår?
Håret är ju henne givet såsom slöja.
Om nu likväl någon vill vara genstridig, så mån han veta att vi för vår del icke hava en sådan sedvänja, ej heller andra Guds församlingar.
Detta bjuder jag eder nu.
Men vad jag icke kan prisa är att I kommen tillsammans, icke till förbättring, utan till försämring.
Ty först och främst hör jag sägas att vid edra församlingsmöten söndringar yppa sig bland eder.
Och till en del tror jag att så är.
Ty partier måste ju finnas bland eder, för att det skall bliva uppenbart vilka bland eder som hålla provet.
När I alltså kommen tillsammans med varandra, kan ingen Herrens måltid hållas;
ty vid måltiden tager var och en i förväg själv den mat han har medfört, och så får den ene hungra, medan den andre får för mycket.
Haven I då icke edra hem, där I kunnen äta ock dricka?
Eller är det så, att I förakten Guds församling och viljen komma dem att blygas, som intet hava?
Vad skall jag då säga till eder?
Skall jag prisa eder?
Nej, i detta stycke prisar jag eder icke.
Ty jag har från Herren undfått detta, som jag ock har meddelat eder: I den natt då Herren Jesus blev förrådd tog han ett bröd
och tackade Gud och bröt det och sade: »Detta är min lekamen, som varder utgiven för eder.
Gören detta till min åminnelse.»
Sammalunda tog han ock kalken, efter måltiden, och sade: »Denna kalk är det nya förbundet, i mitt blod.
Så ofta I dricken den, så gören detta till min åminnelse.»
Ty så ofta I äten detta bröd och dricken kalken, förkunnen I Herrens död, till dess att han kommer.
Den som nu på ett ovärdigt sätt äter detta bröd eller dricker Herrens kalk, han försyndar sig på Herrens lekamen och blod.
Pröve då människan sig själv, och äte så av brödet och dricke av kalken.
Ty den som äter och dricker, utan att göra åtskillnad mellan Herrens lekamen och annan spis, han äter och dricker en dom över sig.
Därför finnas ock bland eder många som äro svaga och sjuka, och ganska många äro avsomnade.
Om vi ginge till doms med oss själva, så bleve vi icke dömda.
Men då vi nu bliva dömda, så är detta en Herrens tuktan, som drabbar oss, för att vi icke skola bliva fördömda tillika med världen.
Alltså, mina bröder, när I kommen tillsammans för att hålla måltid, så vänten på varandra.
Om någon är hungrig, då må han äta hemma, så att eder sammankomst icke bliver eder till en dom.
Om det övriga skall jag förordna, när jag kommer.
Vad nu angår dem som hava andliga gåvor, så vill jag säga eder, mina bröder, huru med dem förhåller sig.
I veten att I, medan I voren hedningar, läten eder blindvis föras bort till de stumma avgudarna.
Därför vill jag nu förklara för eder, att likasom ingen som talar i Guds Ande säger: »Förbannad vare Jesus», så kan ej heller någon säga: »Jesus är Herre» annat än i den helige Ande.
Nådegåvorna äro mångahanda, men Anden är en och densamme.
Tjänsterna äro mångahanda, men Herren är en och densamme.
Kraftverkningarna äro mångahanda, men Gud är en och densamme, han som verkar allt i alla.
Men de gåvor i vilka Anden uppenbarar sig givas åt var och en så, att de kunna bliva till nytta.
Så gives genom Anden åt den ene att tala visdomens ord, åt en annan att efter samme Ande tala kunskapens ord,
åt en annan gives tro i samme Ande, åt en annan givas helbrägdagörelsens gåvor i samme ene Ande,
åt en annan gives gåvan att utföra kraftgärningar, åt en annan att profetera, åt en annan att skilja mellan andar, åt en annan att tala tungomål på olika sätt, åt en annan att uttyda, när någon talar tungomål.
Men allt detta verkar densamme ene Anden, i det han, alltefter sin vilja, tilldelar åt var och en någon särskild gåva.
Ty likasom kroppen är en och likväl har många lemmar, och likasom kroppens alla lemmar, fastän de äro många, likväl utgöra en enda kropp, likaså är det med Kristus.
Ty i en och samme Ande äro vi alla döpta till att utgöra en och samma kropp, vare sig vi äro judar eller greker, vare sig vi äro trälar eller fria; och alla hava vi fått en och samme Ande utgjuten över oss.
Kroppen utgöres ju icke heller av en enda lem, utan av många.
Om foten ville säga: »Jag är icke hand, därför hör jag icke till kroppen», så skulle den icke dess mindre höra till kroppen.
Och om örat ville säga: »Jag är icke öga, därför hör jag icke till kroppen», så skulle det icke dess mindre höra till kroppen.
Om hela kroppen vore öga, var funnes då hörseln?
Och om den hel och hållen vore öra, var funnes då lukten?
Men nu har Gud insatt lemmarna i kroppen, var och en av dem på det sätt som han har velat.
Om åter allasammans utgjorde en enda lem, var funnes då själva kroppen?
Men nu är det så, att lemmarna äro många, och att kroppen dock är en enda.
Ögat kan icke säga till handen: »Jag behöver dig icke», ej heller huvudet till fötterna: »Jag behöver eder icke.»
Nej, just de kroppens lemmar som tyckas vara svagast äro som mest nödvändiga.
Och de delar av kroppen, som tyckas oss vara mindre hedersamma, dem bekläda vi med så mycket större heder; och dem som vi blygas för, dem skyla vi med så mycket större blygsamhet,
under det att de andra icke behöva något sådant.
Men när Gud sammanfogade kroppen av olika delar och därvid lät den ringare delen få en så mycket större heder,
så skedde detta, för att söndring icke skulle uppstå i kroppen, utan alla lemmar endräktigt hava omsorg om varandra.
Om nu en lem lider, så lida alla de andra lemmarna med den; om åter en lem äras, så glädja sig alla de andra lemmarna med den.
Men nu ären I Kristi kropp och hans lemmar, var och en i sin mån.
Och Gud har i församlingen satt först och främst några till apostlar, för det andra några till profeter, för det tredje några till lärare, vidare några till att utföra kraftgärningar, ytterligare några till att hava helbrägdagörelsens gåvor, eller till att taga sig an de hjälplösa, eller till att vara styresmän, eller till att på olika sätt tala tungomål.
Icke äro väl alla apostlar?
Icke äro väl alla profeter?
Icke äro väl alla lärare?
Icke utföra väl alla kraftgärningar?
Icke hava väl alla helbrägdagörelsens gåvor?
Icke tala väl alla tungomål?
Icke kunna väl alla uttyda?
Men varen ivriga att undfå de nådegåvor som äro de största.
Och nu vill jag ytterligare visa eder en väg, en övermåttan härlig väg.
Om jag talade både människors och änglars tungomål, men icke hade kärlek, så vore jag allenast en ljudande malm eller en klingande cymbal.
Och om jag hade profetians gåva och visste alla hemligheter och ägde all kunskap, och om jag hade all tro, så att jag kunde förflytta berg, men icke hade kärlek, så vore jag intet.
Och om jag gåve bort allt vad jag ägde till bröd åt de fattiga, ja, om jag offrade min kropp till att brännas upp, men icke hade kärlek, så vore detta mig till intet gagn.
Kärleken är tålig och mild.
Kärleken avundas icke, kärleken förhäver sig icke, den uppblåses icke.
Den skickar sig icke ohöviskt, den söker icke sitt, den förtörnas icke, den hyser icke agg för en oförrätts skull.
Den gläder sig icke över orättfärdigheten, men har sin glädje i sanningen.
Den fördrager allting, den tror allting, den hoppas allting, den uthärdar allting.
Kärleken förgår aldrig.
Men profetians gåva, den skall försvinna, och tungomålstalandet, det skall taga slut, och kunskapen, den skall försvinna.
Ty vår kunskap är ett styckverk, och vårt profeterande är ett styckverk;
men när det kommer, som är fullkomligt, då skall det försvinna, som är ett styckverk.
När jag var barn, talade jag såsom ett barn, mitt sinne var såsom ett barns, jag hade barnsliga tankar; men sedan jag blev man, har jag lagt bort vad barnsligt var.
Nu se vi ju på ett dunkelt sätt, såsom i en spegel, men då skola vi se ansikte mot ansikte.
Nu är min kunskap ett styckverk, men då skall jag känna till fullo, såsom jag själv har blivit till fullo känd.
Så bliva de då beståndande, tron, hoppet, kärleken, dessa tre; men störst bland dem är kärleken.
Faren efter kärleken, men varen ock ivriga att undfå de andliga gåvorna, framför allt profetians gåva.
Ty den som talar tungomål, han talar icke för människor, utan för Gud; ingen förstår honom ju, han talar i andehänryckning hemlighetsfulla ord.
Men den som profeterar, han talar för människor, dem till uppbyggelse och förmaning och tröst.
Den som talar tungomål uppbygger allenast sig själv, men den som profeterar, han uppbygger en hel församling.
Jag skulle väl vilja att I alla taladen tungomål, men ännu hellre ville jag att I profeteraden.
Den som profeterar är förmer än den som talar tungomål, om nämligen den senare icke därjämte uttyder sitt tal, så att församlingen får någon uppbyggelse.
Ja, mina bröder, om jag komme till eder och talade tungomål, vad gagn gjorde jag eder därmed, såframt jag icke därjämte genom mitt tal meddelade eder antingen någon uppenbarelse eller någon kunskap eller någon profetia eller någon undervisning?
Gäller det icke jämväl om livlösa ting som giva ljud ifrån sig, det må nu vara en flöjt eller en harpa, att vad som spelas på dem icke kan uppfattas, om de icke giva ifrån sig toner som kunna skiljas från varandra?
Likaså, om den signal som basunen giver är otydlig, vem gör sig då redo till strid?
Detsamma gäller nu för eder; om I icke med edra tungor frambringen begripliga ord, huru skall man då kunna förstå vad I talen?
Då bliver det ju ett tal i vädret.
Det finnes här i världen olika språk, vem vet huru många, och bland dem finnes intet vars ljud äro utan mening.
Men om jag nu icke förstår språket, så bliver jag en främling för den som talar, och den som talar bliver en främling för mig.
Detta gäller ock för eder; när I ären ivriga att undfå andliga gåvor, så må eder strävan efter att dessa hos eder skola överflöda hava församlingens uppbyggelse till mål.
Därför må den som talar tungomål bedja om att han ock må kunna uttyda.
Ty om jag talar tungomål, när jag beder, så beder visserligen min ande, men mitt förstånd kommer ingen frukt åstad.
Vad följer då härav?
Jo, jag skall väl bedja med anden, men jag skall ock bedja med förståndet; jag skall väl lovsjunga med anden, men jag skall ock lovsjunga med förståndet.
Eljest, om du lovar Gud med anden, huru skola de som sitta på de olärdas plats då kunna säga sitt »amen» till din tacksägelse?
De förstå ju icke vad du säger.
Om än din tacksägelse är god, så bliva de andra dock icke uppbyggda därav. --
Gud vare tack, jag talar tungomål mer än I alla;
och dock vill jag hellre i församlingen tala fem ord med mitt förstånd, till undervisning jämväl för andra, än tio tusen ord i tungomål.
Mina bröder, varen icke barn till förståndet; nej varen barn i ondskan, men varen fullmogna till förståndet.
Det är skrivet i lagen: »Genom människor med främmande tungomål och genom främlingars läppar skall jag tala till detta folk, men icke ens så skola de höra på mig, säger Herren.»
Alltså äro »tungomålen» ett tecken, ej för dem som tro, utan för dem som icke tro; profetian däremot är ett tecken, ej för dem som icke tro, utan för dem som tro.
Om nu hela församlingen komme tillhopa till gemensamt möte, och alla där talade tungomål, och så några som vore olärda komme ditin, eller några som icke trodde, skulle då icke dessa säga att I voren ifrån edra sinnen?
Om åter alla profeterade, och så någon som icke trodde, eller som vore olärd komme ditin, då skulle denne känna sig avslöjad av alla och av alla utrannsakad.
Vad som vore fördolt i hans hjärta bleve då uppenbart, och så skulle han falla ned på sitt ansikte och tillbedja Gud och betyga att »Gud verkligen är i eder».
Vad följer då härav, mina bröder?
Jo, när I kommen tillsammans, så har var och en något särskilt att meddela: den ene har en psalm, den andre något till undervisning, en annan åter någon uppenbarelse, en talar tungomål, en annan uttyder; allt detta må nu ske så, att det länder till uppbyggelse.
Vill man tala tungomål, så må för var gång två eller högst tre få tala, och av dessa en i sänder, och en må uttyda det.
Är ingen uttydare tillstädes, så må de tiga i församlingen och tala allenast för sig själva och för Gud.
Av dem som vilja profetera må två eller tre få tala, och de andra må döma om det som talas.
Men om någon annan som sitter där får en uppenbarelse, då må den förste tiga.
Ty I kunnen alla få profetera, den ene efter den andre, så att alla bliva undervisade och alla förmanade;
och profeters andar äro profeterna underdåniga.
Gud är ju icke oordningens Gud, utan fridens.
Såsom kvinnorna tiga i alla andra de heligas församlingar, så må de ock tiga i edra församlingar.
Det är dem icke tillstatt att tala, utan de böra underordna sig, såsom lagen bjuder.
Vilja de hava upplysning om något, så må de hemma fråga sina män; ty det är en skam för en kvinna att tala i församlingen. --
Eller är det från eder som Guds ord har utgått?
Eller har det kommit allenast till eder?
Om någon menar sig vara en profet eller en man med andegåva, så må han ock inse att vad jag skriver till eder är Herrens bud.
Men vill någon icke inse detta, så vare det hans egen sak.
Alltså, mina bröder, varen ivriga att undfå profetians gåva och förmenen ej heller någon att tala tungomål.
Men låten allt tillgå på höviskt sätt och med ordning.
Mina bröder, jag vill påminna eder om det evangelium som jag förkunnade för eder, som I jämväl togen emot, och som I ännu stån kvar i,
genom vilket I ock bliven frälsta; jag vill påminna eder om huru jag förkunnade det för eder, såframt I eljest hållen fast därvid -- om nu icke så är att I förgäves haven kommit till tro.
Jag meddelade eder ju såsom ett huvudstycke vad jag själv hade undfått: att Kristus dog för våra synder, enligt skrifterna,
och att han blev begraven, och att han har uppstått på tredje dagen, enligt skrifterna,
och att han visade sig för Cefas och sedan för de tolv.
Därefter visade han sig för mer än fem hundra bröder på en gång, av vilka de flesta ännu leva kvar, medan några äro avsomnade.
Därefter visade han sig för Jakob och sedan för alla apostlarna.
Allra sist visade han sig också för mig, som är att likna vid ett ofullgånget foster.
Ty jag är den ringaste bland apostlarna, ja, icke ens värdig att kallas apostel, jag som har förföljt Guds församling.
Men genom Guds nåd är jag vad jag är, och hans nåd mot mig har icke varit fåfäng, utan jag har arbetat mer än de alla -- dock icke jag, utan Guds nåd, som har varit med mig.
Det må nu vara jag eller de andra, så är det på det sättet vi predika, och på det sättet I haven kommit till tro.
Om det nu predikas om Kristus att han har uppstått från de döda, huru kunna då somliga bland eder säga att det icke finnes någon uppståndelse från de döda?
Om det åter icke finnes någon uppståndelse från de döda, då har icke heller Kristus uppstått.
Men om Kristus icke har uppstått, då är ju vår predikan fåfäng, då är ock eder tro fåfäng;
då befinnas vi ock vara falska Guds vittnen, eftersom vi hava vittnat mot Gud att han har uppväckt Kristus, som han icke har uppväckt, om det är sant att döda icke uppstå.
Ja, om döda icke uppstå, så har ej heller Kristus uppstått.
Men om Kristus icke har uppstått, så är eder tro förgäves; I ären då ännu kvar i edra synder.
Då hava ju ock de gått förlorade, som hava avsomnat i Kristus.
Om vi i detta livet hava i Kristus haft vårt hopp, och därav intet bliver, då äro vi de mest ömkansvärda av alla människor.
Men nu har Kristus uppstått från de döda, såsom förstlingen av de avsomnade.
Ty eftersom döden kom genom en människa, så kom ock genom en människa de dödas uppståndelse.
Och såsom i Adam alla dö, så skola ock i Kristus alla göras levande.
Men var och en i sin ordning: Kristus såsom förstlingen, därnäst, vid Kristi tillkommelse, de som höra honom till.
Därefter kommer änden, då när han överlämnar riket åt Gud och Fadern, sedan han från andevärldens alla furstar och alla väldigheter och makter har tagit all deras makt.
Ty han måste regera »till dess han har lagt alla sina fiender under sina fötter».
Sist bland hans fiender bliver ock döden berövad all sin makt;
ty »allt har han lagt under hans fötter».
Men när det heter att »allt är honom underlagt», då är uppenbarligen den undantagen, som har lagt allt under honom.
Och sedan allt har blivit Sonen underlagt, då skall ock Sonen själv giva sig under den som har lagt allt under honom.
Och så skall Gud bliva allt i alla.
Vad kunna annars de som låta döpa sig för de dödas skull vinna därmed?
Om så är att döda alls icke uppstå, varför låter man då döpa sig för deras skull?
Och varför undsätta vi oss själva var stund för faror?
Ty -- så sant jag i Kristus Jesus, vår Herre, kan berömma mig av eder, mina bröder -- jag lider döden dag efter dag.
Om jag hade tänkt såsom människor pläga tänka, när jag i Efesus kämpade mot vilddjuren, vad gagnade mig då det jag gjorde?
Om döda icke uppstå -- »låtom oss då äta och dricka, ty i morgon måste vi dö».
Faren icke vilse: »För goda seder dåligt sällskap är fördärv.»
Vaknen upp till rätt nykterhet, och synden icke.
Somliga finnas ju, som leva i okunnighet om Gud; eder till blygd säger jag detta.
Nu torde någon fråga: »På vad sätt uppstå då de döda, och med hurudan kropp skola de träda fram?»
Du oförståndige!
Det frö du sår, det får ju icke liv, om det icke först har dött.
Och när du sår, då är det du sår icke den växt som en gång skall komma upp, utan ett naket korn, kanhända ett vetekorn, kanhända något annat.
Men Gud giver det en kropp, en sådan som han vill, och åt vart frö dess särskilda kropp.
Icke allt kött är av samma slag, utan människors har sin art, boskapsdjurs kött en annan art, fåglars kött åter en annan, fiskars återigen en annan.
Så finnas ock både himmelska kroppar och jordiska kroppar, men de himmelska kropparnas härlighet är av ett slag, de jordiska kropparnas av ett annat slag.
En härlighet har solen, en annan härlighet har månen, åter en annan härlighet hava stjärnorna; ja, den ena stjärnan är icke lik den andra i härlighet. --
Så är det ock med de dödas uppståndelse: vad som bliver sått förgängligt, det uppstår oförgängligt;
vad som bliver sått i ringhet, det uppstår i härlighet; vad som bliver sått i svaghet, det uppstår i kraft;
här sås en »själisk» kropp, där uppstår en andlig kropp.
Så visst som det finnes en »själisk» kropp, så visst finnes det ock en andlig.
Så är ock skrivet: »Den första människan, Adam, blev en levande varelse med själ.»
Den siste Adam åter blev en levandegörande ande.
Men icke det andliga är det första, utan det »själiska»; sedan kommer det andliga.
Den första människan var av jorden och jordisk, den andra människan är av himmelen.
Sådan som den jordiska var, sådana äro ock de jordiska; och sådan som den himmelska är, sådana äro ock de himmelska.
Och såsom vi hava burit den jordiskas gestalt, så skola vi ock bära den himmelskas gestalt.
Mina bröder, vad jag nu vill säga är detta, att kött och blod icke kunna få Guds rike till arvedel; ej heller får förgängligheten oförgängligheten till arvedel.
Se, jag säger eder en hemlighet: Vi skola icke alla avsomna, men alla skola vi bliva förvandlade,
och det i ett nu, i ett ögonblick, vid den sista basunens ljud.
Ty basunen skall ljuda, och de döda skola uppstå till oförgänglighet, och då skola vi bliva förvandlade.
Ty detta förgängliga måste ikläda sig oförgänglighet, och detta dödliga ikläda sig odödlighet.
Men när detta förgängliga har iklätt sig oförgänglighet, och detta dödliga har iklätt sig odödlighet, då skall det ord fullbordas, som står skrivet: »Döden är uppslukad och seger vunnen.»
Du död, var är din seger?
Du död, var är din udd?
Dödens udd är synden, och syndens makt kommer av lagen.
Men Gud vare tack, som giver oss segern genom vår Herre Jesus Kristus!
Alltså, mina älskade bröder, varen fasta, orubbliga, alltid överflödande i Herrens verk, eftersom I veten att edert arbete icke är fåfängt i Herren.
Vad nu angår insamlingen till de heliga, så mån I förfara på samma sätt som jag har förordnat för församlingarna i Galatien.
Var och en av eder må spara ihop vad han får tillfälle till, och på första dagen i var vecka må han lägga av detta hemma hos sig, så att insamlingen icke göres först vid min ankomst.
Men när jag kommer, skall jag sända åstad de män som I själva pröven vara lämpliga, med brev till Jerusalem, för att där frambära eder kärleksgåva.
Och om saken befinnes vara värd att också jag reser, så skola de få åtfölja mig.
Jag tänker nämligen komma till eder, sedan jag har farit genom Macedonien.
Ty Macedonien vill jag allenast fara igenom,
men hos eder skall jag kanhända stanna något, möjligen vintern över, för att I därefter mån hjälpa mig till vägs, dit jag kan vilja begiva mig.
Jag vill icke besöka eder nu strax, på genomresa, ty jag hoppas att någon tid få stanna hos eder, om Herren så tillstädjer.
Men i Efesus vill jag stanna ända till pingst.
Ty en dörr till stor och fruktbärande verksamhet har öppnats för mig; jag har ock många motståndare.
Men när Timoteus kommer, så sen till, att han utan fruktan må kunna vistas hos eder.
Han utför ju Herrens verk, han såväl som jag;
må därför ingen förakta honom.
Hjälpen honom sedan till vägs i frid, så att han kommer åter till mig; ty jag väntar honom med bröderna.
Vad angår brodern Apollos, så har jag ivrigt uppmanat honom att med de andra bröderna begiva sig till eder.
Han var dock alls icke hågad att komma just nu; men när det bliver honom lägligt, skall han komma.
Vaken, stån fasta i tron, skicken eder såsom män, varen starka.
Låten allt hos eder ske i kärlek.
Mina bröder, jag vill giva eder en förmaning: I kännen ju Stefanas' husfolk och veten att de äro förstlingen i Akaja, och att de hava ägnat sig åt de heligas tjänst;
därför mån I å eder sida underordna eder under dessa män och under envar som bistår dem i deras arbete och själv gör sig möda.
Jag gläder mig över att Stefanas och Fortunatus och Akaikus hava kommit hit, ty dessa hava givit mig ersättning för vad jag har måst sakna genom att vara skild från eder;
de hava vederkvickt min ande såväl som eder ande.
Så lären eder nu att rätt uppskatta sådana män.
Församlingarna i provinsen Asien hälsar eder.
Akvila och Priska, tillika med den församling som kommer tillhopa i deras hus, hälsa eder mycket i Herren.
Ja, alla bröderna hälsa eder.
Hälsen varandra med en helig kyss.
Här skriver jag, Paulus, min hälsning med egen hand.
Om någon icke har Herren kär, så vare han förbannad.
Marana, ta!
Herren Jesu nåd vare med eder.
Min kärlek är med eder alla, i Kristus Jesus.
Paulus, genom Guds vilja Kristi Jesu apostel, så ock brodern Timoteus, hälsar den Guds församling som finnes i Korint, och tillika alla de heliga som finnas i hela Akaja.
Nåd vare med eder och frid ifrån Gud, vår Fader, och Herren Jesus Kristus.
Lovad vare vår Herres, Jesu Kristi, Gud och Fader, barmhärtighetens Fader och all trösts Gud,
han som tröstar oss i all vår nöd, så att vi genom den tröst vi själva undfå av Gud kunna trösta dem som äro stadda i allahanda nöd.
Ty såsom Kristuslidanden till överflöd komma över oss, så kommer ock genom Kristus tröst till oss i överflödande mått.
Men drabbas vi av nöd, så sker detta till tröst och frälsning för eder.
Undfå vi däremot tröst, så sker ock detta till tröst för eder, en tröst som skall visa sin kraft däri, att I ståndaktigt uthärden samma lidanden som vi utstå.
Och det hopp vi hysa i fråga om eder är fast,
ty vi veta att såsom I delen våra lidanden, så delen I ock den tröst vi undfå.
Vi vilja nämligen icke lämna eder, käre bröder, i okunnighet om vilken nöd vi fingo utstå i provinsen Asien, och huru övermåttan svårt det blev oss, utöver vår förmåga, så att vi till och med misströstade om livet.
Ja, vi hade redan i vårt inre likasom fått vår dödsdom, för att vi icke skulle förtrösta på oss själva, utan på Gud, som uppväcker de döda.
Och ur en sådan dödsnöd frälste han oss, och han skall än vidare frälsa oss; ja, till honom hava vi satt vårt hopp att han allt framgent skall frälsa oss.
Också I stån oss ju bi med eder förbön.
Och så skola många hembära tacksägelse för oss, för den nåd som genom mångas böner har kommit oss till del.
Ty vad vi kunna berömma oss av, och vad vårt samvete bär oss vittnesbörd om, det är att vi i denna världen hava vandrat i Guds helighet och renhet, icke ledda av köttslig vishet, utan av Guds nåd; så framför allt i vårt förhållande till eder.
Ty i vad vi skriva till eder ligger icke något annat än just vad I läsen och väl kunnen förstå.
Och jag hoppas att I skolen komma att till fullo förstå
vad I redan nu delvis förstån om oss: att vi äro eder berömmelse, likasom I ären vår berömmelse, på vår Herre Jesu dag.
Och i denna tillförsikt tänkte jag komma först till eder, för att I skullen få ännu ett kärleksbevis.
Genom eder stad ville jag alltså taga vägen till Macedonien, och jag skulle sedan från Macedonien återigen komma till eder, för att då av eder utrustas för resan till Judeen.
Så tänkte jag; och icke har jag väl därför nu handlat i vankelmod?
Eller plägar jag kanhända fatta mina beslut efter köttet, så att vad jag säger är på samma gång »ja, ja» och »nej, nej»?
Ingalunda; så sant Gud är trofast, vad vi tala till eder är icke »ja och nej».
Guds Son, Jesus Kristus, han som bland eder har blivit predikad genom oss -- genom mig och Silvanus och Timoteus -- han kom ju icke såsom »ja och nej», utan »ja» har kommit i och genom honom.
Ty Guds löften, så många de äro, hava i honom fått sitt »ja»; därför få de ock genom honom sitt »amen», på det att Gud må bliva ärad genom oss.
Men den som befäster oss såväl som eder i Kristus, och den som har smort oss, det är Gud,
han som har låtit oss undfå sitt insegel och givit oss Anden till en underpant i våra hjärtan.
Jag kallar Gud till vittne över min själ, att det är av skonsamhet mot eder som jag ännu icke har kommit till Korint.
(Detta säger jag icke, som om vi vore herrar över eder tro; fastmer äro vi edra medarbetare till att bereda eder glädje, ty i tron stån I fasta.)
Jag satte mig nämligen i sinnet att jag icke åter skulle komma till eder med bedrövelse.
Ty om jag bedrövade eder, vem skulle då bereda mig glädje?
Månne någon annan än den som genom mig hade blivit bedrövad?
Och vad jag skrev, det skrev jag, för att jag icke vid min ankomst skulle få bedrövelse från dem som jag borde få glädje av.
Ty jag har den tillförsikten till eder alla, att min glädje är allas eder glädje.
Och det var i stor nöd och hjärteångest, under många tårar, som jag skrev till eder, icke för att I skullen bliva bedrövade, utan för att I skullen förstå den synnerliga kärlek som jag har till eder.
Men om en viss man har vållat bedrövelse, så är det icke särskilt mig han har bedrövat, utan eder alla, i någon mån -- för att jag nu icke skall tala för strängt.
Nu är det likväl nog med den näpst som han har fått mottaga från de flesta bland eder.
I mån alltså nu tvärtom snarare förlåta och trösta honom, så att han icke till äventyrs går under genom sin alltför stora bedrövelse.
Därför uppmanar jag eder att fatta gemensamt beslut om att bemöta honom med kärlek.
Ty när jag skrev, var det just för att få veta huru I skullen hålla provet, huruvida I voren lydiga i allting.
Den som I förlåten något, honom förlåter ock jag, likasom jag också förut, om jag har haft något att förlåta, har inför Kristi ansikte förlåtit det för eder skull.
Jag vill nämligen icke att vi skola lida förfång av Satan; ty vad han har i sinnet, därom äro vi icke i okunnighet.
Jag kom till Troas för att förkunna evangelium om Kristus, och en dörr till verksamhet i Herren öppnades för mig;
men jag fick ingen ro i min ande, ty jag fann icke där min broder Titus.
Jag tog då avsked av dem som voro där och begav mig till Macedonien.
Men Gud vare tack, som i Kristus alltid för oss fram i segertåg och genom oss allestädes utbreder hans kunskaps vällukt!
Ty vi äro en Kristi välluktande rökelse inför Gud, både ibland dem som bliva frälsta och ibland dem som gå förlorade.
För dessa senare äro vi en lukt från död till död; för de förra äro vi en lukt från liv till liv.
Vem är nu skicklig härtill?
Jo, vi förfalska ju icke av vinningslystnad Guds ord, såsom så många andra göra; utan av rent sinne, drivna av Gud, förkunna vi ordet i Kristus, inför Gud.
Begynna vi nu åter att anbefalla oss själva?
Eller behöva vi kanhända, såsom somliga, ett anbefallningsbrev till eder?
Eller kanhända ifrån eder?
Nej, I ären själva vårt brev, ett brev som är inskrivet i våra hjärtan, känt och läst av alla människor.
Ty det är uppenbart att I ären ett Kristus-brev, avfattat genom oss, skrivet icke med bläck, utan med den levande Gudens Ande, icke på tavlor av sten, utan på tavlor av kött, på människohjärtan.
En sådan tillförsikt hava vi genom Kristus till Gud.
Icke som om vi av oss själva vore skickliga att tänka ut något, såsom komme det från oss själva, utan den skicklighet vi hava kommer från Gud,
som också har gjort oss skickliga till att vara tjänare åt ett nytt förbund, ett som icke är bokstav, utan är ande; ty bokstaven dödar, men Anden gör levande.
Om nu redan dödens ämbete, som var med bokstäver inristat på stenar, framträdde i härlighet, så att Israels barn icke kunde se på Moses' ansikte för hans ansiktes härlighets skull, vilken dock var försvinnande,
huru mycket större härlighet skall då icke Andens ämbete hava!
Ty om redan fördömelsens ämbete var härligt, så måste rättfärdighetens ämbete ännu mycket mer överflöda av härlighet.
Ja, en så översvinnlig härlighet har detta ämbete, att vad som förr hade härlighet här visar sig vara utan all härlighet.
Ty om redan det som var försvinnande framträdde i härlighet, så måste det som bliver beståndande hava en ännu mycket större härlighet.
Då vi nu hava ett sådant hopp, gå vi helt öppet till väga
och göra icke såsom Moses, vilken hängde ett täckelse för sitt ansikte, så att Israels barn icke kunde se huru det som var försvinnande tog en ände.
Men deras sinnen blevo förstockade.
När det gamla förbundets skrifter föreläsas, hänger ju ännu i denna dag samma täckelse oborttaget kvar; ty först i Kristus försvinner det.
Ja, ännu i dag hänger ett täckelse över deras hjärtan, då Moses föreläses.
Men när de en gång omvända sig till Herren, tages täckelset bort.
Och Herren är Anden, och där Herrens Ande är, där är frihet.
Men vi alla som med avhöljt ansikte återspegla Herrens härlighet, vi förvandlas till hans avbilder, i det vi stiga från den ena härligheten till den andra, såsom när den Herre verkar, som själv är ande.
Därför, då vi nu, genom den barmhärtighet som har vederfarits oss, hava detta ämbete, så fälla vi icke modet.
Nej, vi hava frånsagt oss allt skamligt hemlighetsväsen och gå icke illfundigt till väga, ej heller förfalska vi Guds ord, utan framlägga öppet sanningen och anbefalla oss så, inför Gud, hos var människas samvete.
Och om vårt evangelium nu verkligen är bortskymt av ett täckelse, så finnes det täckelset hos dem som gå förlorade.
Ty de otrognas sinnen har denna tidsålders gud så förblindat, att de icke se det sken som utgår från evangelium om Kristi, Guds egen avbilds, härlighet.
Vi predika ju icke oss själva, utan Kristus Jesus såsom Herre, och oss såsom tjänare åt eder, för Jesu skull.
Ty den Gud som sade: »Ljus skall lysa fram ur mörkret», han är den som har låtit ljus gå upp i våra hjärtan, för att kunskapen om Guds härlighet, som strålar fram i Kristi ansikte, skall kunna sprida sitt sken.
Men denna skatt hava vi i lerkärl, för att den översvinnliga kraften skall befinnas vara Guds och icke något som kommer från oss.
Vi äro på allt sätt i trångmål, dock icke utan utväg; vi äro rådvilla, dock icke rådlösa;
vi äro förföljda, dock icke givna till spillo; vi äro slagna till marken, dock icke förlorade.
Alltid bära vi Jesu dödsmärken på vår kropp, för att också Jesu liv skall bliva uppenbarat i vår kropp.
Ja, ännu medan vi leva, överlämnas vi för Jesu skull beständigt åt döden, på det att ock Jesu liv må bliva uppenbarat i vårt dödliga kött.
Så utför nu döden sitt verk i oss, men i eder verkar livet.
Men såsom det är skrivet: »Jag tror, därför talar jag ock», så tro också vi, eftersom vi hava samma trons Ande; därför tala vi ock,
ty vi veta att han som uppväckte Herren Jesus, han skall ock uppväcka oss med Jesus och ställa oss inför sig tillsammans med eder.
Allt sker nämligen för eder skull, på det att nåden, genom att komma allt flera till del, må bliva så mycket större och verka en allt mer överflödande tacksägelse, Gud till ära.
Därför fälla vi icke modet; om ock vår utvärtes människa förgås, så förnyas likväl vår invärtes människa dag efter dag.
Ty vår bedrövelse, som varar ett ögonblick och väger föga, bereder åt oss, i översvinnligen rikt mått, en härlighet som väger översvinnligen tungt och varar i evighet --
åt oss som icke hava till ögonmärke de ting som synas, utan dem som icke synas; ty de ting som synas, de vara allenast en tid, med de som icke synas, de vara i evighet.
Ty vi veta, att om vår kroppshydda, vår jordiska boning, nedbrytes, så hava vi en byggnad som kommer från Gud, en boning som icke är gjord med händer, en evig boning i himmelen.
Därför sucka vi ju ock av längtan att få överkläda oss med vår himmelska hydda;
ty hava vi en gång iklätt oss denna, skola vi sedan icke komma att befinnas nakna.
Ja, vi som ännu leva här i kroppshyddan, vi sucka och äro betungade, eftersom vi skulle vilja undgå att avkläda oss och i stället få överkläda oss, så att det som är dödligt bleve uppslukat av livet.
Och den som har berett oss till just detta, det är Gud, som till en underpant har givit oss Anden.
Så äro vi då alltid vid gott mod.
Vi veta väl att vi äro borta ifrån Herren, så länge vi äro hemma i kroppen;
ty vi vandra här i tro och icke i åskådning.
Men vi äro vid gott mod och skulle helst vilja flytta bort ifrån kroppen och komma hem till Herren.
Därför söka vi ock vår ära i att vara honom till behag, vare sig vi äro hemma eller borta.
Ty vi måste alla, sådana vi äro, träda fram inför Kristi domstol, för att var och en skall få igen sitt jordelivs gärningar, alltefter som han har handlat, vare sig han har gjort gott eller ont.
Då vi alltså veta vad det är att frukta Herren, söka vi att »vinna människor», men för Gud är det uppenbart hurudana vi äro; och jag hoppas att det också är uppenbart för edra samveten.
Vi vilja nu ingalunda åter anbefalla oss själva hos eder, men vi vilja giva eder en anledning att berömma eder i fråga om oss, så att I haven något att svara dem som berömma sig av utvärtes ting och icke av vad som är i hjärtat.
Ty om vi hava varit »från våra sinnen», så har det varit i Guds tjänst; om vi åter äro vid lugn besinning, så är det eder till godo.
Ty Kristi kärlek tvingar oss, eftersom vi tänka så: en har dött för alla, alltså hava de alla dött.
Och han har dött för alla, på det att de som leva icke mer må leva för sig själva, utan leva för honom som har dött och uppstått för dem.
Allt ifrån denna tid veta vi därför för vår del icke av någon efter köttet.
Och om vi än efter köttet hade lärt känna Kristus, så känna vi honom nu icke mer på det sättet.
Alltså, om någon är i Kristus, så är han en ny skapelse.
Det gamla är förgånget; se, något nytt har kommit!
Men alltsammans kommer från Gud, som har försonat oss med sig själv genom Kristus och givit åt oss försoningens ämbete.
Ty det var Gud som i Kristus försonade världen med sig själv; han tillräknar icke människorna deras synder, och han har betrott oss med försoningens ord.
Å Kristi vägnar äro vi alltså sändebud; det är Gud som förmanar genom oss.
Vi bedja å Kristi vägnar: Låten försona eder med Gud.
Den som icke visste av någon synd, honom har han för oss gjort till synd, på det att vi i honom må bliva rättfärdighet från Gud.
Men såsom medarbetare förmana vi eder ock att icke så mottaga Guds nåd, att det bliver utan frukt.
Han säger ju: »Jag bönhör dig i behaglig tid, och jag hjälper dig på frälsningens dag.»
Se, nu är den välbehagliga tiden; se, nu är frälsningens dag.
Härvid vilja vi icke i något stycke vara till någon anstöt, på det att vårt ämbete icke må bliva smädat.
Fastmer vilja vi i allting bevisa oss såsom Guds tjänare, i mycken ståndaktighet, under bedrövelse och nöd och ångest,
under hugg och slag, under fångenskap och upprorslarm, under mödor, vakor och svält,
i renhet, i kunskap, i tålamod och godhet, i helig ande, i oskrymtad kärlek,
med sanning i vårt tal, med kraft från Gud, med rättfärdighetens vapen både i högra handen och i vänstra,
under ära och smälek, under ont rykte och gott rykte, såsom villolärare, då vi dock äro sannfärdiga,
såsom okända, fastän vi äro väl kända, såsom döende, men se, vi leva, såsom tuktade, men likväl icke till döds,
såsom bedrövade, men dock alltid glada, såsom fattiga, medan vi dock göra många rika, såsom utblottade på allt, men likväl ägande allt.
Vi hava nu upplåtit vår mun och talat öppet till eder, I korintier.
Vårt hjärta har vidgat sig för eder.
Ja, det rum I haven i vårt inre är icke litet, men i edra hjärtan är allenast litet rum.
Given oss då lika för lika -- om jag nu får tala såsom till barn -- ja, vidgen också I edra hjärtan.
Gån icke i ok tillsammans med dem som icke tro; det bleve omaka par.
Vad har väl rättfärdighet att skaffa med orättfärdighet, eller vilken gemenskap har ljus med mörker?
Huru förlika sig Kristus och Beliar, eller vad delaktighet har den som tror med den som icke tror?
Eller huru låter ett Guds tempel förena sig med avgudar?
Vi äro ju ett den levande Gudens tempel, ty Gud har sagt: »Jag skall bo i dem och vandra ibland dem; jag skall vara deras Gud, och de skola vara mitt folk.»
Alltså: »Gån ut ifrån dem och skiljen eder ifrån dem, säger Herren; kommen icke vid det orent är.
Då skall jag taga emot eder
och vara en Fader för eder; och I skolen vara mina söner och döttrar, säger Herren, den Allsmäktige.»
Då vi nu hava dessa löften, mina älskade, så låtom oss rena oss från allt som befläckar vare sig kött eller ande, i det vi fullborda vår helgelse i Guds fruktan.
Bereden oss ett rum i edra hjärtan; vi hava icke handlat orätt mot någon, icke varit någon till skada, icke gjort någon något förfång. --
Jag säger icke detta för att döma eder; jag har ju redan sagt att I haven ett rum i vårt hjärta, så att vi skola både dö och leva med varandra.
Stor är den tillit som jag har till eder, mycket berömmer jag mig av eder; jag har fått hugnad i fullt mått och glädje i rikt överflöd, mitt i allt vårt betryck.
Ty väl fingo vi till köttet ingen ro, icke ens sedan vi hade kommit till Macedonien, utan vi voro på allt sätt i trångmål, utifrån genom strider, inom oss genom farhågor;
men Gud, som tröstar dem som äro betryckta, han tröstade oss genom Titus' ankomst,
och icke allenast genom hans ankomst, utan ock därigenom att han hade fått så mycken hugnad av eder.
Han omtalade nämligen för oss eder längtan, eder klagan, eder iver i fråga om mig; och så gladde jag mig ännu mer.
Ty om jag ock bedrövade eder genom mitt brev, så ångrar jag nu icke detta.
Nej, om jag förut ångrade det -- eftersom jag ser att det brevet har bedrövat eder, låt vara allenast för en liten tid --
så gläder jag mig nu i stället, icke därför att I bleven bedrövade, utan därför att eder bedrövelse lände eder till bättring.
Det var ju efter Guds sinne som I bleven bedrövade, och I haven alltså icke genom oss lidit någon skada.
Ty den bedrövelse som är efter Guds sinne kommer åstad en bättring som leder till frälsning, och som man icke ångrar; men världens bedrövelse kommer åstad död.
Se, just detta, att I bleven bedrövade efter Guds sinne, huru mycket nit har det icke framkallat hos eder, ja, huru många ursäkter, huru stor förtrytelse, huru mycken fruktan, huru mycken längtan, huru mycken iver, huru många bestraffningar!
På allt sätt haven I bevisat att I viljen vara rena i den sak det här gäller. --
Om jag skrev till eder, så skedde detta alltså icke för den mans skull, som hade gjort orätt, ej heller för den mans skull, som hade lidit orätt, utan på det att edert nit för oss skulle bliva uppenbart bland eder själva inför Gud.
Så hava vi nu fått hugnad.
Och till den hugnad, som vi redan för egen del fingo, kom den ännu mer överflödande glädje som bereddes oss av den glädje Titus hade fått.
Ty hans ande har fått vederkvickelse genom eder alla.
Och om jag inför honom har berömt mig något i fråga om eder, så har jag icke kommit på skam därmed; utan likasom vi eljest i allting hava talat sanning inför eder, så har också det som vi inför Titus hava sagt till eder berömmelse visat sig vara sanning.
Och hans hjärta överflödar ännu mer av kärlek till eder, då han nu påminner sig allas eder lydnad, huru I villigt togen emot honom, med fruktan och bävan.
Jag gläder mig över att jag, i allt vad eder angår, kan vara vid gott mod.
Vi vilja meddela eder, käre bröder, huru Guds nåd har verkat i Macedoniens församlingar.
Fastän de hava varit prövade av svår nöd, har deras överflödande glädje, mitt under deras djupa fattigdom, så flödat över, att de av gott hjärta hava givit rikliga gåvor.
Ty de hava givit efter sin förmåga, ja, över sin förmåga, och det självmant; därom kan jag vittna.
Mycket enträget bådo de oss om den ynnesten att få vara med om understödet åt de heliga.
Och de gåvo icke allenast vad vi hade hoppats, utan sig själva gåvo de, först och främst åt Herren, och så åt oss, genom Guds vilja.
Så kunde vi uppmana Titus att han skulle fortsätta såsom han hade begynt och föra jämväl detta kärleksverk bland eder till fullbordan.
Ja, då I nu utmärken eder i alla stycken: i tro, i tal, i kunskap, i allsköns nit, i kärlek, den kärlek som av eder har blivit oss bevisad, så mån I se till, att I också utmärken eder i detta kärleksverk.
Detta säger jag dock icke såsom en befallning, utan därför att jag, genom att framhålla andras nit, vill pröva om också eder kärlek är äkta.
I kännen ju vår Herres, Jesu Kristi, nåd, huru han, som var rik, likväl blev fattig för eder skull, på det att I genom hans fattigdom skullen bliva rika.
Det är allenast ett råd som jag härmed giver.
Ty detta kan vara nyttigt för eder.
I voren ju före de andra -- redan under förra året -- icke allenast när det gällde att sätta saken i verket, utan till och med när det gällde att besluta sig för den.
Fullborden nu ock edert verk, så att I, som voren så villiga att besluta det, jämväl, i mån av edra tillgångar, fören det till fullbordan.
Ty om den goda viljan är för handen, så bliver den välbehaglig med de tillgångar den har och bedömes ej efter vad den icke har.
Ty meningen är icke att andra skola hava lättnad och I själva lida nöd.
Nej, en utjämning skall ske,
så att edert överflöd denna gång kommer deras brist till hjälp, för att en annan gång deras överflöd skall komma eder brist till hjälp.
Så skall en utjämning ske,
efter skriftens ord: »Den som hade samlat mycket hade intet till överlopps, och den som hade samlat litet, honom fattades intet.»
Gud vare tack, som också i Titus' hjärta ingiver samma nit för eder.
Ty han mottog villigt vår uppmaning; ja, han var så nitisk, att han nu självmant far åstad till eder.
Med honom sända vi ock här en broder som i alla våra församlingar prisas för sitt nit om evangelium;
dessutom har han ock av församlingarna blivit utvald att vara vår följeslagare, när vi skola begiva oss åstad med den kärleksgåva som nu genom vår försorg kommer till stånd, Herren till ära och såsom ett vittnesbörd om vår goda vilja.
Därmed vilja vi förebygga att man talar illa om oss, i vad som rör det rikliga sammanskott som nu genom vår försorg kommer till stånd.
Ty vi vinnlägga oss om vad som är gott icke allenast inför Herren, utan ock inför människor.
Jämte dessa sända vi en annan av våra bröder, vilkens nit vi ofta och i många stycken hava funnit hålla provet, och som nu på grund av sin stora tillit till eder är ännu mycket mer nitisk.
Om jag nu har anbefallt Titus, så mån I besinna att han är min medbroder och min medarbetare till edert bästa; och om jag har skrivit om andra våra bröder, så mån I besinna att de äro församlingssändebud och Kristi ära.
Given alltså inför församlingarna bevis på eder kärlek, och därmed också på sanningen av det som vi inför dem hava sagt till eder berömmelse.
Om understödet till de heliga är det nu visserligen överflödigt att jag här skriver till eder;
jag känner ju eder goda vilja, och av den plägar jag, i fråga om eder, berömma mig inför macedonierna, i det jag omtalar att Akaja ända sedan förra året har varit redo, och att det är just edert nit som har eggat så många andra.
Likväl sänder jag nu åstad dessa bröder, för att det som jag har sagt till eder berömmelse icke skall i denna del befinnas hava varit tomt tal.
Ty, såsom jag förut har sagt, jag vill att I skolen vara redo.
Eljest, om några macedonier komma med mig och finna eder oberedda, kunna vi -- för att icke säga I -- till äventyrs komma på skam med vår tillförsikt i denna sak.
Jag har därför funnit det vara nödvändigt att uppmana bröderna att i förväg begiva sig till eder och förbereda den rikliga »välsignelsegåva» som I redan haven utlovat.
De skola laga att denna är tillreds såsom en riklig gåva, och icke såsom en gåva i njugghet.
Besinnen detta: den som sår sparsamt, han skall ock skörda sparsamt; men den som sår rikligt, han skall ock skörda riklig välsignelse.
Var och en give efter som han har känt sig manad i sitt hjärta, icke med olust eller av tvång, ty »Gud älskar en glad givare».
Men Gud är mäktig att i överflödande mått låta all nåd komma eder till del, så att I alltid i allo haven allt till fyllest och i överflöd kunnen giva till allt gott verk,
efter skriftens ord: »Han utströr, han giver åt de fattiga, hans rättfärdighet förbliver evinnerligen.»
Och han som giver såningsmannen »säd till att så och bröd till att äta», han skall ock giva eder utsädet och låta det föröka sig och skall bereda växt åt eder rättfärdighets frukt.
I skolen bliva så rika på allt, att I av gott hjärta kunnen giva allahanda gåvor, vilka, när de överlämnas genom oss, skola framkalla tacksägelse till Gud.
Ty det understöd, som kommer till stånd genom denna eder tjänst, skall icke allenast avhjälpa de heligas brist, utan verka ännu långt mer genom att framkalla många tacksägelser till Gud.
De skola nämligen, därför att I visen eder så väl hålla provet i fråga om detta understöd, komma att prisa Gud för att I med så lydaktigt sinne bekännen eder till Kristi evangelium och av så gott hjärta visen dem och alla andra edert deltagande.
De skola ock själva bedja för eder och längta efter eder, för den Guds nåds skull, som i så översvinnligen rikt mått beskäres eder.
Ja, Gud vare tack för hans outsägligt rika gåva!
Jag Paulus själv, som »är så ödmjuk, när jag står ansikte mot ansikte med eder, men visar mig så modig mot eder, när jag är långt borta», jag förmanar eder vid Kristi saktmod och mildhet
och beder eder se till, att jag icke, när jag en gång är hos eder, måste »visa mig modig», i det jag helt oförskräckt tänker våga mig på somliga som mena att vi »vandra efter köttet».
Ty fastän vi vandra i köttet, föra vi dock icke en strid efter köttet.
Våra stridsvapen äro nämligen icke av köttslig art; de äro tvärtom så mäktiga inför Gud, att de kunna bryta ned fästen.
Ja, vi bryta ned tankebyggnader och alla slags höga bålverk, som uppresas mot kunskapen om Gud, och vi taga alla slags tankefunder till fånga och lägga dem under Kristi lydnad.
Och när lydnaden fullt har kommit till väldet bland eder, då äro vi redo att näpsa all olydnad.
Sen då vad som ligger öppet för allas ögon.
Om någon i sitt sinne är viss om att han hör Kristus till, så må han ytterligare besinna inom sig, att lika visst som han själv hör Kristus till, lika visst göra också vi det.
Och om jag än något härutöver berömmer mig, då nu fråga är om vår myndighet -- den som Herren har givit oss, till att uppbygga eder och icke till att nedbryta -- så skall jag dock icke komma på skam därmed.
Jag vill icke att det skall se ut, som om jag med mina brev allenast tänkte skrämma eder.
Ty man säger ju: »Hans brev äro väl myndiga och stränga, men när han kommer själv, uppträder han utan kraft, och på hans ord aktar ingen.»
Den som säger sådant, han må emellertid göra sig beredd på att sådana som vi äro i orden, genom våra brev, när vi äro frånvarande, sådana skola vi ock visa oss i gärningarna, när vi äro närvarande.
Ty vi äro icke nog dristiga att räkna oss till eller jämföra oss med somliga som giva sig själva gott vitsord, men som äro utan förstånd, i det att de mäta sig allenast efter sig själva och jämföra sig allenast med sig själva.
Vi för vår del vilja icke berömma oss till övermått, utan allenast efter måttet av det område som Gud tillmätte åt oss, när han bestämde att vi skulle nå fram jämväl till eder.
Ty vi sträcka oss icke utom vårt område, såsom nådde vi icke rätteligen fram till eder; vi hava ju redan med evangelium om Kristus hunnit fram jämväl till eder.
När vi säga detta, berömma vi oss icke till övermått, icke av andras arbete.
Men väl hava vi det hoppet, att i samma mån som eder tro växer till, vi inom det område som har tillfallit oss skola bland eder vinna framgång, i så överflödande mått,
att vi också få förkunna evangelium i trakter som ligga bortom eder -- och detta utan att vi, inom ett område som tillhör andra, berömma oss i fråga om det som redan där är uträttat.
Men »den som vill berömma sig, han berömme sig av Herren».
Ty icke den håller provet, som giver sig själv gott vitsord, utan den som Herren giver sådant vitsord.
Jag skulle önska att I villen hava fördrag med mig, om jag nu talar något litet efter dårars sätt.
Dock, I haven helt visst fördrag med mig.
Ty jag nitälskar för eder såsom Gud nitälskar, och jag har trolovat eder med Kristus, och ingen annan, för att kunna ställa fram inför honom en ren jungfru.
Men jag fruktar att såsom ormen i sin illfundighet bedrog Eva, så skola till äventyrs också edra sinnen fördärvas och dragas ifrån den uppriktiga troheten mot Kristus.
Om någon kommer och predikar en annan Jesus, än den vi hava predikat, eller om I undfån ett annat slags ande, än den I förut haven undfått, eller ett annat slags evangelium, än det I förut haven mottagit, då fördragen I ju sådant alltför väl.
Jag menar nu att jag icke i något stycke står tillbaka för dessa så övermåttan höga »apostlar».
Om jag än är oförfaren i talkonsten, så är jag det likväl icke i fråga om kunskap.
Tvärtom, vi hava på allt sätt, i alla stycken, lagt vår kunskap i dagen inför eder.
Eller var det väl en synd jag begick, när jag för intet förkunnade Guds evangelium för eder och sålunda ödmjukade mig, på det att I skullen bliva upphöjda?
Andra församlingar plundrade jag, i det jag, för att kunna tjäna eder, tog lön av dem.
Och när jag under min vistelse hos eder led brist, låg jag ändå ingen till last; ty den brist jag led avhjälptes av bröderna, när de kommo från Macedonien.
Ja, på allt sätt aktade jag mig för att vara eder till tunga, och allt framgent skall jag akta mig därför.
Så visst som Kristi sannfärdighet är i mig, den berömmelsen skall icke få tagas ifrån mig i Akajas bygder.
Varför?
Månne därför att jag icke älskar eder?
Gud vet att jag så gör.
Och vad jag nu gör, det skall jag ock framgent göra, för att de som trakta efter tillfälle att bliva likställda med oss i fråga om berömmelse skola genom mig berövas tillfället därtill.
Ty de männen äro falska apostlar, oredliga arbetare, som förskapa sig till Kristi apostlar.
Och detta är icke att undra på.
Satan själv förskapar sig ju till en ljusets ängel.
Det är då icke något märkligt, om jämväl hans tjänare så förskapa sig, att de likna rättfärdighetens tjänare.
Men deras ände skall svara emot deras gärningar.
Åter säger jag: Ingen må mena att jag är en dåre; men om jag vore det, så mån I ändå hålla till godo med mig -- låt vara såsom med en dåre -- så att ock jag får berömma mig något litet.
Vad jag talar, då jag nu med sådan tillförsikt berömmer mig, det talar jag icke efter Herrens sinne, utan efter dårars sätt.
Då så många berömma sig på köttsligt vis, vill ock jag berömma mig;
I haven ju gärna fördrag med dårar, I som själva ären så kloka.
I fördragen ju, om man trälbinder eder, om man utsuger eder, om man fångar eder, om man förhäver sig över eder, om man slår eder i ansiktet.
Till vår skam måste jag tillstå att vi för vår del hava »varit för svaga» till sådant.
Men eljest, vadhelst andra kunna göra sig stora med, det kan också jag göra mig stor med -- om jag nu får tala efter dårars sätt.
Äro de hebréer, så är jag det ock.
Äro de israeliter, så är jag det ock.
Äro de Abrahams säd, så är jag det ock.
Äro de Kristi tjänare, så är jag det ännu mer -- om jag nu får tala såsom vore jag en dåre.
Jag har haft mer arbete, oftare varit i fängelse, fått hugg och slag till överflöd, varit i dödsnöd många gånger.
Av judarna har jag fem gånger fått fyrtio slag, på ett när.
Tre gånger har jag blivit piskad med spön, en gång har jag blivit stenad, tre gånger har jag lidit skeppsbrott, ett helt dygn har jag drivit omkring på djupa havet.
Jag har ofta måst vara ute på resor; jag har utstått faror på floder, faror bland rövare, faror genom landsmän, faror genom hedningar, faror i städer, faror i öknar, faror på havet, faror bland falska bröder --
allt under arbete och möda, under mångfaldiga vakor, under hunger och törst, under svält titt och ofta, under köld och nakenhet.
Och till allt annat kommer det, att jag var dag är överlupen, då jag måste hava omsorg om alla församlingarna.
Vem är svag, utan att också jag bliver svag?
Vem kommer på fall, utan att jag bliver upptänd? --
Om jag nu måste berömma mig, så vill jag berömma mig av min svaghet.
Herren Jesu Gud och Fader, han som är högtlovad i evighet, vet att jag icke ljuger.
I Damaskus lät konung Aretas' ståthållare sätta ut vakt vid damaskenernas stad för att gripa mig;
och jag måste i en korg släppas ned genom en öppning på muren och kom så undan hans händer.
Jag måste ytterligare berömma mig.
Väl är sådant icke eljest nyttigt, men jag kommer nu till syner och uppenbarelser, som hava beskärts mig av Herren.
Jag vet om en man som är i Kristus, att han för fjorton år sedan blev uppryckt ända till tredje himmelen; huruvida det nu var i kroppslig måtto, eller om han var skild från sin kropp, det vet jag icke, Gud allena vet det.
Ja, jag vet om denne man, att han -- huruvida det nu var i kroppslig måtto, eller om han var skild från sin kropp, det vet jag icke, Gud allena vet det --
jag vet om honom, att han blev uppryckt till paradiset och fick höra outsägliga ord, sådana som det icke är lovligt för en människa att uttala.
I fråga om den mannen vill jag berömma mig, men i fråga om mig själv vill jag icke berömma mig, om icke av min svaghet.
Visserligen skulle jag icke vara en dåre, om jag ville berömma mig själv, ty det vore sanning som jag då skulle tala; men likväl avhåller jag mig därifrån, för att ingen skall hava högre tankar om mig än skäligt är, efter vad han ser hos mig eller hör av mig.
Och för att jag icke skall förhäva mig på grund av mina övermåttan höga uppenbarelser, har jag fått en törntagg i mitt kött, en Satans ängel, som skall slå mig i ansiktet, för att jag icke skall förhäva mig.
Att denne måtte vika ifrån mig, därom har jag tre gånger bett till Herren.
Men Herren har sagt till mig; »Min nåd är dig nog, ty kraften fullkomnas i svaghet.»
Därför vill jag hellre med glädje berömma mig av min svaghet, på det att Kristi kraft må komma och vila över mig.
Ja, därför finner jag behag i svaghet, i misshandling, i nöd, i förföljelse, i ångest för Kristi skull; ty när jag är svag, då är jag stark.
Så har jag nu gjort mig till en dåre; I haven själva nödgat mig därtill.
Jag hade ju bort få gott vitsord av eder; ty om jag än är ett intet, så har jag dock icke i något stycke stått tillbaka för dessa så övermåttan höga »apostlar».
De gärningar som äro en apostels kännemärken hava ock med all uthållighet blivit gjorda bland eder, genom tecken och under och kraftgärningar.
Och haven I väl i något stycke blivit tillbakasatta för de andra församlingarna?
Dock, kanhända i det stycket, att jag för min del icke har legat eder till last?
Den oförrätten mån I då förlåta mig.
Se, det är nu tredje gången som jag står redo att komma till eder.
Och jag skall icke ligga eder till last, ty icke edert söker jag, utan eder själva.
Och barnen äro ju icke pliktiga att spara åt föräldrarna, utan föräldrarna åt barnen.
Och för min del vill jag gärna för edra själar både offra vad jag äger och låta mig själv offras hel och hållen.
Om jag nu så högt älskar eder, skall jag väl därför bliva mindre älskad?
Dock, det kunde ju vara så, att jag visserligen icke själv hade betungat eder, men att jag på en listig omväg hade fångat eder, jag som är så illfundig.
Har jag då verkligen, genom någon av dem som jag har sänt till eder, berett mig någon orätt vinning av eder?
Sant är att jag bad Titus fara och sände med honom den andre brodern.
Men icke har väl Titus berett mig någon orätt vinning av eder?
Hava vi icke båda vandrat i en och samme Ande?
Hava vi icke båda gått i samma fotspår?
Nu torden I redan länge hava menat att det är inför eder som vi försvara oss.
Nej, det är inför Gud, i Kristus, som vi tala, men visserligen alltsammans för att uppbygga eder, I älskade.
Ty jag fruktar att jag vid min ankomst till äventyrs icke skall finna eder sådana som jag skulle önska, och att jag själv då av eder skall befinnas vara sådan som I icke skullen önska.
Jag fruktar att till äventyrs kiv, avund, vrede, genstridighet, förtal, skvaller, uppblåsthet och oordning råda bland eder.
Ja, jag fruktar att min Gud skall låta mig vid min ankomst åter bliva förödmjukad genom eder, och att jag skall få sörja över många av dem som förut hava syndat, och som ännu icke hava känt ånger över den orenhet och otukt och lösaktighet som de hava övat.
Det är nu tredje gången som jag skall komma till eder; »efter två eller tre vittnens utsago skall var sak avgöras».
Till dem som förut hava syndat och till alla de andra har jag redan i förväg sagt, och jag säger nu åter i förväg -- nu då jag är borta ifrån eder, likasom förut då jag för andra gången var hos eder -- att jag icke skall visa någon skonsamhet, när jag kommer igen.
I viljen ju hava ett bevis för att det är Kristus som talar i mig, han som icke är svag mot eder, utan är stark bland eder.
Ty om han än blev korsfäst i följd av svaghet, så lever han dock av Guds kraft.
Också vi äro ju svaga i honom, men av Guds kraft skola vi leva med honom och bevisa det på eder.
Rannsaken eder själva, huruvida I ären i tron, ja, pröven eder själva.
Eller kännen I icke med eder själva att Jesus Kristus är i eder?
Varom icke, så hållen I ej provet.
Att vi för vår del icke äro av dem som ej hålla provet, det hoppas jag att I skolen få lära känna.
Men vi bedja till Gud att I icke mån göra något ont, detta icke för att vi å vår sida skola synas hålla provet, utan för att I själva verkligen skolen göra vad gott är.
Sedan må vi å vår sida gärna anses icke hålla provet.
Ty icke mot sanningen, utan allenast för sanningen förmå vi något.
Och vi glädja oss, när vi äro svaga, men I ären starka.
Just detta bedja vi också om, att I mån alltmer fullkomnas.
Och medan jag ännu är borta ifrån eder, skriver jag detta, för att jag icke, när jag är hos eder, skall nödgas uppträda med stränghet, i kraft av den myndighet som Herren har givit mig, till att uppbygga och icke till att nedbryta.
För övrigt, mina bröder, varen glada, låten fullkomna eder, låten förmana eder, varen ens till sinnes, hållen frid; då skall kärlekens och fridens Gud vara med eder.
Hälsen varandra med en helig kyss.
Alla de heliga hälsa eder.
Herrens, Jesu Kristi, nåd och Guds kärlek och den helige Andes delaktighet vare med eder alla.
Paulus, apostel, icke från människor, ej heller genom någon människa, utan genom Jesus Kristus och genom Gud, Fadern, som har uppväckt honom från de döda --
jag, jämte alla de bröder som äro här med mig, hälsar församlingarna i Galatien.
Nåd vare med eder och frid ifrån Gud, vår Fader, och ifrån Herren Jesus Kristus,
som har utgivit sig själv för våra synder, för att rädda oss från den nuvarande onda tidsåldern, efter vår Guds och Faders vilja.
Honom tillhör äran i evigheternas evigheter.
Amen.
Det förundrar mig att I så hastigt avfallen från honom, som har kallat eder till att vara i Kristi nåd, och vänden eder till ett nytt evangelium.
Likväl är detta icke något annat »evangelium»; det är allenast så, att några finnas som vålla förvirring bland eder och vilja förvända Kristi evangelium.
Men om någon, vore det ock vi själva eller en ängel från himmelen, förkunnar evangelium i strid mot vad vi hava förkunnat för eder, så vare han förbannad.
Ja, såsom vi förut hava sagt, så säger jag nu åter: Om någon förkunnar evangelium för eder i strid mot vad I haven undfått, så vare han förbannad.
Är det då människor som jag nu söker vinna för mig, eller är det Gud?
Står jag verkligen efter att »vara människor till behag»?
Nej, om jag ännu ville vara människor till behag, så vore jag icke en Kristi tjänare.
Ty det vill jag säga eder, mina bröder, att det evangelium som har blivit förkunnat av mig icke är någon människolära.
Det är ju icke heller av någon människa som jag har undfått det eller blivit undervisad däri, utan genom en uppenbarelse från Jesus Kristus.
I haven ju hört huru det var med mig, medan jag ännu vandrade i judiskt väsende: att jag då övermåttan våldsamt förföljde Guds församling och ville utrota den,
ja, att jag gick längre i judiskt väsende än många av mina samtida landsmän och ännu ivrigare nitälskade för mina fäders stadgar.
Men när han, som allt ifrån min moders liv har avskilt mig, och som genom sin nåd har kallat mig,
täcktes i mig uppenbara sin Son, för att jag bland hedningarna skulle förkunna evangelium om honom, då begav jag mig strax åstad; jag rådförde mig icke med någon människa,
ej heller for jag upp till Jerusalem, till dem som före mig voro apostlar.
I stället for jag bort till Arabien och vände så åter tillbaka till Damaskus.
Först sedan, tre år därefter, for jag upp till Jerusalem, för att lära känna Cefas, och jag stannade hos honom femton dagar.
Men av de andra apostlarna såg jag ingen; allenast Jakob, Herrens broder, såg jag.
Och Gud vet att jag icke ljuger i vad jag här skriver till eder.
Därefter for jag till Syriens och Ciliciens bygder.
Men för de kristna församlingarna i Judeen var jag personligen okänd.
De hörde allenast huru man sade: »Han som förut förföljde oss, han förkunnar nu evangelium om den tro som han förr ville utrota.»
Och de prisade Gud för min skull.
Efter fjorton års förlopp for jag sedan åter upp till Jerusalem, åtföljd av Barnabas; jag tog då också Titus med mig.
Men det var på grund av en uppenbarelse som jag for dit.
Och för bröderna där framlade jag det evangelium som jag predikar bland hedningarna; särskilt framlade jag det för de män som stodo högst i anseende -- detta av oro för att mitt strävande nu vore förgäves eller förut hade varit det.
Men icke ens Titus, min följeslagare, som var grek, blev nödgad att låta omskära sig.
Det var nämligen så, att några falska bröder hade kommit att upptagas i församlingen, dit de hade smugit sig in för att bespeja vår frihet, den som vi hava i Kristus Jesus, varefter de ville trälbinda oss.
Dock gåvo vi icke ens ett ögonblick vika för dem genom en sådan underkastelse; ty vi ville att evangelii sanning skulle bliva bevarad hos eder.
Och vad angår dem som ansågos något vara -- hurudana de nu voro, det kommer icke mig vid; Gud har icke anseende till personen -- så sökte icke dessa män, de som stodo högst i anseende, att pålägga mig några nya förpliktelser.
Tvärtom; de sågo att jag hade blivit betrodd med att förkunna evangelium för de oomskurna, likasom Petrus hade fått de omskurna på sin del --
ty densamme som hade stått Petrus bi vid hans apostlaverksamhet bland de omskurna, han hade ock stått mig bi bland hedningarna --
och när de nu förnummo vilken nåd som hade blivit mig given, räckte de mig och Barnabas handen till samarbete, både Jakob och Cefas och Johannes, de män som räknades för själva stödjepelarna; vi skulle verka bland hedningarna, och de bland de omskurna.
Allenast skulle vi tänka på de fattiga; och just detta har jag också vinnlagt mig om att göra.
Men när Cefas kom till Antiokia, trädde jag öppet upp mot honom, ty han hade befunnits skyldig till en försyndelse.
Förut hade han nämligen ätit tillsammans med hedningarna; men så kommo några män dit från Jakob, och efter deras ankomst drog han sig tillbaka och höll sig undan, av fruktan för de omskurna.
Till samma skrymteri gjorde sig också de andra judarna skyldiga, och så blev till och med Barnabas indragen i deras skrymteri.
Men när jag såg att de icke vandrade med fasta steg, enligt evangelii sanning, sade jag till Cefas i allas närvaro: »Om du, som är en jude, kan leva efter hednisk sed i stället för efter judisk, varför vill du då nödga hedningarna att leva efter judiskt sätt?»
Vi för vår del äro väl på grund av vår härkomst judar och icke »hedniska syndare»;
men då vi nu veta att en människa icke bliver rättfärdig av laggärningar, utan genom tro på Kristus Jesus, hava också vi satt vår tro till Jesus Kristus, för att vi skola bliva rättfärdiga av tro på Kristus, och icke av laggärningar.
Ty av laggärningar bliver intet kött rättfärdigt.
Men om nu jämväl vi, i det vi sökte att bliva rättfärdiga i Kristus, hava befunnits vara syndare, då är ju Kristus en syndatjänare?
Bort det!
Om så vore att jag byggde upp igen detta samma som jag redan har brutit ned, då bevisade jag därmed, att jag var en överträdare.
Ty jag för min del har genom lagen dött bort ifrån lagen, för att jag skall leva för Gud.
Jag är korsfäst med Kristus,
och nu lever icke mer jag, utan Kristus lever i mig; och det liv som jag nu lever i köttet, det lever jag i tron på Guds Son, som har älskat mig och utgivit sig själv för mig.
Jag förkastar icke Guds nåd.
Om rättfärdighet kunde vinnas genom lagen, då hade ju Kristus icke behövt lida döden.
I oförståndige galater!
Vem har så dårat eder, I som dock haven fått Jesus Kristus målad för edra ögon såsom korsfäst?
Allenast det vill jag att I skolen svara mig på: Kom det sig av laggärningar att I undfingen Anden, eller kom det sig därav att I lyssnaden i tro?
Ären I så oförståndiga?
I, som haven begynt i Anden, viljen I nu sluta i köttet?
Haven I då upplevat så mycket förgäves -- om det nu verkligen har varit förgäves?
Alltså, att han som förlänade eder Anden och utförde kraftgärningar bland eder gjorde detta, kom det sig av laggärningar eller därav att I lyssnaden i tro,
i enlighet med det ordet: »Abraham trodde Gud, och det räknades honom till rättfärdighet»?
Så mån I nu veta att de som låta det bero på tro, de äro Abrahams barn.
Och eftersom skriften förutsåg att det var av tro som hedningarna skulle bliva rättfärdiggjorda av Gud, så gav den i förväg åt Abraham detta glada budskap: »I dig skola alla folk varda välsignade.»
Alltså bliva de som låta det bero på tro välsignade tillika med Abraham, honom som trodde.
Ty alla de som låta det bero på laggärningar, de äro under förbannelse.
Det är nämligen skrivet: »Förbannad vare var och en som icke förbliver vid allt som är skrivet i lagens bok, och icke gör därefter.»
Och att ingen i kraft av lag bliver rättfärdig inför Gud, det är uppenbart, eftersom det heter: »Den rättfärdige skall leva av tro.»
Men i lagen beror det icke på tro; tvärtom heter det: »Den som gör efter dessa stadgar skall leva genom dem.»
Kristus friköpte oss från lagens förbannelse, när han blev en förbannelse för vår skull.
Det är ju skrivet: »Förbannad är var och en som är upphängd på trä.»
Vi friköptes, för att den välsignelse som hade givits åt Abraham skulle i Jesus Kristus komma också hedningarna till del, så att vi genom tron skulle undfå den utlovade Anden.
Mina bröder, jag vill taga ett exempel från vad som gäller bland människor.
Icke ens när fråga är om en människas testamentsförordnande, kan någon upphäva det eller lägga något därtill, sedan det en gång har vunnit gällande kraft.
Nu gåvos löftena åt Abraham, så ock åt hans »säd».
Det heter icke: »och åt dem som komma av din säd», såsom när det talas om många; utan det heter, såsom när det talas om en enda: »och åt din säd», vilken är Kristus.
Vad jag alltså vill säga är detta: Ett förordnande som Gud redan hade givit gällande kraft kan icke genom en lag, som utgavs fyra hundra trettio år därefter, hava blivit ogiltigt, så att löftet därmed har gjorts om intet.
Om det nämligen vore på grund av lag som arvet skulle undfås, så vore det icke på grund av löfte.
Men åt Abraham har Gud skänkt det genom ett löfte.
Vartill tjänade då lagen?
Jo, på det att överträdelserna skulle komma i dagen, blev den efteråt given, för att gälla till dess att »säden» skulle komma, han åt vilken löftet hade blivit givet; och den utgavs genom änglar och överlämnades i en medlares hand.
Men den som är medlare är icke medlare för allenast en enda.
Men Gud är en.
Är då lagen emot Guds löften?
Bort det!
Om en lag hade blivit given, som kunde göra levande, då skulle rättfärdigheten verkligen komma av lagen.
Men nu har skriften inneslutit alltsammans under synd, för att det som var utlovat skulle, av tro på Jesus Kristus, komma dem till del som tro.
Men förrän tron kom, voro vi inneslutna under lagen och höllos i förvar under den, i förbidan på den tro som en gång skulle uppenbaras.
Så har lagen blivit vår uppfostrare till Kristus, för att vi skola bliva rättfärdiga av tro.
Men sedan tron har kommit, stå vi icke mer under uppfostrare.
Alla ären I Guds barn genom tron, i Kristus Jesus;
ty I alla, som haven blivit döpta till Kristus, haven iklätt eder Kristus.
Här är icke jude eller grek, här är icke träl eller fri, här är icke man och kvinna: alla ären I ett i Kristus Jesus.
Hören I nu Kristus till, så ären I därmed ock Abrahams säd, arvingar enligt löftet.
Vad jag vill säga är detta: Så länge arvingen är barn, finnes ingen skillnad mellan honom och en träl, fastän han är herre över alla ägodelarna;
ty han står under förmyndare och förvaltare, intill den tid som fadern har bestämt.
Sammalunda höllos ock vi, när vi voro barn, i träldom under världens »makter».
Men när tiden var fullbordad, sände Gud sin Son, född av kvinna och ställd under lagen,
för att han skulle friköpa dem som stodo under lagen, så att vi skulle få söners rätt.
Och eftersom I nu ären söner, har han sänt i våra hjärtan sin Sons Ande, som ropar: »Abba!
Fader!»
Så är du nu icke mer träl, utan son; och är du son, så är du ock arvinge, insatt därtill av Gud.
Förut, innan I ännu känden Gud, voren I trälar under gudar som till sitt väsende icke voro gudar.
Men nu, sedan I haven lärt känna Gud och, vad mer är, haven blivit kända av Gud, huru kunnen I nu vända tillbaka till de svaga och arma »makter», under vilka I åter på nytt viljen bliva trälar?
I akten ju på dagar och på månader och på särskilda tider och år. --
Jag är bekymrad för eder och fruktar att jag till äventyrs har arbetat förgäves för eder.
Jag beder eder, mina bröder: Bliven såsom jag är, eftersom jag har blivit såsom I voren.
I haven icke gjort mig något för när.
I veten ju att det var på grund av kroppslig svaghet som jag första gången kom att förkunna evangelium för eder.
Och fastän mitt kroppsliga tillstånd då väl hade kunnat innebära en frestelse för eder, så sågen I det ändå icke med ringaktning eller leda, utan togen emot mig såsom en Guds ängel, ja, såsom Kristus Jesus själv.
När hör man eder nu prisa eder saliga?
Det vittnesbördet kan jag nämligen giva eder, att I då, om så hade varit möjligt, skullen hava rivit ut edra ögon och givit dem åt mig.
Så har jag då blivit eder ovän därigenom att jag säger eder sanningen!
Man söker med iver att vinna eder för sig, men icke med en god iver; nej, del vilja avspärra eder från andra, för att I med så mycket större iver skolen hålla eder till dem.
Och det är nu gott att I bliven omfattade med ivrig omsorg, i en god sak, alltid, och icke allenast när jag är tillstädes hos eder,
I mina barn, som jag nu åter med vånda måste föda till livet, intill dess att Kristus har tagit gestalt i eder.
Jag skulle önska att jag just nu vore hos eder och kunde göra min röst rätt bevekande.
Ty jag vet mig knappt någon råd med eder.
Sägen mig, I som viljen stå under lagen: haven I icke hört vad lagen säger?
Det är ju skrivet att Abraham fick två söner, en med sin tjänstekvinna, och en med sin fria hustru.
Men tjänstekvinnans son är född efter köttet, då däremot den fria hustruns son är född i kraft av löftet.
Dessa ord hava en djupare mening; ty de båda kvinnorna beteckna två förbund.
Av dessa kommer det ena från berget Sina och föder sina barn till träldom, och detta har sin förebild i Agar.
Berget Sina kallas nämligen i Arabien för Agar och svarar emot det nuvarande Jerusalem, ty detta lever med sina barn i träldom.
Men det Jerusalem som är därovan, det är fritt, och det är vår moder.
Så är ju skrivet: »Jubla, du ofruktsamma, du som icke föder barn; brist ut och ropa, du som icke bliver moder, Ty den ensamma skall hava många barn, flera än den som har man.»
Och I, mina bröder, ären löftets barn, likasom Isak var.
Men likasom förr i tiden den son som var född efter köttet förföljde den som var född efter Anden, så är det ock nu.
Dock, vad säger skriften? »Driv ut tjänstekvinnan och hennes son; ty tjänstekvinnans son skall förvisso icke ärva med den fria hustruns son.»
Alltså, mina bröder, vi äro icke barn av en tjänstekvinna, utan av den fria hustrun.
För att vi skola vara fria, har Kristus frigjort oss.
Stån därför fasta, och låten icke något nytt träldomsok läggas på eder.
Se, jag säger eder, jag Paulus, att om I låten omskära eder, så bliver Kristus eder till intet gagn.
Och för var och en som låter omskära sig betygar jag nu åter att han är pliktig att fullgöra hela lagen.
I haven kommit bort ifrån Kristus, I som viljen bliva rättfärdiga i kraft av lagen; I haven fallit ur nåden.
Vi vänta nämligen genom ande, av tro, den rättfärdighet som är vårt hopp.
Ty i Kristus Jesus betyder det intet huruvida någon är omskuren eller oomskuren; allt beror på huruvida han har en tro som är verksam genom kärlek.
I begynten edert lopp väl.
Vem har nu lagt hinder i eder väg, så att I icke mer lyden sanningen?
Till sådant kom ingen maning från honom som har kallat eder.
Litet surdeg syrar hela degen.
För min del har jag i Herren den tillförsikten till eder, att I icke häri skolen tänka på annat sätt; men den som vållar förvirring bland eder, han skall bära sin dom, vem han än må vara.
Om så vore, mina bröder, att jag själv ännu predikade omskärelse, varför skulle jag då ännu alltjämt lida förföljelse?
Då vore ju korsets stötesten röjd ur vägen. --
Jag skulle önska att de män som uppvigla eder läte omskära sig ända till avstympning.
I ären ju kallade till frihet, mina bröder; bruken dock icke friheten så, att köttet får något tillfälle.
Fastmer mån I tjäna varandra genom kärleken.
Ty hela lagens uppfyllelse ligger i ett enda budord, nämligen detta: »Du skall älska din nästa såsom dig själv.»
Men om I bitens inbördes och äten på varandra, så mån I se till, att I icke bliven uppätna av varandra.
Vad jag vill säga är detta: Vandren i ande, så skolen I förvisso icke göra vad köttet har begärelse till.
Ty köttet har begärelse mot Anden, och Anden mot köttet; de två ligga ju i strid med varandra, för att hindra eder att göra vad I viljen.
Men om I drivens av ande, så stån I icke under lagen.
Men köttets gärningar äro uppenbara: de äro otukt, orenhet, lösaktighet,
avgudadyrkan, trolldom, ovänskap, kiv, avund, vrede, genstridighet, tvedräkt, partisöndring,
missunnsamhet, mord, dryckenskap, vilt leverne och annat sådant, varom jag säger eder i förväg, såsom jag redan förut har sagt, att de som göra sådant, de skola icke få Guds rike till arvedel.
Andens frukt åter är kärlek, glädje, frid, tålamod, mildhet, godhet, trofasthet,
saktmod, återhållsamhet.
Mot sådant är icke lagen.
Och de som höra Kristus Jesus till hava korsfäst sitt kött tillika med dess lustar och begärelser.
Om vi nu hava liv genom ande, så låtom oss ock vandra i ande.
Låtom oss icke söka fåfänglig ära, i det att vi utmana varandra och avundas varandra.
Mina bröder, om så händer att någon ertappas med att begå en försyndelse, då mån I, som ären andliga människor, upprätta honom i saktmods ande.
Och du må hava akt på dig själv, att icke också du bliver frestad.
Bären varandras bördor; så uppfyllen I Kristi lag.
Ty om någon tycker sig något vara, fastän han intet är, så bedrager han sig själv.
Må var och en pröva sina egna gärningar; han skall då tillmäta sig berömmelse allenast efter vad han själv är, och icke efter vad andra äro.
Ty var och en har sin egen börda att bära.
Den som får undervisning i ordet, han låte den som undervisar honom få del med sig i allt gott.
Faren icke vilse.
Gud låter icke gäcka sig.
Ty vad människan sår, det skall hon ock skörda.
Den som sår i sitt kötts åker, han skall av köttet skörda förgängelse, men den som sår i Andens åker, han skall av Anden skörda evigt liv.
Och låtom oss icke förtröttas att göra vad gott är; ty om vi icke uppgivas, så skola vi, när tiden är inne, få inbärga vår skörd.
Må vi alltså, medan vi hava tillfälle, göra vad gott är mot var man, och först och främst mot dem som äro våra medbröder i tron.
Sen här med vilka stora bokstäver jag egenhändigt skriver till eder!
Alla de som eftersträva ett gott anseende här i köttet, de vilja nödga eder till omskärelse, detta allenast för att de själva skola undgå att bliva förföljda för Kristi kors' skull.
Ty icke ens dessa omskurna själva hålla lagen.
Nej, det är för att kunna berömma sig av edert kött som de vilja att I skolen låta omskära eder.
Men vad mig angår, så vare det fjärran ifrån mig att berömma mig av något annat än av vår Herres, Jesu Kristi, kors, genom vilket världen för mig är korsfäst, och jag för världen.
Ty det kommer icke an på om någon är omskuren eller oomskuren; allt beror på huruvida han är en ny skapelse.
Och över alla dem som komma att vandra efter detta rättesnöre, över dem vare frid och barmhärtighet, ja, över Guds Israel.
Må nu ingen härefter vålla mig oro; ty jag bär Jesu märken på min kropp.
Vår Herres, Jesu Kristi, nåd vare med eder ande, mina bröder.
Amen.
Paulus, genom Guds vilja Kristi Jesu apostel, hälsar de heliga som bo i Efesus, de i Kristus Jesus troende.
Nåd vare med eder och frid ifrån Gud, vår Fader, och Herren Jesus Kristus.
Välsignad vare vår Herres, Jesu Kristi, Gud och Fader, som i Kristus har välsignat oss med all den himmelska världens andliga välsignelse,
såsom han ju, förrän världens grund var lagd, har utvalt oss i honom till att vara heliga och ostraffliga inför sig.
Ty i sin kärlek förutbestämde han oss till barnaskap hos sig, genom Jesus Kristus, efter sin viljas behag,
den nådeshärlighet till pris, varmed han har benådat oss i den älskade.
I honom hava vi förlossning genom hans blod, förlåtelse för våra synder, efter hans nåds rikedom.
Och denna nåd har han i överflödande mått låtit komma oss till del, med all vishet och allt förstånd,
i det att han för oss har kungjort sin viljas hemlighet, enligt det beslut som han efter sitt behag hade fattat inom sig själv,
om en ordning som i tidernas fullbordan skulle komma till stånd, det beslutet att i Kristus sammanfatta allt som finnes i himmelen och på jorden.
I honom hava vi ock undfått vår arvslott, vi som förut voro bestämda därtill genom dens beslut, som verkar allting efter sin egen viljas råd.
Så skulle vi, hans härlighet till pris, vara de som i Kristus redan i förväg hava ägt ett hopp.
I honom haven jämväl I, sedan I haven fått höra sanningens ord, eder frälsnings evangelium, ja, i honom haven I, sedan I nu ock haven kommit till tron, såsom ett insegel undfått den utlovade helige Ande,
vilken är en underpant på vårt arv, till förvissning om att hans egendomsfolk skall förlossas, hans härlighet till pris.
Sedan jag fick höra om eder tro i Herren Jesus och om eder kärlek till alla de heliga,
har därför jag å min sida icke upphört att tacka Gud för eder, när jag tänker på eder i mina böner.
Och min bön är att vår Herres, Jesu Kristi, Gud, härlighetens Fader, må giva eder en visdomens och uppenbarelsens ande till kunskap om sig,
och att han må upplysa edra hjärtans ögon, så att I förstån hurudant det hopp är, vartill han har kallat eder, huru rikt på härlighet hans arv är bland de heliga,
och huru översvinnligt stor hans makt är på oss som tro -- allt i enlighet med den väldiga styrkas kraft,
varmed han har verkat i Kristus, i det att han uppväckte honom från de döda och satte honom på sin högra sida i den himmelska världen,
över alla andevärldens furstar och väldigheter och makter och herrar, ja, över allt som kan nämnas, icke allenast i denna tidsålder, utan ock i den tillkommande.
»Allt lade han under hans fötter.»
Och honom gav han åt församlingen till att vara ett huvud över allting --
åt församlingen, ty den är hans kropp och är uppfylld av honom som uppfyller allt i alla.
Så har han ock gjort eder levande, eder som voren döda genom de överträdelser och synder
i vilka I förut vandraden, efter denna världs och tidsålders sätt, i det I följden fursten över luftens härsmakt, över den andemakt som nu är verksam i de ohörsamma.
Bland dessa voro förut också vi allasammans, där vi vandrade i vårt kötts begärelser och gjorde vad köttet och sinnet ville; och vi voro genom vår natur hemfallna åt vredesdomen, vi likasom de andra.
Men Gud, som är rik på barmhärtighet, har, för den stora kärleks skull, varmed han har älskat oss,
gjort oss levande med Kristus, oss som voro döda genom våra synder.
Av nåd ären I frälsta!
Ja, han har uppväckt oss med honom och satt oss med honom i den himmelska världen, i Kristus Jesus,
för att i de kommande tidsåldrarna bevisa sin nåds översvinnliga rikedom, genom godhet mot oss i Kristus Jesus.
Ty av nåden ären I frälsta genom tro -- och det icke av eder själva, Guds gåva är det --
icke av gärningar, för att ingen skall berömma sig.
Ty hans verk äro vi, skapade i Kristus Jesus till goda gärningar, vilka Gud förut har berett, för att vi skola vandra i dem.
Kommen därför ihåg att I förut, I som voren hedningar i köttet och bleven kallade oomskurna av dem som kallas omskurna, efter den omskärelse som med händer göres på köttet --
kommen ihåg att I på den tiden, då när I voren utan Kristus, voren utestängda från medborgarskap i Israel och främmande för löftets förbund, utan hopp och utan Gud i världen.
Nu däremot, då I ären i Kristus Jesus, haven I, som förut voren fjärran, kommit nära, i och genom Kristi blod.
Ty han är vår frid, han som av de båda har gjort ett och brutit ned den skiljemur som stod emellan oss, nämligen ovänskapen.
Ty i sitt kött gjorde han om intet budens stadgelag, för att han skulle av de två i sig skapa en enda ny människa och så bereda frid,
och för att han skulle åt dem båda, förenade i en enda kropp, skaffa försoning med Gud, sedan han genom korset hade i sin person dödat ovänskapen.
Och han har kommit och har förkunnat det glada budskapet om frid för eder, I som voren fjärran, och om frid för dem som voro nära.
Ty genom honom hava vi, de ena såväl som de andra, i en och samme Ande tillträde till Fadern.
Alltså ären I nu icke mer främlingar och gäster, utan I haven medborgarskap med de heliga och ären Guds husfolk,
uppbyggda på apostlarnas och profeternas grundval, där hörnstenen är Kristus Jesus själv,
i vilken allt det som uppbygges bliver sammanslutet och så växer upp till ett heligt tempel i Herren.
I honom bliven också I med de andra uppbyggda till en Guds boning, i Anden.
Fördenskull böjer jag mina knän, jag Paulus, som till gagn för eder, I hedningar, är Kristi Jesu fånge.
I haven väl hört om det nådesuppdrag av Gud, som är mig givet för eder räkning,
huru genom uppenbarelse den hemlighet blev för mig kungjord, varom jag ovan har i korthet skrivit.
Och när I läsen detta, kunnen I därav förstå vilken insikt jag har i Kristi hemlighet,
som under förgångna släktens tider icke hade blivit kungjord för människors barn, såsom den nu genom andeingivelse har blivit uppenbarad för hans heliga apostlar och profeter.
Jag menar den hemligheten, att hedningarna i Kristus Jesus äro våra medarvingar och jämte oss lemmar i en och samma kropp och jämte oss delaktiga i löftet -- detta genom evangelium,
vars tjänare jag har blivit i följd av den Guds nåds gåva som blev mig given genom hans mäktiga kraft.
Ja, åt mig, den ringaste bland alla heliga, blev den nåden given att för hedningarna förkunna evangelium om Kristi outrannsakliga rikedom,
och att lägga i dagen huru det rådslut har blivit utfört, som tidsåldrarna igenom hade såsom en hemlighet varit fördolt i Gud, alltings skapare.
Ty Gud ville att hans mångfaldiga visdom nu, i och genom församlingen, skulle bliva kunnig för furstarna och väldigheterna i den himmelska världen.
Sådant hade hans beslut varit från tidsåldrarnas begynnelse, det som han utförde i Kristus Jesus, vår Herre.
Och i honom kunna vi med tillförsikt frimodigt träda fram, genom tron på honom.
Därför beder jag eder att icke fälla modet vid mina lidanden för eder; de lända ju eder till ära.
Fördenskull böjer jag mina knän för Fadern --
honom från vilken allt vad fader heter i himmelen och på jorden har sitt namn --
och beder att han ville efter sin härlighets rikedom förläna eder, att I genom hans Ande växen till i kraft till eder invärtes människa,
och att Kristus genom tron må bo i edra hjärtan, och att I mån vara rotade och grundade i kärleken,
så att I, tillika med alla de heliga, till fullo förmån fatta vad bredden och längden och höjden och djupet är
och så lära känna Kristi kärlek, som övergår all kunskap.
Ty så skolen I bliva helt uppfyllda av all Guds fullhet.
Men honom, som förmår göra mer, ja, långt mer än allt vad vi bedja eller tänka, efter den kraft som är verksam i oss,
honom tillhör äran i församlingen och i Kristus Jesus alla släkten igenom i evigheternas evighet, amen.
Så förmanar jag nu eder, jag som är en fånge i Herren, att föra en vandel som är värdig den kallelse I haven undfått,
med all ödmjukhet och allt saktmod, med tålamod, så att I haven fördrag med varandra i kärlek
och vinnläggen eder om att bevara Andens enhet genom fridens band:
en kropp och en Ande, likasom I ock bleven kallade till att leva i ett och samma hopp, det som tillhör eder kallelse --
en Herre, en tro, ett dop, en Gud, som är allas Fader,
han som är över alla, genom alla och i alla.
Men åt var och en särskild av oss blev nåden given, alltefter som Kristus tillmätte honom sin gåva.
Därför heter det: »Han for upp i höjden, han tog fångar, han gav människorna gåvor.»
Men detta ord »han for upp», vad innebär det, om icke att han förut hade farit hit ned till jordens lägre rymder?
Den som for ned, han är ock den som for upp över alla himlar, för att han skulle uppfylla allt.
Och han gav oss somliga till apostlar, somliga till profeter, somliga till evangelister, somliga till herdar och lärare.
Ty han ville göra de heliga skickliga till att utföra sitt tjänarvärv, att uppbygga Kristi kropp,
till dess att vi allasammans komma fram till enheten i tron och i kunskapen om Guds Son, till manlig mognad, och så bliva fullvuxna, intill Kristi fullhet.
Så skulle vi icke mer vara barn, icke såsom havets vågor drivas omkring av vart vindkast i läran, vid människornas bedrägliga spel, när de illfundigt söka främja villfarelsens listiga anslag.
Nej, vi skulle då hålla oss till sanningen, och i alla stycken i kärlek växa upp till honom som är huvudet, Kristus.
Ty från honom hämtar hela kroppen sin tillväxt, till att bliva uppbyggd i kärlek, i det att den sammanslutes och får sammanhållning genom det bistånd var led giver, med en kraft som är avmätt efter var särskild dels uppgift.
Jag tillsäger eder alltså och uppmanar eder allvarligt i Herren, att icke mer vandra såsom hedningarna i sitt sinnes fåfänglighet vandra,
hedningarna, vilka, i följd av den okunnighet som råder hos dem genom deras hjärtans förstockelse, äro förmörkade till förståndet och bortkomna från det liv som är av Gud.
Ty i sin försoffning hava de överlämnat sig åt lösaktighet, så att de i girighet bedriva alla slags orena gärningar.
Men I haven icke fått en sådan undervisning om Kristus,
om I eljest så haven hört om honom och så blivit lärda i honom, som sanning är i Jesus:
att I -- då detta nu krävdes på grund av eder förra vandel -- haven avlagt den gamla människan, som fördärvar sig genom att följa sina begärelsers bedrägliga lockelser,
och nu förnyens genom Anden som bor i edert sinne,
och att I haven iklätt eder den nya människan, som är skapad till likhet med Gud i sanningens rättfärdighet och helighet.
Läggen därför bort lögnen, och talen sanning med varandra, eftersom vi äro varandras lemmar.
»Vredgens, men synden icke»; låten icke solen gå ned över eder vrede,
och given icke djävulen något tillfälle.
Den som har stulit, han stjäle icke mer, utan arbete hellre, och uträtte med sina händer vad gott är, så att han har något varav han kan dela med sig åt den som lider brist.
Låten intet ohöviskt tal utgå ur eder mun, utan allenast det som är gott, till uppbyggelse, där sådan behöves, så att det bliver till välsignelse för dem som höra det.
Och bedröven icke Guds helige Ande, vilken I haven undfått såsom ett insegel, för förlossningens dag.
All bitterhet och häftighet och vrede, allt skriande och smädande, ja, allt vad ondska heter vare fjärran ifrån eder.
Varen i stället goda och barmhärtiga mot varandra, och förlåten varandra, såsom Gud i Kristus har förlåtit eder.
Bliven alltså Guds efterföljare, såsom hans älskade barn,
och vandren i kärlek, såsom Kristus älskade eder och utgav sig själv för oss till en gåva och ett offer, »Gud till en välbehaglig lukt».
Men otukt och orenhet, av vad slag det vara må, och girighet skolen I, såsom det anstår heliga, icke ens låta nämnas bland eder,
ej heller ohöviskt väsende och dåraktigt tal och gyckel; sådant är otillbörligt.
Låten fastmer tacksägelse höras.
Ty det bören I veta, och det insen I också själva, att ingen otuktig eller oren människa har arvedel i Kristi och Guds rike, ej heller någon girig, ty en sådan är en avgudadyrkare.
Låten ingen bedraga eder med tomma ord; ty för sådana synder kommer Guds vrede över de ohörsamma.
Haven alltså ingen del i sådant.
I voren ju förut mörker, men nu ären I ljus i Herren; vandren då såsom ljusets barn.
Ty ljusets frukt består i allt vad godhet och rättfärdighet och sanning är.
Ja, vandren så, i det att I pröven vad som är välbehagligt för Herren.
Och haven ingen delaktighet i mörkrets gärningar, som icke giva någon frukt, utan avslöjen dem fastmer.
Vad av sådana människor i hemlighet förövas, därom är det skamligt till och med att tala;
men alltsammans bliver uppenbart, när det avslöjas genom ljuset.
Ty varhelst något bliver uppenbart, där är ljus.
Därför heter det: »Vakna upp, du som sover, och stå upp ifrån de döda, så skall Kristus lysa fram för dig.»
Sen därför noga till, huru I vandren: att I vandren icke såsom ovisa människor, utan såsom visa;
och tagen väl i akt vart lägligt tillfälle.
Ty tiden är ond.
Varen alltså icke oförståndiga, utan förstån vad som är Herrens vilja.
Och dricken eder icke druckna av vin; ty därav kommer ett oskickligt leverne.
Låten eder fastmer uppfyllas av ande,
och talen till varandra i psalmer och lovsånger och andliga visor, och sjungen och spelen till Herrens ära i edra hjärtan,
och tacken alltid Gud och Fadern för allt, i vår Herres, Jesu Kristi, namn.
Underordnen eder varandra i Kristi fruktan.
I hustrur, underordnen eder edra män, såsom I underordnen eder Herren;
ty en man är sin hustrus huvud, såsom Kristus är församlingens huvud, han som ock är denna sin kropps Frälsare.
Ja, såsom församlingen underordnar sig Kristus, så skola ock hustrurna i allt underordna sig sina män.
I män, älsken edra hustrur, såsom Kristus har älskat församlingen och utgivit sig själv för henne
till att helga henne, genom att rena henne medelst vattnets bad, i kraft av ordet.
Ty så ville han själv ställa fram församlingen inför sig i härlighet, utan fläck och skrynka och annat sådant; fastmer skulle hon vara helig och ostrafflig.
På samma sätt äro männen pliktiga att älska sina hustrur, då dessa ju äro deras egna kroppar; den som älskar sin hustru, han älskar sig själv.
Ingen har någonsin hatat sitt eget kött; i stället när och omhuldar man det, såsom Kristus gör med församlingen,
eftersom vi äro lemmar av hans kropp.
»Fördenskull skall en man övergiva sin fader och sin moder och hålla sig till sin hustru, och de tu skola varda ett kött.» --
Den hemlighet som ligger häri är stor; jag säger detta med tanke på Kristus och församlingen.
Dock gäller också om eder att var och en skall älska sin hustru såsom sig själv; men hustrun å sin sida skall visa sin man vördnad.
I barn, varen edra föräldrar lydiga i Herren, ty detta är rätt och tillbörligt.
»Hedra din fader och din moder.»
Det är ju först detta bud som har ett löfte med sig:
»för att det må gå dig väl och du må länge leva på jorden».
Och I fäder, reten icke edra barn till vrede, utan fostren dem i Herrens tukt och förmaning.
I tjänare, varen edra jordiska herrar lydiga, med fruktan och bävan, av uppriktigt hjärta, såsom gällde det Kristus;
icke med ögontjänst, av begär att behaga människor, utan såsom Kristi tjänare, som av hjärtat göra Guds vilja;
och gören eder tjänst med villighet, såsom tjänaden I Herren och icke människor.
I veten ju att vad gott var och en gör, det skall han få igen av Herren, vare sig han är träl eller fri.
Och I herrar, handlen på samma sätt mot dem, och upphören att bruka hårda ord; I veten ju att i himmelen finnes den som är Herre över både dem och eder, och att hos honom icke finnes anseende till personen.
För övrigt, bliven allt starkare i Herren och i hans väldiga kraft.
Ikläden eder hela Guds vapenrustning, så att I kunnen hålla stånd emot djävulens listiga angrepp.
Ty den kamp vi hava att utkämpa är en kamp icke mot kött och blod, utan mot furstar och väldigheter och världshärskare, som råda här i mörkret, mot ondskans andemakter i himlarymderna.
Tagen alltså på eder hela Guds vapenrustning, så att I kunnen stå emot på den onda dagen och, sedan I haven fullgjort allt, behålla fältet.
Stån därför omgjordade kring edra länder med sanningen, och »varen iklädda rättfärdighetens pansar»,
och haven såsom skor på edra fötter den beredvillighet som fridens evangelium giver.
Och tagen alltid trons sköld, varmed I skolen kunna utsläcka den ondes alla brinnande pilar.
Och låten giva eder »frälsningens hjälm» och Andens svärd, som är Guds ord.
Gören detta under ständig åkallan och bön, så att I alltjämt bedjen i Anden och fördenskull vaken, under ständig uthållighet och ständig bön för alla de heliga.
Bedjen ock för mig, att min mun må upplåtas, och att det jag skall tala må bliva mig givet, så att jag frimodigt kungör evangelii hemlighet,
för vars skull jag är ett sändebud i kedjor; ja, bedjen att jag må frimodigt tala därom med de rätta orden.
Men för att ock I skolen få veta något om mig, huru det går mig, kommer Tykikus, min älskade broder och trogne tjänare i Herren, att underrätta eder om allt.
Honom sänder jag till eder, just för att I skolen få veta huru det är med oss, och för att han skall hugna edra hjärtan.
Frid vare med bröderna och kärlek tillika med tro, från Gud, Fadern, och Herren Jesus Kristus.
Nåd vare med alla som älska vår Herre Jesus Kristus -- nåd i oförgängligt liv.
Paulus och Timoteus, Kristi Jesu tjänare, hälsa alla de heliga i Kristus Jesus som bo i Filippi, tillika med församlingsföreståndare och församlingstjänare.
Nåd vare med eder och frid ifrån Gud, vår Fader, och Herren Jesus Kristus.
Jag tackar min Gud, så ofta jag tänker på eder,
i det jag alltid i alla mina böner med glädje beder för eder alla.
Jag tackar honom för att I, allt ifrån första dagen intill nu, haven deltagit i arbetet för evangelium.
Och jag har den tillförsikten, att han som i eder har begynt ett gott verk, han skall ock fullborda det, intill Kristi Jesu dag.
Och det är ju rätt och tillbörligt att jag tänker så om eder alla, eftersom jag, både när jag ligger i bojor, och när jag försvarar och befäster evangelium, har eder i mitt hjärta såsom alla med mig delaktiga i nåden.
Ty Gud är mitt vittne, han vet huru jag längtar efter eder alla med Kristi Jesu kärlek.
Och därom beder jag, att eder kärlek må allt mer och mer överflöda av kunskap och förstånd i allt,
så att I kunnen döma om vad rättast är, på det att I mån bliva rena och för ingen till stötesten, i väntan på Kristi dag,
och bliva rika på rättfärdighetens frukt, vilken kommer genom Jesus Kristus, Gud till ära och pris.
Jag vill att I, mina bröder, skolen veta att det som har vederfarits mig snarare har länt till evangelii framgång.
Det har nämligen så blivit uppenbart för alla i pretoriet och för alla andra, att det är i Kristus som jag bär mina bojor;
och de flesta av bröderna hava genom mina bojor blivit så frimodiga i Herren, att de med allt större dristighet våga oförskräckt förkunna Guds ord.
Somliga finnas väl ock, som av avund och trätlystnad predika Kristus, men det finnes också andra som göra det av god vilja.
Dessa senare göra det av kärlek, eftersom de veta att jag är satt till att försvara evangelium.
De förra åter förkunna Kristus av genstridighet, icke med rent sinne, i tanke att de skola tillskynda mig ytterligare bedrövelse i mina bojor.
Vad mer?
Kristus bliver dock på ena eller andra sättet förkunnad, det må nu ske för syns skull eller i uppriktighet; och däröver gläder jag mig.
Ja, jag skall ock framgent få glädja mig;
ty jag vet att detta skall lända mig till frälsning, genom eder förbön och därigenom att Jesu Kristi Ande förlänas mig.
Det är nämligen min trängtan och mitt hopp att jag i intet skall komma på skam, utan att Kristus, nu såsom alltid, skall av mig med all frimodighet bliva förhärligad i min kropp, det må ske genom liv eller genom död.
Ty att leva, det är för mig Kristus, och att dö, det är för mig en vinning.
Men om det att leva i köttet för mig är att utföra ett arbete som bär frukt, vilketdera skall jag då välja?
Det kan jag icke säga.
Jag drages åt båda hållen.
Ty väl åstundar jag att bryta upp och vara hos Kristus, vilket ju vore mycket bättre;
men att jag lever kvar i köttet är för eder skull mer av nöden.
Och då jag är förvissad härom, vet jag att jag skall leva kvar och förbliva hos eder alla, eder till förkovran och glädje i tron,
för att eder berömmelse skall överflöda i Kristus Jesus, i fråga om mig, därigenom att jag ännu en gång kommer till eder.
Fören allenast en sådan vandel som är värdig Kristi evangelium, så att jag -- vare sig jag kommer och besöker eder, eller jag förbliver frånvarande -- får höra om eder att I stån fasta i en och samme Ande och endräktigt kämpen tillsammans för tron på evangelium,
utan att i något stycke låta skrämma eder av motståndarna.
Ty att I så skicken eder är för dem ett vittnesbörd om att de själva gå mot fördärvet, men att I skolen bliva frälsta, och detta av Gud.
Åt eder har ju förunnats icke allenast att tro på Kristus, utan ock att lida för hans skull,
i det att I haven samma kamp som I förr sågen mig hava och nu hören att jag har.
Om nu förmaning i Kristus, om uppmuntran i kärlek, om gemenskap i Anden, om hjärtlig godhet och barmhärtighet betyda något,
gören då min glädje fullkomlig, i det att I ären ens till sinnes, uppfyllda av samma kärlek, endräktiga, liksinnade,
fria ifrån genstridighet och ifrån begär efter fåfänglig ära.
Fasthellre må var och en i ödmjukhet akta den andre förmer än sig själv.
Och sen icke var och en på sitt eget bästa, utan var och en också på andras.
Varen så till sinnes som Kristus Jesus var,
han som var till i Guds-skepnad, men icke räknade jämlikheten med Gud såsom ett byte,
utan utblottade sig själv, i det han antog tjänare-skepnad, när han kom i människogestalt.
Så befanns han i utvärtes måtto vara såsom en människa
och ödmjukade sig och blev lydig intill döden, ja, intill döden på korset.
Därför har ock Gud upphöjt honom över allting och givit honom det namn som är över alla namn
för att i Jesu namn alla knän skola böja sig, deras som äro i himmelen, och deras som äro på jorden, och deras som äro under jorden,
och för att alla tungor skola bekänna, Gud, Fadern, till ära, att Jesus Kristus är Herre.
Därför, mina älskade, såsom I alltid förut haven varit lydiga, så mån I också nu med fruktan och bävan arbeta på eder frälsning, och det icke allenast såsom I gjorden, då jag var närvarande, utan ännu mycket mer nu, då jag är frånvarande.
Ty Gud är den som verkar i eder både vilja och gärning, för att hans goda vilja skall ske.
Gören allt utan att knorra och tveka,
så att I bliven otadliga och rena, Guds ostraffliga barn mitt ibland »ett vrångt och avogt släkte», inom vilket I lysen såsom himlaljus i världen,
i det att I hållen fast vid livets ord.
Bliven mig så till berömmelse på Kristi dag, till ett vittnesbörd om att jag icke har strävat förgäves och icke förgäves har arbetat.
Men om än mitt blod bliver utgjutet såsom ett drickoffer, när jag förrättar min tempeltjänst och därvid frambär offret av eder tro, så gläder jag mig dock och deltager i allas eder glädje.
Sammalunda mån ock I glädjas och deltaga i min glädje.
Jag hoppas nu i Herren Jesus att snart kunna sända Timoteus till eder, så att ock jag får känna hugnad genom det som jag då hör om eder.
Ty jag har ingen av samma sinne som han, ingen som av så uppriktigt hjärta kommer att hava omsorg om eder.
Allasammans söka de sitt eget, icke vad som hör Kristus Jesus till.
Men hans beprövade trohet kännen I; I veten huru han med mig har verkat i evangelii tjänst, såsom en son tjänar sin fader.
Honom hoppas jag alltså kunna sända, så snart jag har fått se huru det går med min sak.
Och i Herren är jag viss om att jag också själv snart skall få komma.
Emellertid har jag funnit det nödvändigt att sända brodern Epafroditus, min medarbetare och medkämpe, tillbaka till eder, honom som I haven skickat hit, för att å edra vägnar överlämna åt mig vad jag kunde behöva.
Ty han längtar efter eder alla och har ingen ro, därför att I haven hört honom vara sjuk.
Han har också verkligen varit sjuk, ja, nära döden, men Gud förbarmade sig över honom; och icke allenast över honom, utan också över mig, för att jag icke skulle få bedrövelse på bedrövelse.
Därför är jag så mycket mer angelägen att sända honom, både för att I skolen få glädjen att återse honom, och för att jag själv därigenom skall få lättnad i min bedrövelse.
Tagen alltså emot honom i Herren, med all glädje, och hållen sådana män i ära.
Ty för Kristi verks skull var han nära döden, i det han satte sitt liv på spel, för att giva mig ersättning för den tjänst som jag måste sakna från eder personligen.
För övrigt, mina bröder, glädjen eder i Herren.
Att skriva till eder detsamma som förut, det räknar jag icke för något besvär, och det är för eder tryggare.
Given akt på de hundarna, given akt på de onda arbetarna, given akt på »de sönderskurna».
Ty vi äro »de omskurna», vi som genom Guds Ande tjäna Gud och berömma oss av Kristus Jesus och icke förtrösta på köttet --
fastän jag för min del väl också kunde hava skäl att förtrösta på köttet.
Ja, om någon menar sig kunna förtrösta på köttet, så kan jag det ännu mer,
jag som blev omskuren, när jag var åtta dagar gammal, jag som är av Israels folk och av Benjamins stam, en hebré, född av hebréer, jag som i fråga om lagen har varit en farisé,
i fråga om nitälskan varit en församlingens förföljare, i fråga om rättfärdighet -- den som vinnes i kraft av lagen -- varit en ostrafflig man.
Men allt det som var mig en vinning, det har jag för Kristi skull räknat såsom en förlust.
Ja, jag räknar i sanning allt såsom förlust mot det som är långt mer värt: kunskapen om Kristus Jesus, min Herre.
Ty det är för hans skull som jag har gått förlustig alltsammans och nu räknar det såsom avskräde, på det att jag må vinna Kristus
och bliva funnen i honom, icke med min egen rättfärdighet, den som kommer av lag, utan med den rättfärdighet som kommer genom tro på Kristus, rättfärdigheten av Gud, på grund av tron.
Ty jag vill lära känna honom och hans uppståndelses kraft och få känna delaktighet i hans lidanden, i det jag bliver honom lik genom en död sådan som hans,
om jag så skulle kunna nå fram till uppståndelsen från de döda.
Icke som om jag redan hade vunnit det eller redan hade blivit fullkomlig, men jag far efter att vinna det, eftersom jag själv har blivit vunnen av Kristus Jesus.
Ja, mina bröder, jag håller icke före att jag ännu har vunnit det, men ett gör jag: jag förgäter det som är bakom mig och sträcker mig mot det som är framför mig
och jagar mot målet, för att få den segerlön som hålles framför oss genom Guds kallelse ovanifrån, i Kristus Jesus.
Må därför vi alla som äro »fullkomliga» hava ett sådant tänkesätt.
Men om så är, att I i något stycke haven andra tankar, så skall Gud också däröver giva eder klarhet.
Dock, såvitt vi redan hava hunnit något framåt, så låtom oss vandra vidare på samma väg.
Mina bröder, varen ock I mina efterföljare, och sen på dem som vandra på samma sätt som jag, eftersom I ju haven oss till föredöme.
Ty det är såsom jag ofta har sagt eder och nu åter måste säga under tårar: många vandra såsom fiender till Kristi kors,
och deras ände är fördärv; de hava buken till sin Gud och söka sin ära i det som är deras skam, och deras sinne är vänt till det som hör jorden till.
Vi åter hava vårt medborgarskap i himmelen, och därifrån vänta vi ock Herren Jesus Kristus såsom Frälsare,
vilken skall så förvandla vår förnedringskropp, att den bliver lik hans härlighetskropp -- genom den kraft varmed han ock kan underlägga sig allt.
Därför, mina älskade och efterlängtade bröder, min glädje och min krona, stån fasta i Herren med detta sinne, I mina älskade.
Evodia förmanar jag, och Syntyke förmanar jag att de skola vara ens till sinnes i Herren.
Ja, också till dig, min Synsygus -- du som med rätta bär det namnet -- har jag en bön: Var dessa kvinnor till hjälp, ty jämte mig hava de kämpat i evangelii tjänst, de såväl som Klemens och mina andra medarbetare, vilkas namn äro skrivna i livets bok.
Glädjen eder i Herren alltid.
Åter vill jag säga: Glädjen eder.
Låten edert saktmod bliva kunnigt för alla människor.
Herren är nära!
Gören eder intet bekymmer, utan låten i allting edra önskningar bliva kunniga inför Gud, genom åkallan och bön, med tacksägelse.
Så skall Guds frid, som övergår allt förstånd, bevara edra hjärtan och edra tankar, i Kristus Jesus.
För övrigt, mina bröder, vad sant är, vad värdigt, vad rätt, vad rent är, vad som är älskligt och värt att akta, ja, allt vad dygd heter, och allt som förtjänar att prisas -- tänken på allt sådant.
Detta, som I haven lärt och inhämtat och haven hört av mig och sett hos mig, det skolen I göra; och så skall fridens Gud vara med eder.
Det har varit för mig en stor glädje i Herren att I nu omsider haven kommit i en så god ställning, att I haven kunnat tänka på mitt bästa.
Dock, I tänkten nog också förut därpå, men I haden icke tillfälle att göra något.
Icke som om jag härmed ville säga att något har fattats mig; ty jag har lärt mig att vara nöjd med de omständigheter i vilka jag är.
Jag vet att finna mig i ringhet, jag vet ock att finna mig i överflöd.
Med vilken ställning och vilka förhållanden som helst är jag förtrogen: jag kan vara mätt, och jag kan vara hungrig; jag kan hava överflöd, och jag kan lida brist.
Allt förmår jag i honom som giver mig kraft.
Dock gjorden I väl däri att I visaden mig deltagande i mitt betryck.
I veten ju ock själva, I filipper, att under evangelii första tid, då när jag hade dragit bort ifrån Macedonien, ingen annan församling än eder trädde i sådan förbindelse med mig, att räkning kunde föras över »utgivet och mottaget».
Ty medan jag ännu var i Tessalonika, sänden I mig både en och två gånger vad jag behövde. --
Icke som om jag skulle åstunda själva gåvan; nej, vad jag åstundar är en sådan frukt därav, som rikligen kommer eder själva till godo.
Jag har nu fått ut allt, och det i överflödande mått.
Jag har fullt upp, sedan jag av Epafroditus har mottagit eder gåva, »en välbehaglig lukt», ett offer som täckes Gud och behagar honom väl.
Så skall ock min Gud, efter sin rikedom, i fullt mått och på ett härligt sätt i Kristus Jesus giva eder allt vad I behöven.
Men vår Gud och Fader tillhör äran i evigheternas evigheter.
Amen.
Hälsen var och en av de heliga i Kristus Jesus.
De bröder som äro här hos mig hälsa eder.
Alla de heliga hälsa eder, först och främst de som höra till kejsarens hus.
Herrens, Jesu Kristi, nåd vare med eder ande.
Paulus, genom Guds vilja Kristi Jesu apostel, så ock brodern Timoteus,
hälsar de heliga som bo i Kolosse, de troende bröderna i Kristus.
Nåd vare med eder och frid ifrån Gud, vår Fader.
Vi tacka Gud, vår Herres, Jesu Kristi, Fader, alltid för eder i våra böner,
ty vi hava hört om eder tro i Kristus Jesus och om den kärlek som I haven till alla de heliga;
vi tacka honom för det hopps skull, som är förvarat åt eder i himmelen.
Om detta hopp haven I redan förut fått höra, genom sanningens ord i det evangelium
som har kommit till eder, likasom det ock är att finna överallt i världen och där bär frukt och växer till, på samma sätt som det har gjort bland eder, allt ifrån den dag, då I hörden det och lärden i sanning känna Guds nåd.
Det var ju en sådan undervisning I mottogen av Epafras, vår älskade medtjänare, som i vårt ställe är eder en trogen Kristi tjänare;
det är också han som för oss har omtalat eder kärlek i Anden.
Allt ifrån den dag då vi fingo höra härom, hava vi därför, å vår sida, icke upphört att bedja för eder och bönfalla om att I mån bliva uppfyllda av kunskap om Guds vilja, i allt slags andlig vishet och andligt förstånd.
Så skolen I kunna föra en vandel som är värdig Herren, honom i allt till behag, och genom kunskapen om Gud bära frukt och växa till i allt gott verk.
Och genom hans härliga makt skolen I på allt sätt uppfyllas av kraft till att bevisa ståndaktighet och tålamod i allt;
och I skolen med glädje tacka Fadern, som har gjort eder skickliga till delaktighet i den arvslott som de heliga hava i ljuset.
Ty han har frälst oss från mörkrets välde och försatt oss i sin älskade Sons rike.
I honom hava vi förlossningen, förlåtelsen för våra synder,
i honom som är den osynlige Gudens avbild och förstfödd före allt skapat.
Ty i honom skapades allt i himmelen och på jorden, synligt såväl som osynligt, både tronänglar och herrar och furstar och väldigheter i andevärlden.
Alltsammans har blivit skapat genom honom och till honom.
Ja, han är till före allt annat, och alltsammans äger bestånd i honom.
Och han är huvudet för kroppen, det är församlingen, han som är begynnelsen, den förstfödde ifrån de döda.
Så skulle han i allt vara den främste.
Ty det behagade Gud att låta all fullhet taga sin boning i honom
och att genom honom försona allt med sig, sedan han genom blodet på hans kors hade berett frid.
Ja, genom honom skulle så ske med allt vad på jorden och i himmelen är.
Också åt eder, som förut voren bortkomna från honom och genom edert sinnelag hans fiender, i det att I gjorden vad ont var,
också åt eder har han nu skaffat försoning i hans jordiska kropp, genom hans död, för att kunna ställa eder fram inför sig heliga och obefläckade och ostraffliga --
om I nämligen förbliven i tron, väl grundade och fasta, utan att låta rubba eder från det hopp som tillbjudes oss i evangelium, det evangelium som I haven hört, och som blivit predikat bland allt skapat under himmelen, det vars tjänare jag, Paulus, har blivit.
Nu gläder jag mig mitt i mina lidanden för eder; och vad som fattas i det mått av Kristus-bedrövelser som jag i mitt kött måste utstå, det uppfyller jag nu för hans kropp, som är församlingen.
Ty dennas tjänare har jag blivit, i enlighet med det uppdrag av Gud, som har blivit mig givet, att jag nämligen överallt skall för eder förkunna Guds ord,
den hemlighet som tidsåldrar och släkten igenom hade varit fördold, men som nu har blivit uppenbarad för hans heliga.
Ty för dem ville Gud kungöra huru rik på härlighet den är bland hedningarna, denna hemlighet, vilken är »Kristus i eder, vårt härlighetshopp».
Och honom förkunna vi för vår del, i det vi förmana var människa och undervisa var människa med all vishet, för att kunna ställa fram var människa såsom fullkomlig i Kristus.
Och för det målet arbetar och kämpar jag, i enlighet med hans kraft, som mäktigt verkar i mig.
Jag vill nämligen, att I skolen veta, vilken kamp jag har att utstå för eder och för församlingen i Laodicea och för alla de andra som icke personligen hava sett mitt ansikte.
Ty jag önskar, att deras hjärtan skola få hugnad, därigenom att de slutas tillsammans i kärlek och komma till en full förståndsvisshets hela rikedom, till en rätt kunskap om Guds hemlighet, vilken är Kristus;
ty i honom finnas visdomens och kunskapens alla skatter fördolda.
Detta säger jag, för att ingen skall bedraga eder med skenfagert tal.
Ty om jag ock till kroppen är frånvarande, så är jag dock i anden hos eder och gläder mig, när jag ser den ordning, som råder bland eder, och när jag ser fastheten i eder tro på Kristus.
Såsom I nu haven mottagit Kristus Jesus, Herren, så vandren i honom
och varen rotade i honom och låten eder uppbyggas i honom och befästas i tron, i enlighet med den undervisning I haven fått, och överflöden i tacksägelse.
Sen till, att ingen får bortföra eder såsom ett segerbyte genom sin tomma och bedrägliga »vishetslära», i det att han åberopar fäderneärvda människomeningar och håller sig till världens »makter» och icke till Kristus.
Ty i honom bor gudomens hela fullhet lekamligen,
och i honom haven I blivit delaktiga av den fullheten, i honom som är huvudet för alla andevärldens furstar och väldigheter.
I honom haven I ock blivit omskurna genom en omskärelse, som icke skedde med händer, en som bestod däri att I bleven avklädda eder köttsliga kropp; jag menar omskärelsen i Kristus.
I haven ju med honom blivit begravna i dopet; I haven ock i dopet blivit uppväckta med honom, genom tron på Guds kraft, hans som uppväckte honom från de döda.
Ja, också eder som voren döda genom edra synder och genom edert kötts oomskurenhet, också eder har han gjort levande med honom; ty han har förlåtit oss alla våra synder.
Han har nämligen utplånat den handskrift som genom sina stadgar anklagade oss och låg oss i vägen; den har han skaffat undan genom att nagla den fast vid korset.
Han har avväpnat andevärldens furstar och väldigheter och låtit dem bliva till skam inför alla, i det att han i honom har triumferat över dem.
Låten därför ingen döma eder i fråga om mat och dryck eller angående högtid eller nymånad eller sabbat.
Sådant är allenast en skuggbild av vad som skulla komma, men verkligheten själv finnes hos Kristus.
Låten icke segerlönen tagas ifrån eder av någon som har sin lust i »ödmjukhet» och ängladyrkan och gör sig stor med sina syner, någon som utan orsak är uppblåst genom sitt köttsliga sinne
och icke håller sig till honom som är huvudet, honom från vilken hela kroppen vinner sin tillväxt i Gud, i det att den av sina ledgångar och senor får bistånd och sammanhållning.
Om I nu haven dött med Kristus och så blivit frigjorda ifrån världens »makter», varför låten I då allahanda stadgar läggas på eder, likasom levden I ännu i världen:
»Det skall du icke taga i», »Det skall du icke smaka», »Det skall du icke komma vid»,
och detta när det gäller ting, som alla äro bestämda till att gå under genom förbrukning -- allt till åtlydnad av människobud och människoläror?
Visserligen har allt detta fått namn om sig att vara »vishet», eftersom däri ligger ett självvalt gudstjänstväsende och ett slags »ödmjukhet» och en kroppens späkning; men ingalunda ligger däri »en viss heder», det tjänar allenast till att nära det köttsliga sinnet.
Om I alltså ären uppståndna med Kristus, så söken det som är därovan, där varest Kristus är och sitter på Guds högra sida.
Ja, haven edert sinne vänt till det som är därovan, icke till det som är på jorden.
Ty I haven dött, och edert liv är fördolt med Kristus i Gud.
När Kristus, han som är vårt liv, bliver uppenbarad, då skolen ock I med honom bliva uppenbarade i härlighet.
Så döden nu edra lemmar, som höra jorden till: otukt, orenhet, lusta, ond begärelse, så ock girigheten, som ju är avgudadyrkan;
ty för sådant kommer Guds vrede.
I de synderna vandraden också I förut, då I ännu haden edert liv i dem.
Men nu skolen också I lägga bort alltsammans; vrede, häftighet, ondska, smädelse och skamligt tal ur eder mun;
I skolen icke ljuga på varandra.
I haven ju avklätt eder den gamla människan med hennes gärningar
och iklätt eder den nya, den som förnyas till sann kunskap och så bliver en avbild av honom som har skapat henne.
Och därvid kommer det icke an på om någon är grek eller jude, omskuren eller oomskuren, barbar eller skyt, träl eller fri; nej, Kristus är allt och i alla.
Så kläden eder nu såsom Guds utvalda, hans heliga och älskade, i hjärtlig barmhärtighet, godhet, ödmjukhet, saktmod, tålamod.
Och haven fördrag med varandra och förlåten varandra, om någon har något att förebrå en annan.
Såsom Herren har förlåtit eder, så skolen ock I förlåta.
Men över allt detta skolen I ikläda eder kärleken, ty den är fullkomlighetens sammanhållande band.
Och låten Kristi frid regera i edra hjärtan; ty till att äga den ären I ock kallade såsom lemmar i en och samma kropp.
Och varen tacksamma.
Låten Kristi ord rikligen bo ibland eder; undervisen och förmanen varandra i all vishet, med psalmer och lovsånger och andliga visor, och sjungen med tacksägelse till Guds ära i edra hjärtan.
Och allt, vadhelst I företagen eder i ord eller gärning, gören det allt i Herren Jesu namn och tacken Gud, Fadern, genom honom.
I hustrur, underordnen eder edra män, såsom tillbörligt är i Herren.
I män, älsken edra hustrur och varen icke bittra mot dem.
I barn, varen edra föräldrar lydiga i allt, ty detta är välbehagligt i Herren.
I fäder, reten icke edra barn, på det att de icke må bliva klenmodiga.
I tjänare, varen i allt edra jordiska herrar lydiga, icke med ögontjänst, av begär att behaga människor, utan av uppriktigt hjärta, i Herrens fruktan.
Vadhelst I gören, gören det av hjärtat, såsom tjänaden I Herren och icke människor.
I veten ju, att I till vedergällning skolen av Herren få eder arvedel; den herre I tjänen är Kristus.
Den som gör orätt, han skall få igen den orätt han har gjort, utan anseende till personen.
I herrar, given edra tjänare, vad rätt och billigt är; I veten ju, att också I haven en herre i himmelen.
Varen uthålliga i bönen och vaken i den under tacksägelse.
Och bedjen jämväl för oss, att Gud må åt oss öppna en dörr för ordet, så att vi få förkunna Kristi hemlighet, den hemlighet, för vars skull jag också är en fånge;
ja, bedjen, att jag må uppenbara den med de rätta orden.
Skicken eder visligt mot dem som stå utanför och tagen väl i akt vart lägligt tillfälle.
Edert tal vare alltid välbehagligt, kryddat med salt; I bören förstå, huru I skolen svara var och en.
Om allt vad mig angår skall min älskade broder Tykikus, min trogne tjänare och min medtjänare i Herren, underrätta eder.
Honom sänder jag till eder, just för att I skolen få veta, huru det är med oss, och för att han skall hugna edra hjärtan.
Tillika sänder jag Onesimus, min trogne och älskade broder, eder landsman.
De skola underrätta eder om allting här.
Aristarkus, min medfånge, hälsar eder; så gör ock Markus, Barnabas syskonbarn.
Angående honom haven I redan fått föreskrifter; och om han kommer till eder, så tagen vänligt emot honom.
Också Jesus, som kallas Justus, hälsar eder.
Av de omskurna äro dessa mina enda medarbetare för Guds rike, och de hava varit mig till hugnad.
Epafras, eder landsman, hälsar eder, en Kristi Jesu tjänare, som i sina böner alltid kämpar för eder, för att I skolen stå fasta och vara fullkomliga och fullt vissa i allt som är Guds vilja.
Ty jag giver honom det vittnesbördet, att han har stor möda för eder likasom ock för dem som bo i Laodicea och i Hierapolis.
Lukas, läkaren, den älskade brodern, hälsar eder; så gör ock Demas.
Hälsen bröderna i Laodicea, så ock Nymfas tillika med den församling som kommer tillhopa i hans hus.
Sedan detta brev har blivit uppläst hos eder, så sörjen för att det ock bliver uppläst i laodicéernas församling och att jämväl I fån läsa det brev, som kommer från Laodicea.
Sägen ock detta till Arkippus: »Hav akt på det ämbete, som du har undfått i Herren, så att du fullgör, vad därtill hör.»
Här skriver jag, Paulus, min hälsning med egen hand.
Tänken på mina bojor.
Nåd vare med eder.
Paulus och Silvanus och Timoteus hälsa tessalonikernas församling i Gud, Fadern, och Herren Jesus Kristus.
Nåd och frid vare med eder.
Vi tacka Gud alltid för eder alla, när vi tänka på eder i våra böner.
Ty oavlåtligen ihågkomma vi inför vår Gud och Fader edra gärningar i tron och edert arbete i kärleken och eder ståndaktighet i hoppet, i vår Herre Jesus Kristus.
Vi veta ju, käre bröder, i Guds älskade, huru det var, när I bleven utvalda:
vårt evangelium kom till eder icke med ord allenast, utan i kraft och helig ande och med full visshet.
I veten ock på vad sätt vi uppträdde bland eder, till edert bästa.
Och I å eder sida bleven våra efterföljare och därmed Herrens, i det att I, mitt under stort betryck, togen emot ordet med glädje i helig ande.
Så bleven I själva ett föredöme för alla de troende i Macedonien och Akaja.
Ty från eder har genljudet av Herrens ord gått vidare ut; icke allenast i Macedonien och Akaja, utan allestädes har eder tro på Gud blivit känd, så att vi för vår del icke behöva tala något därom.
Ty själva förkunna de om oss, med vilken framgång vi begynte vårt arbete hos eder, och huru I från avgudarna omvänden eder till Gud, till att tjäna den levande och sanne Guden,
och till att vänta hans Son från himmelen, honom som han har uppväckt från de döda, Jesus, som frälsar oss undan den kommande vredesdomen.
I veten ju själva, käre bröder, att det icke var utan kraft vi begynte vårt arbete hos eder.
Nej, fastän vi, såsom i veten, i Filippi förut hade fått utstå lidande och misshandling, hade vi dock frimodighet i vår Gud till att förkunna för eder Guds evangelium, under mycken kamp.
Ty vad vi tala till tröst och förmaning, det har icke sin grund i villfarelse eller i orent uppsåt, ej heller sker det med svek;
utan därför att vi av Gud hava prövats värdiga att få evangelium oss betrott, tala vi i enlighet därmed, icke för att vara människor till behag, utan för att vara Gud till behag, honom som prövar våra hjärtan.
Aldrig någonsin hava vi uppträtt med smickrets ord, det veten I, ej heller så, att vi skulle få en förevändning att bereda oss vinning -- Gud är vårt vittne.
Ej heller hava vi sökt pris av människor, vare sig av eder eller av andra,
fastän vi såsom Kristi apostlar väl hade kunnat uppträda med myndighet.
Tvärtom hava vi visat oss milda bland eder, såsom när en moder omhuldar sina späda barn.
I sådan ömhet om eder ville vi gärna icke allenast göra också eder delaktiga av Guds evangelium, utan till och med offra våra liv för eder, ty I haden blivit oss kära.
I kommen ju ihåg, käre bröder, vårt arbete och vår möda, huru vi, under det att vi predikade för eder Guds evangelium, strävade natt och dag, för att icke bliva någon av eder till tunga.
I själva ären våra vittnen, och Gud är vårt vittne, I veten, och han vet huru heligt och rättfärdigt och ostraffligt vi förhöllo oss mot eder, I som tron.
Likaledes veten I huru vi förmanade och uppmuntrade var och en av eder, såsom en fader sina barn,
och huru vi uppfordrade eder att föra en vandel som vore värdig Gud, honom som kallar eder till sitt rike och sin härlighet.
Därför tacka vi ock oavlåtligen Gud för att I, när I undfingen det Guds ord som vi predikade, icke mottogen det såsom människoord, utan såsom Guds ord, vilket det förvisso är, ett ord som ock är verksamt i eder som tron.
I, käre bröder, haven ju blivit efterföljare till de Guds församlingar i Kristus Jesus som äro i Judeen.
Ty I haven av edra egna landsmän fått lida detsamma som de hava lidit av judarna --
av dem som dödade både Herren Jesus och profeterna och förjagade oss, och som äro misshagliga för Gud och fiender till alla människor,
i det att de söka hindra oss att tala till hedningarna, så att dessa kunna bliva frälsta.
Så uppfylla de alltjämt sina synders mått.
Dock, vredesdomen har kommit över dem i all sin stränghet.
Men då vi nu hava måst vara skilda från eder, käre bröder -- visserligen allenast för en kort tid och i utvärtes måtto, icke till hjärtat -- hava vi blivit så mycket mer angelägna att få se edra ansikten och känt stor åstundan därefter.
Ty vi hava varit redo att komma till eder -- jag, Paulus, för min del både en och två gånger -- men Satan har hindrat oss.
Ty vem är vårt hopp och vår glädje och vår berömmelses krona inför vår Herre Jesus vid hans tillkommelse, vem, om icke just I?
Ja, I ären vår ära och vår glädje.
Därför, när vi icke mer kunde uthärda, beslöto vi att stanna ensamma kvar i Aten,
och sände åstad Timoteus, vår broder och Guds tjänare vid förkunnandet av evangelium om Kristus, för att han skulle styrka och uppmuntra eder i eder tro,
så att ingen bleve vacklande under dessa lidanden.
Ty I veten själva att sådana äro oss förelagda.
Redan när vi voro hos eder, sade vi ju eder förut att vi skulle komma att utstå lidanden.
Så har nu ock skett, det veten I.
Det var också därför som jag sände honom åstad, när jag icke mer kunde uthärda; ty jag ville veta något om eder tro, eftersom jag fruktade att frestaren till äventyrs hade så frestat eder, att vårt arbete skulle bliva utan frukt.
Men nu, då Timoteus har kommit till oss från eder och förkunnat för oss det glada budskapet om eder tro och kärlek, och sagt oss att I alltjämt haven oss i god hågkomst, och att I längten efter att se oss, likasom vi längta efter eder,
nu hava vi i fråga om eder, käre bröder, genom eder tro fått hugnad i all vår nöd och allt vårt lidande.
Ty nu leva vi, eftersom I stån fasta i Herren.
Ja, huru skola vi nog kunna tacka Gud för eder, till gengäld för all den glädje som vi genom eder hava inför vår Gud?
Natt och dag är det vår innerligaste bön, att vi må få se edra ansikten och avhjälpa vad som kan brista i eder tro.
Men vår Gud och Fader själv och vår Herre Jesus må för oss jämna vägen till eder.
Och eder må Herren giva en allt större och mer överflödande kärlek till varandra, ja, till alla människor, en sådan kärlek som vi hava till eder,
så att edra hjärtan styrkas till att vara ostraffliga i helighet inför vår Gud och Fader vid vår Herre Jesu tillkommelse, när han kommer med alla sina heliga.
Ytterligare, käre bröder, bedja vi nu och förmana eder i Herren Jesus att allt mer förkovra eder i en sådan vandel som I haven fått lära av oss att I skolen föra, Gud till behag -- en sådan vandel som I redan fören.
I veten ju vilka bud vi hava givit eder genom Herren Jesus.
Ty detta är Guds vilja, detta som hör till eder helgelse, att I avhållen eder från otukt,
och att var och en av eder vet att hava sin egen maka i helgelse och ära,
icke i begärelses lusta såsom hedningarna -- vilka icke känna Gud --
och att ingen i sitt förhållande till sin broder kränker honom eller gör honom något förfång, ty Herren är en hämnare över allt detta, såsom vi redan förut hava sagt och betygat för eder.
Gud har ju icke kallat oss till orenhet, utan till att leva i helgelse.
Den som icke vill veta av detta, han förkastar alltså icke en människa, utan Gud, honom som giver sin helige Ande till att bo i eder.
Om broderlig kärlek är det icke behövligt att skriva till eder, ty I haven själva fått lära av Gud att älska varandra;
så handlen I ju ock mot alla bröderna i hela Macedonien.
Men vi förmana eder, käre bröder, att allt mer förkovra eder häri
och att sätta eder ära i att leva i stillhet och sköta vad eder åligger och arbeta med edra händer, enligt vad vi hava bjudit eder,
så att I skicken eder höviskt mot dem som stå utanför och icke behöven anlita någons hjälp.
Vi vilja icke lämna eder, käre bröder, i okunnighet om huru det förhåller sig med dem som avsomna, för att I icke skolen sörja såsom de andra, de som icke hava något hopp.
Ty lika visst som Jesus, såsom vi tro, har dött och har uppstått, lika visst skall ock Gud genom Jesus föra dem som äro avsomnade fram jämte honom.
Såsom ett ord från Herren säga vi eder nämligen detta, att vi som leva och lämnas kvar till Herrens tillkommelse ingalunda skola komma före dem som äro avsomnade.
Ty Herren skall själv stiga ned från himmelen, och ett maktbud skall ljuda, en överängels röst och en Guds basun.
Och först skola de i Kristus döda uppstå;
sedan skola vi som då ännu leva och hava lämnats kvar bliva jämte dem bortryckta på skyar upp i luften, Herren till mötes; och så skola vi alltid få vara hos Herren.
Så trösten nu varandra med dessa ord.
Vad åter angår tid och stund härför, så är det icke behövligt att därom skriva till eder, käre bröder.
Ty I veten själva nogsamt att Herrens dag kommer såsom en tjuv om natten.
Bäst de säga: »Allt står väl till, och ingen fara är på färde», då kommer plötsligt fördärv över dem, såsom födslovåndan över en havande kvinna, och de skola förvisso icke kunna fly undan.
Men I, käre bröder, I leven icke mörker, så att den dagen kan komma över eder såsom en tjuv;
I ären ju alla ljusets barn och dagens barn.
Ja, vi höra icke natten eller mörkret till;
låtom oss alltså icke sova såsom de andra, utan låtom oss vaka och vara nyktra.
De som sova, de sova om natten, och de som dricka sig druckna, de äro druckna om natten;
men vi som höra dagen till, vi må vara nyktra, iklädda trons och kärlekens pansar, med frälsningens hopp såsom hjälm.
Ty Gud har icke bestämt oss till att drabbas av vrede, utan till att vinna frälsning genom vår Herre, Jesus Kristus,
som har dött för oss, på det att vi må leva tillika med honom, vare sig vi ännu äro vakna eller vi äro avsomnade.
Trösten därför varandra, och uppbyggen varandra inbördes, såsom I ock redan gören.
Vi bedja eder, käre bröder, att rätt uppskatta de män som arbeta bland eder, och som äro edra föreståndare i Herren och förmana eder.
Låten dem vara eder övermåttan kära, för det verks skull som de utföra.
Hållen frid inbördes.
Vi bjuda eder, käre bröder: Förmanen de oordentliga, uppmuntren de klenmodiga, tagen eder an de svaga, visen tålamod mot var man.
Sen till, att ingen vedergäller någon med ont för ont; faren fastmer alltid efter att göra vad gott är mot varandra och mot var man.
Varen alltid glada.
Bedjen oavlåtligen.
Tacken Gud i alla livets förhållanden.
Ty att I så gören är Guds vilja i Kristus Jesus.
Utsläcken icke Anden,
förakten icke profetisk tal,
men pröven allt, behållen vad gott är,
avhållen eder från allt ont, av vad slag det vara må.
Men fridens Gud själv helge eder till hela eder varelse, så att hela eder ande och eder själ och eder kropp finnas bevarade ostraffliga vid vår Herres, Jesu Kristi, tillkommelse.
Trofast är han som kallar eder; han skall ock utföra sitt verk.
Käre bröder, bedjen för oss.
Hälsen alla bröderna med en helig kyss.
Jag besvär eder vid Herren att låta uppläsa detta brev för alla bröderna.
Vår Herres, Jesu Kristi, nåd vare med eder.
Paulus och Silvanus och Timoteus hälsa tessalonikernas församling i Gud, vår Fader, och Herren Jesus Kristus.
Nåd vare med eder och frid ifrån Gud, Fadern, och Herren Jesus Kristus.
Vi äro pliktiga att alltid tacka Gud för eder, käre bröder, såsom tillbörligt är, därför att eder tro så mäktigt tillväxer, och den kärlek I haven till varandra mer och mer förökas hos eder alla och hos envar av eder.
Därför kunna vi själva i Guds församlingar berömma oss av eder, i fråga om eder ståndaktighet och eder tro under alla edra förföljelser, och under de lidanden I måsten uthärda.
Sådant är ett vittnesbörd om att Guds dom bliver rättvis.
Så skolen I aktas värdiga Guds rike; för dess skull är det ock som I liden.
Guds rättfärdighet kräver ju att de som vålla eder lidande få lidande till vedergällning,
men att I som utstån lidanden fån hugnad tillsammans med oss, när Herren Jesus uppenbarar sig från himmelen med sin makts änglar,
»i lågande eld», och låter straffet drabba dem som icke känna Gud, och dem som icke äro vår Herre Jesu evangelium lydiga.
Dessa skola då bliva straffade med evigt fördärv, bort undan Herrens ansikte och hans överväldigande härlighet,
när han kommer för att förhärligas i sina heliga och visa sig underbar i alla dem som hava kommit till att tro; ty det vittnesbörd vi hava framburit till eder haven I trott.
Så skall ske på den dagen.
Fördenskull bedja vi ock alltid för eder, att vår Gud må akta eder värdiga sin kallelse, och att han må med kraft fullborda i eder allt vad en god vilja kan åstunda, och vad tro kan verka,
så att vår Herre Jesu namn bliver förhärligat i eder, och I i honom, efter vår Guds och Herrens, Jesu Kristi, nåd.
I fråga om vår Herres, Jesu Kristi, tillkommelse, och huru vi skola församlas till honom, bedja vi eder, käre bröder,
att I icke -- vare sig genom någon »andeingivelse» eller på grund av något ord eller något brev, som förmenas komma från oss -- så hastigt låten eder bringas ur fattningen och förloren besinningen, som om Herrens dag redan stode för dörren.
Låten ingen bedraga eder om vad sätt det vara må.
Ty först måste avfallet hava skett och »Laglöshetens människa», fördärvets man, hava trätt fram,
vedersakaren, som upphäver sig över allt vad gud heter, och allt som kallas heligt, så att han tager sitt säte i Guds tempel och föregiver sig vara Gud.
Kommen I icke ihåg att jag sade eder detta, medan jag ännu var hos eder?
Och I veten vad det är som nu håller honom tillbaka, så att han först när hans tid är inne kan träda fram.
Redan är ju laglöshetens hemlighet verksam; allenast måste den som ännu håller tillbaka först skaffas ur vägen.
Sedan skall »den Laglöse» träda fram, och honom skall då Herren Jesus döda med sin muns anda och tillintetgöra genom sin tillkommelses uppenbarelse --
honom som efter Satans tillskyndelse kommer med lögnens alla kraftgärningar och tecken och under
och med orättfärdighetens alla bedrägliga konster, för att bedraga dem som gå förlorade, till straff därför att de icke gåvo kärleken till sanningen rum, så att de kunde bliva frälsta.
Därför sänder ock Gud över dem villfarelsens makt, så att de sätta tro till lögnen,
för att de skola bliva dömda, alla dessa som icke hava satt tro till sanningen, utan funnit behag i orättfärdigheten.
Men vi för vår del äro pliktiga att alltid tacka Gud för eder käre bröder, I Herrens älskade, därför att Gud från begynnelsen har utvalt eder till frälsning, i helgelse i Anden och i tro på sanningen.
Härtill har han ock genom vårt evangelium kallat eder, för att I skolen bliva delaktiga av vår Herres, Jesu Kristi, härlighet.
Stån alltså fasta, käre bröder, och hållen eder vid de lärdomar som I haven mottagit av oss, vare sig muntligen eller genom brev.
Och vår Herre Jesus Kristus själv och Gud, vår Fader, som har älskat oss och i nåd berett oss en evig hugnad och givit oss ett gott hopp,
han hugne edra hjärtan, och styrke eder till allt vad gott är, både i gärning och i ord.
För övrigt, käre bröder, bedjen för oss, att Herrens ord må hava framgång och komma till ära hos andra likasom hos eder,
så ock att vi må bliva frälsta ifrån vanartiga och onda människor.
Ty tron är icke var mans.
Men Herren är trofast, och han skall styrka eder och bevara eder från det onda.
Och vi hava den tillförsikten till eder i Herren, att I både nu gören och framgent skolen göra vad vi bjuda eder.
Ja, Herren styre edra hjärtan till Guds kärlek och Kristi ståndaktighet.
Men vi bjuda eder, käre bröder, i vår Herres, Jesu Kristi, namn, att I dragen eder ifrån var broder som för en oordentlig vandel och icke lever efter de lärdomar han har mottagit av oss.
I veten ju själva huru man bör efterfölja oss.
Ty vi förhöllo oss icke oordentligt bland eder,
ej heller åto vi någons bröd för intet; tvärtom åto vi vårt bröd under arbete och möda, och vi strävade natt och dag, för att icke bliva någon av eder till tunga.
Icke som om vi ej hade haft rätt därtill, men vi ville låta eder i oss få ett föredöme, för att I skullen efterfölja oss.
Redan när vi voro hos eder, gåvo vi ju eder det budet: om någon icke vill arbeta, så skall han icke heller äta.
Vi höra nämligen att somliga bland eder föra en oordentlig vandel och icke arbeta, utan allenast syssla med sådant som icke kommer dem vid.
Sådana människor bjuda och förmana vi i Herren Jesus Kristus, att de arbeta i stillhet, så att de kunna äta sitt eget bröd.
Och I, käre bröder, mån icke förtröttas att göra vad gott är.
Men om någon icke lyder vad vi hava sagt i detta brev, så märken ut för eder den mannen, och haven intet umgänge med honom, på det att han må blygas.
Hållen honom dock icke för en ovän, utan förmanen honom såsom en broder.
Men fridens Herre själv give eder sin frid alltid och på allt sätt.
Herren vare med eder alla.
Här skriver jag, Paulus, min hälsning med egen hand.
Detta är ett kännetecken i alla mina brev; så skriver jag.
Vår Herres, Jesu Kristi, nåd vare med eder alla.
Paulus, Kristi Jesu apostel, förordnad av Gud, vår Frälsare, och Kristus Jesus, vårt hopp,
hälsar Timoteus, sin sannskyldige son i tron.
Nåd, barmhärtighet och frid ifrån Gud, Fadern, och Kristus Jesus, vår Herre!
Jag bjuder dig, nu såsom när jag for åstad till Macedonien, att stanna kvar i Efesus och där förmana somliga att icke förkunna främmande läror
eller akta på fabler och släktledningshistorier utan ände, som ju snarare vålla ordstrider än främja den Guds ordning som kommer till fullbordan i tron.
Och förmaningens ändamål är kärlek av ett rent hjärta och av ett gott samvete och av en oskrymtad tro.
Från dessa stycken hava somliga farit vilse och vänt sin håg till fåfängligt tal --
människor som vilja vara lärare i lagen, fastän de icke förstå ens vad de själva tala, eller vad de ting äro, som de med sådan säkerhet orda om.
Men vi veta att lagen är god, om man nämligen brukar den såsom lagen bör brukas,
och om man förstår detta, att lagen är till icke för rättfärdiga människor, utan för dem som trotsa lag och myndighet, för ogudaktiga och syndare, oheliga och oandliga människor, fadermördare och modermördare, för mandråpare,
för dem som öva otukt och onaturlig vällustsynd, för dem som äro människosäljare, lögnare, menedare eller något annat som strider mot den sunda läran --
detta i enlighet med det evangelium om den salige Gudens härlighet, varmed jag har blivit betrodd.
Vår Herre Kristus Jesus, som har givit mig kraft, tackar jag för att han har tagit mig i sin tjänst och funnit mig vara förtroende värd,
mig som förut var en hädare och förföljare och våldsverkare.
Men barmhärtighet vederfors mig, eftersom jag icke bättre visste, när jag i min otro handlade så.
Och vår Herres nåd blev så mycket mer överflödande, med tron och kärleken i Kristus Jesus.
Det är ett fast ord och i allo värt att mottagas, att Kristus Jesus har kommit i världen för att frälsa syndare, bland vilka jag är den främste.
Men att barmhärtighet vederfors mig, det skedde just för att Kristus Jesus skulle främst på mig bevisa all sin långmodighet, och låta mig bliva en förstlingsbild av dem som skulle komma att tro på honom och så vinna evigt liv.
Men evigheternas konung, den oförgänglige, osynlige, ende Guden, vare ära och pris i evigheternas evigheter!
Amen.
Att så förmana dem, det ålägger jag dig, min son Timoteus, i enlighet med de profetord som en gång uttalades över dig.
Må du i kraft av dem strida den goda striden,
rustad med tro och med ett gott samvete.
Detta hava nu visserligen somliga skjutit å sido, men de hava därigenom lidit skeppsbrott i tron.
Till dem höra Hymeneus och Alexander, vilka jag har överlämnat åt Satan, för att de skola bliva så tuktade, att de icke vidare smäda.
Så uppmanar jag nu framför allt därtill att man må bedja, åkalla, anropa och tacka Gud för alla människor,
för konungar och all överhet, så att vi kunna föra ett lugnt och stilla liv, på ett i allo fromt och värdigt sätt.
Sådant är gott och välbehagligt inför Gud, vår Frälsare,
som vill att alla människor skola bliva frälsta och komma till kunskap om sanningen.
Ty en enda är Gud, och en enda är medlare emellan Gud och människor: en människa, Kristus Jesus,
han som gav sig själv till lösen för alla, varom ock vittnesbördet skulle frambäras, när tiden var inne.
Och själv har jag blivit satt till att vara dess förkunnare och apostel -- det säger jag med sanning, jag ljuger icke -- ja, till att i tro och sanning vara en lärare för hedningar.
Jag vill alltså att männen allestädes skola förrätta bön, i det att de, fria ifrån vrede och disputerande, upplyfta heliga händer.
Likaledes vill jag att kvinnorna skola uppträda i hövisk dräkt, att de blygsamt och tuktigt pryda sig, icke med hårflätningar och guld eller pärlor eller dyrbara kläder,
utan med goda gärningar, såsom det höves kvinnor som vilja räknas för gudfruktiga.
Kvinnan bör i stillhet låta sig undervisas och därvid helt underordna sig.
Däremot kan jag icke tillstädja en kvinna att själv uppträda såsom lärare, ej heller att råda över sin man; fastmer må hon leva i stillhet.
Adam blev ju först skapad och sedan Eva.
Och Adam blev icke bedragen, men kvinnan blev svårt bedragen och förleddes till överträdelse.
Dock skall kvinnan, under det hon föder sina barn, vinna frälsning, om hon förbliver i tro och kärlek och helgelse, med ett tuktigt väsende.
Det är ett visst ord, att om någons håg står till en församlingsföreståndares ämbete, så är det en god verksamhet han åstundar.
En församlingsföreståndare bör därför vara oförvitlig; han bör vara en enda kvinnas man, nykter och tuktig, hövisk i sitt skick, gästvänlig, väl skickad att undervisa,
icke begiven på vin, icke våldsam, utan foglig, icke stridslysten, fri ifrån penningbegär.
Han bör väl förestå sitt eget hus och hålla sina barn i lydnad, med all värdighet;
ty huru skulle dem som icke vet att förestå sitt eget hus kunna sköta Guds församling?
Han bör icke vara nyomvänd, för att han icke skall förblindas av högmod och så hemfalla under djävulens dom.
Han bör ock hava gott vittnesbörd om sig av dem som stå utanför, så att han icke utsättes för smälek och faller i djävulens snara.
Församlingstjänarna böra likaledes skicka sig värdigt, icke vara tvetaliga, icke benägna för mycket vindrickande, icke snikna efter slem vinning;
de böra äga trons hemlighet i ett rent samvete.
Men också dessa skola först prövas; därefter må de, om de befinnas oförvitliga, få tjäna församlingen.
Är det kvinnor, så böra dessa likaledes skicka sig värdigt, icke gå omkring med förtal, men vara nyktra och trogna i allt.
En församlingstjänare skall vara en enda kvinnas man; han skall hålla god ordning på sina barn och väl förestå sitt hus.
Ty de som hava väl skött en församlingstjänares syssla, de vinna en aktad ställning och kunna i tron, den tro de hava i Kristus Jesus, uppträda med mycken frimodighet.
Detta skriver jag till dig, fastän jag hoppas att snart få komma till dig.
Jag vill nämligen, om jag likväl skulle dröja, att du skall veta huru man bör förhålla sig i Guds hus, som ju är den levande Gudens församling, sanningens stödjepelare och grundfäste.
Och erkänt stor är gudaktighetens hemlighet: »Han som blev uppenbarad i köttet, rättfärdigad i anden, sedd av änglar, predikad bland hedningarna, trodd i världen, upptagen i härligheten.»
Men Anden säger uttryckligen, att i kommande tider somliga skola avfalla från tron och hålla sig till villoandar och till onda andars läror.
Så skall ske genom lögnpredikanters skrymteri, människors som i sina egna samveten äro brännmärkta såsom brottslingar,
och som förbjuda äktenskap och vilja att man skall avhålla sig från allahanda mat, som Gud har skapat till att med tacksägelse mottagas av dem som tro och hava lärt känna sanningen.
Ty allt vad Gud har skapat är gott, och intet är förkastligt, när det mottages med tacksägelse:
det bliver nämligen helgat genom Guds ord och genom bön.
Om du framlägger detta för bröderna, så bevisar du dig såsom en god Kristi Jesu tjänare, då du ju hämtar din näring av trons och den goda lärans ord, den läras som du troget har efterföljt.
Men de oandliga käringfablerna må du visa ifrån dig.
Öva dig i stället själv i gudsfruktan.
Ty lekamlig övning gagnar till litet, men gudsfruktan gagnar till allt; den har med sig löfte om liv, både för denna tiden och för den tillkommande.
Detta är ett fast ord och i allo värt att mottagas.
Ja, därför arbeta och kämpa vi, då vi nu hava satt vårt hopp till den levande Guden, honom som är alla människors Frälsare, först och främst deras som tro.
Så skall du bjuda och undervisa.
Låt ingen förakta dig för din ungdoms skull; fastmer må du för dem som tro bliva ett föredöme i tal och i vandel, i kärlek, i tro och i renhet.
Var nitisk i att föreläsa skriften och i att förmana och undervisa, till dess jag kommer.
Försumma icke att vårda den nådegåva som finnes i dig, och som gavs dig i kraft av profetord, under handpåläggning av de äldste.
Tänk på detta, lev i detta, så att din förkovran bliver uppenbar för alla.
Hav akt på dig själv och på din undervisning, och håll stadigt ut därmed; ty om du så gör, frälsar du både dig själv och dem som höra dig.
En äldre man må du icke tillrättavisa med hårda ord; du bör tala till honom såsom till en fader.
Till yngre män må du tala såsom till bröder,
till äldre kvinnor såsom till mödrar, till yngre kvinnor såsom till systrar, i all renhet.
Änkor må du bevisa ära, om de äro rätta, värnlösa änkor.
Men om en änka har barn eller barnbarn, då må i första rummet dessa lära sig att med tillbörlig vördnad taga sig an sina närmaste och så återgälda sina föräldrar vad de äro dem skyldiga; ty sådant är välbehagligt inför Gud.
En rätt, värnlös änka, som sitter ensam, hon har sitt hopp i Gud och håller ut i bön och åkallan natt och dag.
Men en sådan som allenast gör sig goda dagar, hon är död, fastän hon lever. --
Förehåll dem också detta, så att man icke får något att förevita dem.
Men om någon icke drager försorg om sina egna, först och främst om sina närmaste, så har denne förnekat sin tro och är värre än en otrogen.
Såsom »församlingsänka» må ingen annan uppföras än den som är minst sextio år gammal, och som har varit allenast en mans hustru,
en som har det vittnesbördet om sig, att hon har övat goda gärningar, uppfostrat barn, givit härbärge åt husvilla, tvagit heligas fötter, understött nödlidande, korteligen, beflitat sig om allt gott verk.
Unga änkor skall du däremot icke antaga.
Ty när de hava njutit nog av Kristus, vilja de åter gifta sig;
och de äro då hemfallna åt dom, eftersom de hava brutit sin första tro.
Därtill lära de sig ock att vara lättjefulla, i det att de löpa omkring i husen; ja, icke allenast att vara lättjefulla, utan ock att vara skvalleraktiga och att syssla med sådant som icke kommer dem vid, allt medan de tala vad otillbörligt är.
Därför vill jag att unga änkor gifta sig, föda barn, förestå var och en sitt hus och icke giva någon motståndare anledning att smäda.
Redan hava ju några vikit av och följt efter Satan.
Om någon troende, vare sig man eller kvinna, har änkor att sörja för, då må han understödja dem utan att församlingen betungas, för att denna så må kunna understödja rätta, värnlösa änkor.
Sådana äldste som äro goda församlingsföreståndare må aktas dubbel heder värda, först och främst de som arbeta med predikande och undervisning.
Skriften säger ju: »Du skall icke binda munnen till på oxen som tröskar», så ock: »Arbetaren är värd sin lön.» --
Upptag intet klagomål mot någon av de äldste, om det icke styrkes av två eller tre vittnen.
Men begår någon en synd, så skall du inför alla förehålla honom den, så att också de andra känna fruktan.
Jag uppmanar dig allvarligt inför Gud och Kristus Jesus och de utvalda änglarna att iakttaga detta, utan någon förutfattad mening och utan att i något stycke förfara partiskt.
Förhasta dig icke med handpåläggning, och gör dig icke delaktig i en annans synder.
Bevara dig själv ren.
Drick nu icke längre allenast vatten, utan bruka något litet vin för din mages skull, eftersom du så ofta lider av svaghet.
Somliga människors synder ligga i öppen dag och komma i förväg fram till dom; andras åter komma först efteråt fram.
Sammalunda pläga ock goda gärningar ligga i öppen dag; och när så icke är, kunna de ändå icke bliva fördolda.
De som äro trälar och tjäna under andra må akta sina herrar all heder värda, så att Guds namn och läran icke bliva smädade.
Men de som hava troende herrar må icke, därför att de äro deras bröder, akta dem mindre; fastmer må de tjäna dem så mycket villigare, just därför att de äro troende och kära bröder, dessa som vinnlägga sig om att göra vad gott är.
Så skall du undervisa och förmana.
Om någon förkunnar främmande läror och icke håller sig till sunda ord -- vår Herres, Jesu Kristi, ord -- och till den lära som hör gudsfruktan till,
då är han förblindad av högmod, och detta fastän han intet förstår, utan är såsom från vettet i sitt begär efter disputerande och ordstrider, vilka vålla avund, kiv, smädelser, ondskefulla misstankar
och ständiga tvister mellan människor som äro fördärvade i sitt sinne och hava tappat bort sanningen, människor som mena att gudsfruktan är ett medel till vinning.
Ja, gudsfruktan i förening med förnöjsamhet är verkligen en stor vinning.
Vi hava ju icke fört något med oss till världen, just därför att vi icke kunna föra något med oss ut därifrån.
Hava vi föda och kläder, så må vi låta oss nöja därmed.
Men de som vilja bliva rika, de råka in i frestelser och snaror och hemfalla åt många dåraktiga och skadliga begärelser, som sänka människorna ned i fördärv och undergång.
Ty penningbegäret är en rot till allt ont; och somliga hava låtit sig så drivas därav, att de hava villats bort ifrån tron och därigenom tillskyndat sig själva många kval.
Men fly sådant, du gudsmänniska, och far efter rättfärdighet, gudsfruktan, tro, kärlek, ståndaktighet, saktmod.
Kämpa trons goda kamp, sök att vinna det eviga livet, vartill du har blivit kallad, du som ock inför många vittnen har avlagt den goda bekännelsen.
Inför Gud, som giver liv åt allt, och inför Kristus Jesus, som under Pontius Pilatus vittnade med den goda bekännelsen, manar jag dig
att, själv utan fläck och tadel, hålla vad jag har bjudit, intill vår Herres, Jesu Kristi, uppenbarelse,
vilken den salige, ende härskaren skall låta oss se, när tiden är inne, han som är konungarnas konung och herrarnas herre,
han som allena har odödlighet och bor i ett ljus dit ingen kan komma, han som ingen människa har sett eller kan se.
Honom vare ära och evigt välde!
Amen.
Bjud dem som äro rika i den tidsålder som nu är att icke högmodas, och att icke sätta sitt hopp till ovissa rikedomar, utan till Gud, som rikligen giver oss allt till att njuta därav;
bjud dem att göra gott, att vara rika på goda gärningar, att vara givmilda och gärna dela med sig.
Må de så lägga av åt sig skatter som kunna bliva en god grundval för det tillkommande, så att de vinna det verkliga livet.
O Timoteus, bevara vad som har blivit dig betrott; och vänd dig bort ifrån de oandliga, tomma ord och gensägelser som komma från den falskeligen så kallade »kunskapen»,
vilken några föregiva sig äga, varför de ock hava farit vilse i fråga om tron.
Nåd vare med eder.
Paulus, genom Guds vilja Kristi Jesu apostel -- sänd enligt det löfte som gavs oss om liv, livet i Kristus Jesus --
hälsar Timoteus, sin älskade son.
Nåd, barmhärtighet och frid ifrån Gud, Fadern, och Kristus Jesus, vår Herre!
Jag tackar Gud, som jag i likhet med mina förfäder tjänar, och det med rent samvete, såsom jag ock oavlåtligen har dig i åtanke i mina böner, både natt och dag.
Och när jag kommer ihåg dina tårar, längtar jag efter att se dig, för att så bliva uppfylld av glädje,
då jag erinras om din oskrymtade tro, samma tro som förut bodde i din mormoder Lois och din moder Eunice, och som nu -- därom är jag förvissad -- jämväl bor i dig.
Fördenskull påminner jag dig att du må uppliva den nådegåva från Gud, som i följd av min handpåläggning finnes i dig.
Ty Gud har icke givit oss en försagdbetens ande, utan en kraftens och kärlekens och tuktighetens ande.
Blygs därför icke för vittnesbördet om vår Herre, ej heller för mig, hans fånge, utan bär också du ditt lidande för evangelium, genom den kraft som Gud giver,
han som har frälst oss och kallat oss med en helig kallelse, icke på grund av våra gärningar, utan efter sitt eget rådslut och sin nåd, den nåd som redan för evärdliga tider sedan gavs oss i Kristus Jesus,
men som nu har blivit uppenbar genom vår Frälsares, Kristi Jesu, uppenbarelse.
Ty han har gjort dödens makt om intet och fört liv och oförgänglighet fram i ljuset genom evangelium,
till vars förkunnare och apostel och lärare jag har blivit satt.
Fördenskull lider jag också detta, men jag blyges dock icke därför.
Ty jag vet på vem jag tror, och jag är viss om att han är mäktig att för »den dagen» bevara vad som har blivit mig betrott.
Såsom förebild i fråga om sunda ord må du, i tron och kärleken i Kristus Jesus, hava de ord som du har hört av mig.
Bevara genom den helige Ande, vilken bor i oss, det goda som har blivit dig betrott.
Det vet du, att alla i provinsen Asien hava vänt sig ifrån mig, bland dem också Fygelus och Hermogenes.
Må Herren visa barmhärtighet mot Onesiforus' hus, eftersom han ofta var mig till vederkvickelse och icke blygdes för mina kedjor;
fastmer, när han kom till Rom, sökte han efter mig med all iver, till dess han fann mig.
Ja, Herren give att han må finna barmhärtighet hos Herren på »den dagen».
Till huru stor tjänst han var i Efesus, det vet du själv bäst.
Så bliv nu du, min son, allt starkare i den nåd som är i Kristus Jesus.
Och vad du har hört av mig och fått betygat av många vittnen, det må du betro åt män som äro förtroende värda, och som kunna bliva skickliga att i sin ordning undervisa andra.
Bär ock du ditt lidande såsom en god Kristi Jesu stridsman.
Ingen som tjänar i krig låter sig insnärjas i näringsomsorger, ty han vill vara den till behag, som har tagit honom i sin sold.
Likaså, om någon deltager i en tävlingskamp, så vinner han icke segerkransen, ifall han icke kämpar efter stadgad ordning.
Åkermannen, han som gör arbetet, bör främst av alla få njuta av frukten.
Fatta rätt vad jag säger; Herren skall giva dig förstånd i allt.
Tänk på Jesus Kristus, som är uppstånden från de döda, av Davids säd, enligt det evangelium som jag förkunnar,
och i vars tjänst jag jämväl utstår lidande, ja, till och med måste bära bojor såsom en ogärningsman.
Men Guds ord bär icke bojor.
Därför uthärdar jag ståndaktigt allting för de utvaldas skull, på det att också de må vinna frälsningen i Kristus Jesus och därmed evig härlighet.
Detta är ett fast ord; ty hava vi dött med honom, så skola vi ock leva med honom;
äro vi ståndaktiga, så skola vi ock få regera med honom Men förneka vi honom, så skall ock han förneka oss;
äro vi trolösa, så står han troget fast vid sitt ord Ty han kan icke förneka sig själv.
Påminn dem om detta, och uppmana dem allvarligt inför Gud att icke befatta sig med ordstrider; ty sådana gagna till intet, utan äro allenast till fördärv för dem som höra därpå.
Sträva med all flit efter att själv kunna träda fram inför Gud såsom en som håller provet, en arbetare som icke behöver blygas, utan rätt förvaltar sanningens ord.
Men undfly oandligt och tomt prat.
Ty de som befatta sig med sådant komma att gå allt längre i ogudaktighet,
och deras tal skall fräta omkring sig såsom ett kräftsår.
Av det slaget äro Hymeneus och Filetus;
ty när dessa säga att uppståndelsen redan har skett, hava de farit vilse från sanningen, och de förvända så tron hos somliga.
Dock, Guds fasta grundval förbliver beståndande och har ett insegel med dessa ord: »Herren känner de sina», och: »Var och en som åkallar Herrens namn, han vände sig bort ifrån orättfärdighet.»
Men i ett stort hus finnas kärl icke allenast av guld och silver, utan ock av trä och lera; och somliga äro till hedersamt bruk, andra till mindre hedersamt.
Om nu någon håller sig ren och obesmittad av sådant folk, då bliver han ett kärl till hedersamt bruk, helgat, gagneligt för sin herre, tjänligt till allt vad gott är.
Fly ungdomens onda begärelser, och far efter rättfärdighet, tro och kärlek, och frid med dem som av rent hjärta åkalla Herren.
Men undvik dåraktiga och barnsliga tvistefrågor; du vet ju att de föda av sig strider.
Och en Herrens tjänare bör icke strida, utan vara mild mot alla, väl skickad att undervisa, tålig när han får lida.
Han bör med saktmod tillrättavisa de motspänstiga, i hopp att Gud till äventyrs skall förläna dem bättring, så att de komma till kunskap om sanningen,
och i hopp att de så skola bliva nyktra och därigenom befrias ur djävulens snara; ty av honom äro de fångade, så att de göra hans vilja
Men det må du veta, att i de yttersta dagarna svåra tider skola komma.
Ty människorna skola då vara själviska, penningkära, stortaliga, övermodiga, smädelystna, olydiga mot sina föräldrar, otacksamma, gudlösa,
kärlekslösa mot sina närmaste, trolösa, begivna på förtal, omåttliga, tygellösa, fientliga mot det goda,
förrädiska, besinningslösa, förblindade av högmod; de skola älska vällust mer än Gud,
de skola hava ett sken av gudsfruktan, men skola icke vilja veta av dess kraft.
Vänd dig bort ifrån sådana.
Ty till dem höra de män som innästla sig i husen och fånga svaga kvinnor, som äro tyngda av synder och drivas av allahanda begärelser,
kvinnor som alltjämt hålla på med att lära, men aldrig kunna komma till kunskap om sanningen.
Och såsom Jannes och Jambres stodo emot Moses, så stå dessa män emot sanningen; de äro människor som äro fördärvade i sitt sinne och icke hålla provet i fråga om tron.
Men de skola icke tillstädjas att gå längre, ty deras galenskap skall bliva uppenbar för alla, såsom det skedde med de männens.
Du åter har blivit min efterföljare lära, i vandel, i strävanden, i tro, tålamod, i kärlek, i ståndaktighet,
under förföljelser och lidanden, sådana som drabbade mig i Antiokia, Ikonium och Lystra.
Ja, sådana förföljelser har jag fått utstå, men ur alla har Herren frälst mig.
Så skola ock alla de, som vilja leva gudfruktigt i Kristus Jesus, få lida förföljelse.
Men onda människor och bedragare skola gå allt längre i ondska; de skola förvilla andra och själva bliva förvillade.
Men förbliv du vid det som du har lärt, och som du har fått visshet om.
Du vet ju av vilka du har lärt det,
och du känner från barndomen de heliga skrifter som kunna giva dig vishet, så att du bliver frälst genom den tro du har i Kristus Jesus.
All skrift som är ingiven av Gud är ock nyttig till undervisning, till bestraffning, till upprättelse, till fostran i rättfärdighet,
så att en gudsmänniska kan bliva fullt färdig, väl skickad till allt gott verk.
Jag uppmanar dig allvarligt inför Gud och Kristus Jesus, inför honom som skall döma levande och döda, jag uppmanar dig vid hans tillkommelse och hans rike:
Predika ordet, träd upp i tid och otid, bestraffa tillrättavisa, förmana med allt tålamod och med undervisning i alla stycken.
Ty den tid kommer, då de icke längre skola fördraga den sunda läran, utan efter sina egna begärelser skola samla åt sig lärare hoptals, alltefter som det kliar dem i öronen,
en tid då de skola vända sina öron från sanningen, och i stället vända sig till fabler.
Men du, var nykter i allting, bär ditt lidande, utför en evangelists verk, fullgör i allo vad som tillhör ditt ämbete.
Ty själv är jag nu på väg att offras, och tiden är inne, då jag skall bryta upp.
Jag har kämpat den goda kampen, jag har fullbordat mitt lopp, jag har bevarat tron.
Nu ligger rättfärdighetens segerkrans tillreds åt mig, och Herren, den rättfärdige domaren, skall giva den åt mig på »den dagen», och icke åt mig allenast, utan åt alla som hava älskat hans tillkommelse.
Låt dig angeläget vara att snart komma till mig.
Ty av kärlek till denna tidsålders väsende har Demas övergivit mig och har begivit sig till Tessalonika; Krescens har begivit sig till Galatien och Titus till Dalmatien.
Lukas är den ende som är kvar hos mig.
Tag Markus med dig hit; ty han kan i mycket vara mig till gagn och tjäna mig.
Tykikus har jag sänt till Efesus.
När du kommer, så hav med dig den mantel som jag lämnade kvar hos Karpus i Troas, så ock böckerna, först och främst pergamentskrifterna.
Alexander, smeden, har gjort mig mycket ont; Herren kommer att vedergälla honom efter hans gärningar.
Också du må taga dig till vara för honom, ty han har häftigt trätt upp emot det som vi hava talat.
Vid mitt första försvar inför rätta kom ingen mig till hjälp, utan alla övergåvo mig; må det icke bliva dem tillräknat.
Men Herren stod mig bi och gav mig kraft, för att genom mig ordet överallt skulle bliva predikat, så att alla hedningar finge höra det; och så blev jag räddad ur lejonets gap.
Ja, Herren skall rädda mig från alla ondskans tilltag och frälsa mig till sitt himmelska rike.
Honom tillhör äran i evigheternas evigheter.
Amen.
Hälsa Priska och Akvila, så ock Onesiforus' hus.
Erastus stannade kvar i Korint, men Trofimus lämnade jag sjuk efter mig i Miletus.
Låt dig angeläget vara att komma hit före vintern.
Eubulus och Pudens och Linus och Klaudia och alla bröderna hälsa dig.
Herren vare med din ande.
Nåd vare med eder.
Paulus, Guds tjänare och Jesu Kristi apostel, sänd att verka för Guds utvaldas tro och för kunskapen om den sanning som hör gudsfruktan till,
sänd, därför att det finnes ett hopp om evigt liv -- ty evigt liv har Gud, som icke kan ljuga, för evärdliga tider sedan utlovat,
och när tiden var inne, uppenbarade han sitt ord i den predikan varmed jag genom Guds, vår Frälsares, befallning blev betrodd --
jag, Paulus, hälsar Titus, min sannskyldige son på grund av gemensam tro.
Nåd och frid ifrån Gud, Fadern, och Kristus Jesus, vår Frälsare!
När jag lämnade dig kvar på Kreta, var det för att du skulle ordna vad som ännu återstod att ordna, och för att du, på det sätt som jag har ålagt dig, skulle i var särskild stad tillsätta äldste,
varhelst någon oförvitlig man funnes, en enda kvinnas man, en som hade troende barn, vilka icke vore i vanrykte för oskickligt leverne eller vore uppstudsiga.
Ty en församlingsföreståndare bör vara oförvitlig, såsom det höves en Guds förvaltare, icke självgod, icke snar till vrede, icke begiven på vin, icke våldsam, icke sniken efter slem vinning.
Han bör fastmer vara gästvänlig, nitälska för vad gott är, leva tuktigt, rättfärdigt, heligt och återhållsamt;
han bör hålla sig stadigt vid det fasta ordet, såsom han har fått lära det, så att han är mäktig både att förmana medelst den sunda läran och att vederlägga dem som säga emot.
Ty många finnas som icke vilja veta av någon myndighet, många som föra fåfängligt tal och bedraga människors sinnen; så göra i synnerhet de omskurna.
På sådana bör man tysta munnen, ty de förvilla hela hus genom att för slem vinnings skull förkunna otillbörliga läror.
En av dem, en profet av deras eget folk, har sagt: »Kreterna, lögnare jämt, äro odjur, glupska och lata.»
Och det vittnesbördet är sant.
Du skall därför strängt tillrättavisa dem, så att de bliva sunda i tron
och icke akta på judiska fabler och vad som påbjudes av människor som vända sig från sanningen.
Allt är rent för dem som äro rena; men för de orena och otrogna är intet rent, utan hos dem äro både förstånd och samvete orenade.
De säga sig känna Gud, men med sina gärningar förneka de det; ty de äro vederstyggliga och ohörsamma människor, odugliga till allt gott verk.
Du åter må tala vad som är den sunda läran värdigt.
Förmana de äldre männen att vara nyktra, att skicka sig värdigt och tuktigt, att vara sunda i tro, i kärlek, i ståndaktighet.
Förmana likaledes de äldre kvinnorna att skicka sig såsom det höves heliga kvinnor, att icke gå omkring med förtal, icke vara trälar under begäret efter vin, utan lära andra vad gott är, för att fostra dem till tuktighet.
Förmana de yngre kvinnorna att älska sina män och sina barn,
att föra en tuktig och ren vandel, att vara goda husmödrar och att underordna sig sina män, så att Guds ord icke bliver smädat.
Förmana likaledes de yngre männen att skicka sig tuktigt.
Bliv dem i allo ett föredöme i goda gärningar, och låt dem i din undervisning finna oförfalskad renhet och värdighet,
med sunt, ostraffligt tal, så att den som står oss emot måste blygas, då han nu icke har något ont att säga om oss.
Förmana tjänarna att i allt underordna sig sina herrar, att skicka sig dem till behag och icke vara gensvariga,
att icke begå någon oärlighet, utan på allt sätt visa dem redbar trohet, så att de i alla stycken bliva en prydnad för Guds, vår Frälsares, lära.
Ty Guds nåd har uppenbarats till frälsning för alla människor;
den fostrar oss till att avsäga oss all ogudaktighet och alla världsliga begärelser, och till att leva tuktigt och rättfärdigt och gudfruktigt i den tidsålder som nu är,
medan vi vänta på vårt saliga hopps fullbordan och på den store Gudens och vår Frälsares, Kristi Jesu, härlighets uppenbarelse --
hans som har utgivit sig själv för oss, till att förlossa oss från all orättfärdighet, och till att rena åt sig ett egendomsfolk, som beflitar sig om att göra vad gott är.
Så skall du tala; och du skall förmana och tillrättavisa dem med all myndighet.
Låt ingen förakta dig.
Lägg dem på minnet att de böra vara underdåniga överheten, dem som hava myndighet, att de böra visa lydnad och vara redo till allt gott verk,
att de icke må smäda någon, icke vara stridslystna, utan vara fogliga, och att de i allt skola visa sig saktmodiga mot alla människor.
Vi voro ju själva förut oförståndiga, ohörsamma och vilsefarande, vi voro trälar under allahanda begärelser och lustar, vi levde i ondska och avund, vi voro värda att avskys, och vi hatade varandra.
Men när Guds, vår Frälsares, godhet och kärlek till människorna uppenbarades,
då frälste han oss, icke på grund av rättfärdighetsgärningar som vi hade gjort, utan efter sin barmhärtighet, genom ett bad till ny födelse och förnyelse i helig ande,
som han rikligen utgöt över oss genom Jesus Kristus, vår Frälsare,
för att vi, rättfärdiggjorda genom hans nåd, skulle, såsom vårt hopp är, få evigt liv till arvedel.
Detta är ett fast ord, och jag vill att du med kraft vittnar härom, för att de som sätta tro till Gud må beflita sig om att rätt utöva goda gärningar.
Sådant är gott och gagneligt för människorna.
Men dåraktiga tvistefrågor och släktledningshistorier må du undfly, så ock trätor och strider om lagen; ty sådant är gagnlöst och fåfängligt.
En man som kommer partisöndring åstad må du visa ifrån dig, sedan du en eller två gånger har förmanat honom;
ty du vet att en sådan är förvänd och begår synd, ja, han har själv fällt domen över sig.
När jag framdeles sänder Artemas eller Tykikus till dig, låt dig då angeläget vara att komma till mig i Nikopolis, ty jag har beslutit att stanna där över vintern.
Senas, den lagkloke, och Apollos må du med all omsorg utrusta för deras resa, så att intet fattas dem.
Och må jämväl våra bröder, för att icke bliva utan frukt, lära sig att rätt utöva goda gärningar, där hjälp är av nöden.
Alla som äro här hos mig hälsa dig.
Hälsa dem som älska oss i tron.
Nåd vare med eder alla.
Paulus, Kristi Jesu fånge, och brodern Timoteus hälsa Filemon, vår älskade broder och medarbetare,
och Appfia, vår syster, och Arkippus, vår medkämpe, och den församling som kommer tillhopa i ditt hus.
Nåd vare med eder och frid ifrån Gud, vår Fader, och Herren Jesus Kristus.
Jag tackar min Gud alltid, när jag tänker på dig i mina böner,
ty jag har hört om den kärlek och den tro som du har till Herren Jesus, och som du bevisar mot alla de heliga.
Och min bön är att den tro du har gemensam med oss må visa sig verksam, i det att du fullt inser huru mycket gott vi hava i Kristus.
Ty jag har fått mycken glädje och hugnad av den kärlek varmed du, min broder, har vederkvickt de heligas hjärtan.
Därför, fastän jag med mycken frimodighet i Kristus kunde befalla dig att göra vad du nu bör göra,
beder jag dig dock hellre därom för kärlekens skull -- jag, sådan jag nu är, den gamle Paulus, han som därtill nu är en Kristi Jesu fånge;
ja, jag beder dig för min son, den som jag har fött i min fångenskap, för Onesimus,
som förut var ingalunda var dig till »till gagn», men som nu är både dig och mig till stort gagn.
Denne sänder jag här tillbaka till dig; och när jag så gör, är det såsom sände jag åstad mitt eget hjärta.
Jag hade väl själv velat behålla honom hos mig, så att han å dina vägnar kunde hava betjänat mig i den fångenskap som jag utstår för evangelii skull.
Men utan ditt samtycke ville jag intet göra, ty det goda du gjorde skulle ju icke ske såsom av tvång, utan göras av fri vilja.
När han för en liten tid blev skild från dig, skedde detta till äventyrs just för att du skulle få honom igen för alltid,
nu icke längre såsom en träl, utan såsom något vida mer än en träl: såsom en älskad broder.
Detta är han redan för mig i högsta måtto; huru mycket mer då för dig, han, din broder både efter köttet och i Herren!
Om du alltså håller mig för din medbroder, så tag emot honom såsom du skulle taga emot mig själv.
Har han gjort dig någon orätt, eller är han dig något skyldig, så för upp det på min räkning.
Jag, Paulus, skriver här med egen hand: »Jag skall själv betala det.»
Jag skulle också kunna säga: »För upp det på din räkning.»
Ty du har ju en ännu större skuld till mig, nämligen -- dig själv.
Ja, min broder, måtte jag »få gagn» av dig i Herren!
Vederkvick mitt hjärta i Kristus.
Det är därför att jag är viss om din lydaktighet som jag har skrivit detta till dig.
Och jag vet att du kommer att göra ännu mer än jag begär.
Och så tillägger jag: bered dig på att giva mig härbärge.
Jag hoppas nämligen att jag genom edra böner skall bliva skänkt åt eder.
Epafras, min medfånge i Kristus Jesus, hälsar dig;
så göra ock Markus, Aristarkus, Demas och Lukas, mina medarbetare.
Herrens, Jesu Kristi, nåd vare med eder ande.
Sedan Gud fordom många gånger och på många sätt hade talat till fäderna genom profeterna,
har han nu, på det yttersta av denna tid, talat till oss genom sin Son, som han har insatt till arvinge av allt, genom vilken han ock har skapat världen.
Och eftersom denne är hans härlighets återsken och hans väsens avbild och genom sin makts ord bär allt, har han -- sedan han hade utfört en rening från synderna -- satt sig på Majestätets högra sida i höjden.
Och han har blivit så mycket större än änglarna som det namn han har ärvt är förmer än deras.
Ty till vilken av änglarna har han någonsin sagt: »Du är min Son, jag har i dag fött dig»? eller: »Jag skall vara hans Fader, och han skall vara min Son»?
Likaså säger han, med tanke på den tid då han åter skall låta den förstfödde inträda i världen: »Och alla Guds änglar skola tillbedja honom.»
Och medan han om änglarna säger: »Han gör sina änglar till vindar och sina tjänare till eldslågor»,
säger han om Sonen: »Gud, din tron förbliver alltid och evinnerligen, och rättvisans spira är ditt rikes spira.
Du har älskat rättfärdighet och hatat orättfärdighet; därför, o Gud, har din Gud smort dig med glädjens olja mer än dina medbröder»;
så ock: »Du, Herre, lade i begynnelsen jordens grund, och himlarna äro dina händers verk;
de skola förgås, men du förbliver; de skola alla nötas ut såsom en klädnad,
och såsom en mantel skall du hoprulla dem; såsom en klädnad skola de ock bytas om.
Men du är densamme, och dina år skola icke hava någon ände.»
Och till vilken av änglarna har han någonsin sagt: »Sätt dig på min högra sida, till dess jag har lagt dina fiender dig till en fotapall»?
Äro de icke allasammans tjänsteandar, som sändas ut till tjänst för deras skull som skola få frälsning till arvedel?
Därför böra vi så mycket mer akta på det som vi hava hört, så att vi icke gå förlorade.
Ty om det ord som talades genom änglar blev beståndande, och all överträdelse och olydnad fick sin rättvisa lön,
huru skola då vi kunna undkomma, om vi icke taga vara på en sådan frälsning? -- en frälsning som ju först förkunnades genom Herren och sedan bekräftades för oss av dem som hade hört honom,
varjämte Gud själv ytterligare gav sitt vittnesbörd genom tecken och under och allahanda kraftgärningar, och genom att utdela helig ande, allt efter sin vilja.
Ty det var icke under änglars välde som han lade den tillkommande världen, den som vi tala om.
Däremot har någon någonstädes betygat och sagt: »Vad är en människa, att du tänker på henne, eller en människoson, att du låter dig vårda om honom?
En liten tid lät du honom vara ringare än änglarna, men krönte honom sedan med härlighet och ära och satte honom till herre över dina händers verk;
allt lade du under hans fötter.»
När han underlade honom allting, undantog han nämligen intet från att bliva honom underlagt -- om vi ock ännu icke se allting vara honom underlagt.
Men honom som en liten tid hade blivit gjord »ringare än änglarna», honom, Jesus, se vi för sitt dödslidandes skull hava blivit krönt med härlighet och ära, för att det genom Guds nåd skulle komma alla till godo att han smakade döden.
Ty den för vilkens skull allting är, och genom vilken allting är, honom hövdes det, att när han ville föra många sina barn till härlighet, genom lidanden fullkomna deras frälsnings hövding.
Han som helgar och de som bliva helgade hava nämligen alla en och samme Fader.
Fördenskull blyges han icke för att kalla dem bröder;
han säger ju: »Jag skall förkunna ditt namn för mina bröder, mitt i församlingen skall jag prisa dig»;
så ock: »Jag vill sätta min förtröstan till honom»; så ock: »Se här äro jag och barnen som Gud har givit mig.»
Då nu barnen hade blivit delaktiga av kött och blod, blev ock han på ett liknande sätt delaktig därav, för att han genom sin död skulle göra dens makt om intet, som hade döden i sitt våld, det är djävulen,
och göra alla dem fria, som av fruktan för döden hela sitt liv igenom hade varit hemfallna till träldom.
Ty det är ju icke änglar som han tager sig an; det är Abrahams säd som han tager sig an.
Därför måste han i allt bliva lik sina bröder, för att han skulle bliva barmhärtig och en trogen överstepräst i sin tjänst inför Gud, till att försona folkets synder.
Ty därigenom att han har lidit, i det han själv blev frestad, kan han hjälpa dem som frestas.
Därför, I helige bröder, I som haven blivit delaktiga av en himmelsk kallelse, skolen I akta på vår bekännelses apostel och överstepräst, Jesus,
huru han var trogen mot den som hade insatt honom, likasom Moses var »trogen i hela hans hus».
Ty han har blivit aktad värdig så mycket större härlighet än Moses, som uppbyggaren av ett hus åtnjuter större ära än själva huset.
Vart och ett hus bygges ju av någon, men Gud är den som har byggt allt.
Och väl var Moses »trogen i hela hans hus», såsom »tjänare», till ett vittnesbörd om vad som framdeles skulle förkunnas;
men Kristus var trogen såsom »son», en son satt över hans hus.
Och hans hus äro vi, såframt vi intill änden hålla fast vår frimodighet och vår berömmelse i hoppet.
Så säger den helige Ande: »I dag, om I fån höra hans röst,
mån I icke förhärda edra hjärtan, såsom när de förbittrade mig på frestelsens dag i öknen,
där edra fäder frestade mig och prövade mig, fastän de hade sett mina verk i fyrtio år.
Därför blev jag förtörnad på det släktet och sade: 'Alltid fara de vilse med sina hjärtan.'
Men de ville icke veta av mina vägar.
Så svor jag då i min vrede: De skola icke komma in i min vila.»
Sen därför till, mina bröder, att icke hos någon bland eder finnes ett ont otroshjärta, så att han avfaller från den levande Guden,
utan förmanen varandra alla dagar, så länge det heter »i dag», på det att ingen av eder må bliva förhärdad genom syndens makt att bedraga.
Ty vi hava blivit delaktiga av Kristus, såframt vi eljest intill änden hålla fast vår första tillförsikt.
När det nu säges: »I dag, om I fån höra hans röst, mån I icke förhärda edra hjärtan, såsom när de förbittrade mig»,
vilka voro då de som förbittrade honom, fastän de hade hört hans ord?
Var det icke alla de som under Moses hade dragit ut ur Egypten?
Och vilka voro de som han var förtörnad på i fyrtio år?
Var det icke de som hade syndat, de »vilkas kroppar föllo i öknen»?
Och vilka gällde den ed som han svor, att de »icke skulle komma in i hans vila», vilka, om icke dem som hade varit ohörsamma?
Så se vi då att det var för otros skull som de icke kunde komma ditin.
Eftersom nu ett löfte att få komma in i hans vila ännu står kvar, må vi alltså med fruktan se till, att icke någon bland eder en gång befinnes hava blivit efter på vägen.
Ty det glada budskapet hava vi mottagit såväl som de; men för dem blev det löftesord de fingo höra till intet gagn, eftersom det icke genom tron hade blivit upptaget i dem som hörde det.
Vi som hava kommit till tro, vi få ju komma in i vilan.
Det heter också: »Så svor jag då i min vrede: De skola icke komma in i min vila», och detta fastän hans verk stodo där färdiga allt ifrån den tid då världen var skapad.
Ty om den sjunde dagen heter det någonstädes så: »Och Gud vilade på sjunde dagen från alla sina verk»;
här åter heter det: »De skola icke komma in i min vila.»
Eftersom det alltså står kvar att några skola få komma in i den, och eftersom de som först mottogo det glada budskapet för sin ohörsamhets skull icke kommo ditin,
så bestämmer han genom ordet »i dag» åter en viss dag, nu då han så lång tid därefter säger hos David, såsom förut är nämnt: »I dag, om I fån höra hans röst, mån I icke förhärda edra hjärtan.»
Ty om Josua hade fört dem in i vilan, så skulle Gud icke hava talat om en annan, senare dag.
Alltså står en sabbatsvila ännu åter för Guds folk.
Ty den som har kommit in i hans vila, han har funnit vila från sina verk, likasom Gud från sina.
Så låtom oss nu med all flit sträva efter att få komma in i den vilan, för att ingen må, såsom de, falla och bliva ett varnande exempel på ohörsamhet.
Ty Guds ord är levande och kraftigt och skarpare än något tveeggat svärd, och tränger igenom, så att det åtskiljer själ och ande, märg och ben; och det är en domare över hjärtats uppsåt och tankar.
Intet skapat är fördolt för honom, utan allt ligger blottat och uppenbart för hans ögon; och inför honom skola vi göra räkenskap.
Eftersom vi nu hava en stor överstepräst, som har farit upp genom himlarna, nämligen Jesus, Guds Son, så låtom oss hålla fast vid bekännelsen.
Ty vi hava icke en sådan överstepräst som ej kan hava medlidande med våra svagheter, utan en som har varit frestad i allting, likasom vi, dock utan synd.
Låtom oss därför med frimodighet gå fram till nådens tron, för att vi må undfå barmhärtighet och finna nåd, till hjälp i rätt tid.
Ty var och en som skall bliva överstepräst uttages bland människor och tillsättes för att till människors bästa göra tjänst inför Gud, genom att frambära gåvor och offer för synder.
Och han kan hava undseende med de okunniga och vilsefarande, just därför att han själv är behäftad med svaghet
och, för denna sin svaghets skull, måste offra för sina egna synder likaväl som för folkets.
Och ingen tager sig själv denna värdighet, utan han måste, såsom Aron, kallas därtill av Gud.
Så tog sig icke heller Kristus själv äran att bliva överstepräst, utan den äran tillföll honom genom den som sade till honom: »Du är min Son, jag har i dag fött dig»,
likasom han ock på ett annat ställe säger: »Du är en präst till evig tid, efter Melkisedeks sätt.»
Och med starkt rop och tårar frambar han, under sitt kötts dagar, böner och åkallan till den som kunde frälsa honom från döden; och han blev bönhörd och tagen ur sin ångest.
Så lärde han, fastän han var »Son», lydnad genom sitt lidande;
och när han hade blivit fullkomnad, blev han, för alla dem som äro honom lydiga, upphovet till evig frälsning
och hälsades av Gud såsom överstepräst »efter Melkisedeks sätt».
Härom hava vi mycket att säga, mycket som är svårt att göra tydligt i ord, eftersom I haven blivit så tröga till att höra.
Ty fastän det kunde vara på tiden att I själva voren lärare, behöves det snarare att man nu åter undervisar eder i de allra första grunderna av Guds ord; det har kommit därhän med eder, att I behöven mjölk i stället för stadig mat.
Men om någon är sådan att han ännu måste leva av mjölk, då är han oskicklig att förstå en undervisning om rättfärdighet; han är ju ännu ett barn.
Ty den stadiga maten tillhör de fullmogna, dem som genom vanan hava sina sinnen övade till att skilja mellan gott och ont.
Låtom oss därför lämna bakom oss de första grunderna av läran om Kristus och gå framåt mot det som hör till fullkomningen; låtom oss icke åter lägga grunden med bättring från döda gärningar och med tro på Gud,
med undervisning om dop och handpåläggning, om de dödas uppståndelse och en evig dom.
Ja, detta vilja vi göra, såframt Gud eljest tillstädjer det.
Ty dem till vilka ljuset en gång har kommit, och som hava smakat den himmelska gåvan och blivit delaktiga av helig ande,
och som hava fått smaka det goda gudsordet och den tillkommande tidsålderns krafter,
men som ändå hava avfallit -- dem är det omöjligt att återföra till ny bättring, eftersom de på nytt korsfästa Guds Son åt sig och utsätta honom för bespottelse.
Det är ju så, att den jord som indricker regnet, när det titt och ofta strömmar ned däröver, och som framalstrar växter, dem till gagn för vilkas räkning den brukas, den jorden får välsignelse från Gud.
Den åter som bär törne och tistel, den är ingenting värd och är förbannelsen nära, och slutet bliver att den avbrännes med eld.
Men i fråga om eder, I älskade, äro vi vissa om vad bättre är, och vad som länder till frälsning, om vi ock nu tala på detta sätt.
Ty Gud är icke orättvis, så att han förgäter vad I haven verkat, och vilken kärlek I bevisaden mot hans namn, då I tjänaden de heliga, såsom I ännu gören.
Men vår åstundan är att var och en av eder visar samma nit att intill änden bevara full visshet i sitt hopp,
så att I icke bliven tröga, utan bliven efterföljare åt dem som genom tro och tålamod få till arvedel vad utlovat är.
Ty när Gud gav löftet åt Abraham, svor han vid sig själv -- eftersom han icke hade någon högre att svärja vid --
och sade: »Sannerligen, jag skall rikligen välsigna dig och storligen föröka dig.»
Och när denne tåligt förbidade, fick han så vad utlovat var.
Människor svärja ju vid den som är högre än de, och eden tjänar dem till bekräftelse och gör en ände på all tvist.
Därför, när Gud ville för dem som skulle få till arvedel vad löftet innebar ännu kraftigare bevisa oryggligheten av sitt rådslut, lade han därtill en ed.
Så skulle vi genom två oryggliga utsagor, i vilka Gud omöjligen kunde ljuga, undfå en kraftig uppmuntran, vi som hava sökt vår räddning i att hålla fast vid det hopp som ligger framför oss.
I det hoppet hava vi ett säkert och fast själens ankare, som når innanför förlåten,
dit Jesus, såsom vår förelöpare, har gått in för oss, i det han blev en överstepräst »efter Melkisedeks sätt, till evig tid».
Denne Melkisedek, som var konung i Salem och präst åt Gud den Högste -- han som gick Abraham till mötes, när denne var stadd på återvägen, sedan han hade slagit konungarna, och som välsignade honom,
varvid Abraham å sin sida gav honom tionde av allt; denne, som när man uttyder vad han kallas, är först och främst »rättfärdighetens konung», men därjämte ock »Salems konung», det är »fridens konung»,
denne som står där utan fader, utan moder och utan släktledning, utan begynnelse på sina dagar och utan ände på sitt liv och likställes med Guds Son -- denne förbliver en präst för beständigt.
Och sen nu huru stor han är, denne åt vilken vår stamfader Abraham gav tionde av det förnämsta bytet.
Medan de av Levi söner, som undfå prästämbetet, hava befallning att enligt lagen taga tionde av folket, det är av sina bröder, fastän dessa hava utgått från Abrahams länd,
tog denne, som icke var av deras släkt, tionde av Abraham och välsignade honom, densamme som hade fått löftena.
Nu lär ingen kunna neka att det plägar vara den ringare som mottager välsignelse av den som står högre.
Och medan det här är dödliga människor som taga tionde, är det där en som får det vittnesbördet att han förbliver levande.
Genom Abraham har på visst sätt också Levi, som tager tionde, fått giva tionde;
ty han var ännu i sin stamfaders länd, när Melkisedek gick denne till mötes.
Vore det nu så, att fullkomning kunde vinnas genom det levitiska prästadömet -- och på detta var ju folkets lagstiftning byggd -- varför hade det då behövts att en präst av annat slag, »efter Melkisedeks sätt», skulle uppstå, en som icke nämnes »efter Arons sätt»?
(Om prästadömet förändras, måste ju med nödvändighet också lagen förändras.)
Den som detta säges om hörde nämligen till en annan stam, en stam från vilken ingen har utgått, som har gjort tjänst vid altaret.
Ty det är en känd sak att han som är vår Herre har trätt fram ur Juda stam; och med avseende på den har Moses icke talat något om präster.
Och ännu mycket tydligare blir detta, då nu en präst av annat slag uppstår, lik Melkisedek däri,
att han har blivit präst icke på grund av en lag som stadgar härstamning efter köttet, utan på grund av en kraft som kommer av oförgängligt liv.
Han får nämligen det vittnesbördet: »Du är en präst till evig tid, efter Melkisedeks sätt.»
Så upphäves nu visserligen en föregående stadga, därför att den var svag och gagnlös --
eftersom lagen icke kunde åstadkomma något fullkomligt -- men ett bättre hopp sättes i stället, ett hopp genom vilket vi få nalkas Gud.
Och i så måtto som detta icke har kommit till stånd utan edlig bekräftelse -- det är nämligen så, att medan de andra hava blivit präster utan edlig bekräftelse,
har denne blivit det med sådan bekräftelse, genom den som sade till honom: »Herren har svurit och skall icke ångra sig: 'Du är en präst till evig tid'» --
i så måtto är också det förbund bättre, som har Jesus till löftesman.
Och medan de förra prästerna hava måst bliva flera, därför att de genom döden hindrades från att förbliva i sin tjänst,
har däremot denne ett oförgängligt prästadöme, eftersom han förbliver »till evig tid».
Därför kan han ock till fullo frälsa dem som genom honom komma till Gud, ty han lever alltid för att mana gott för dem.
En sådan överstepräst hövdes oss också att hava, en som vore helig, oskyldig, obesmittad, skild från syndare och upphöjd över himmelen,
en som icke var dag behövde frambära offer, såsom de andra översteprästerna, först för sina egna synder och sedan för folkets; detta gjorde han nämligen en gång för alla, när han offrade sig själv.
Ty lagen insätter till överstepräster människor som äro behäftade med svaghet, men det löftesord, som efter lagens utgivande gavs under edlig bekräftelse, insätter en »Son» som är fullkomnad »till evig tid».
Men en huvudpunkt i vad vi vilja säga är detta: Vi hava en överstepräst som sitter på högra sidan om Majestätets tron i himmelen,
för att göra tjänst i det allraheligaste, i det sannskyldiga tabernaklet, vilket Herren har upprättat, och icke någon människa.
Ty var och en som bliver överstepräst tillsättes för att frambära gåvor och offer; därför måste också denne hava något att frambära.
Om han nu vore på jorden, så vore han icke ens präst, då andra där finnas, som efter lagens bud hava att frambära gåvorna,
i det att de tjäna i den helgedom som är en avbild och en skugga av den himmelska.
Om en sådan fick ock Moses befallning genom en uppenbarelse, när han skulle förfärdiga tabernaklet. »Se till», heter det, »att du gör allt efter den mönsterbild som har blivit dig visad på berget.»
Men nu har denne fått ett så mycket förnämligare ämbete, som han är medlare för ett bättre förbund, vars ordning vilar på bättre löften.
Ty om det förra förbundet hade varit utan brist, så skulle väl plats icke hava sökts för ett annat.
Men nu förebrår Gud dem och säger: »Se, dagar skola komma, säger Herren, då jag skall sluta ett nytt förbund med Israels hus och med Juda hus;
icke ett sådant förbund som det jag gjorde med deras fäder, på den dag då jag tog dem vid handen till att föra dem ut ur Egyptens land.
Ty de förblevo icke i mitt förbund, och därför frågade icke heller jag efter dem, säger Herren.
Nej, detta är det förbund som jag skall sluta med Israels hus i kommande dagar, säger Herren: Jag skall lägga mina lagar i deras sinnen, och i deras hjärtan skall jag skriva dem, och jag skall vara deras Gud, och de skola vara mitt folk.
Då skall den ene medborgaren aldrig behöva undervisa den andre, icke den ene brodern den andre och säga: 'Lär känna Herren'; ty de skola alla känna mig, från den minste bland dem till den störste.
Ty jag skall i nåd förlåta deras missgärningar, och deras synder skall jag aldrig mer komma ihåg.»
När han säger »ett nytt förbund», har han därmed givit till känna att det förra är föråldrat; men det som föråldras och bliver gammalt, det är nära att försvinna.
Nu hade visserligen också det förra förbundet sina gudstjänststadgar och sin jordiska helgedom.
Ty i tabernaklet inrättades ett främre rum, vari stodo ljusstaken och bordet med skådebröden; och detta rum kallas »det heliga».
Men bakom den andra förlåten var ett annat rum i tabernaklet, ett som kallas »det allraheligaste»,
med ett gyllene rökelsealtare och förbundets ark, på alla sidor överdragen med guld.
I denna förvarades ett gyllene ämbar med mannat, så ock Arons stav, som hade grönskat, och därtill förbundets tavlor.
Därovanpå stodo härlighetskeruber, som överskyggde nådastolen.
Men om vart särskilt av dessa föremål är nu icke tillfälle att tala.
Så blev detta inrättat.
Och i det främre tabernakelrummet gå prästerna ständigt in och förrätta vad som hör till gudstjänsten,
men i det andra går allenast översteprästen in en gång om året, och då aldrig utan blod; och han frambär blodet för sig själv och för folkets ouppsåtliga synder.
Därmed giver den helige Ande till känna att vägen till det allraheligaste ännu icke har blivit uppenbarad, så länge det främre tabernakelrummet fortfarande äger bestånd.
Ty detta är en sinnebild som avser den nuvarande tiden, och i enlighet härmed frambäras gåvor och offer, vilka dock icke kunna fullkomna, efter samvetets krav, den som förrättar sin gudstjänst,
utan allenast äro utvärtes stadgar -- de såväl som föreskrifterna om mat och dryck och allahanda tvagningar -- stadgar pålagda intill dess tiden vore inne för en bättre ordning.
Men Kristus kom såsom överstepräst för det tillkommande goda; och genom det större och fullkomligare tabernakel som icke är gjort med händer, det är, som icke tillhör den skapelse som nu är,
gick han, icke med bockars och kalvars blod, utan med sitt eget blod, en gång för alla in i det allraheligaste och vann en evig förlossning.
Ty om redan blod av bockar och tjurar och aska av en ko, stänkt på dem som hava blivit orenade, helgar till utvärtes renhet,
huru mycket mer skall icke Kristi blod -- då han nu genom evig ande har framburit sig själv såsom ett felfritt offer åt Gud -- rena våra samveten från döda gärningar till att tjäna den levande Guden!
Så är han medlare för ett nytt förbund, på det att de som voro kallade skulle få det utlovade eviga arvet, därigenom att en led döden till förlossning ifrån överträdelserna under det förra förbundet.
Ty där ett testamente finnes, där måste det styrkas att den som har gjort testamentet är död.
Först genom döden bliver ju ett testamente giltigt, varemot det icke äger gällande kraft, så länge den som har gjort det ännu lever.
Därför har icke heller det förra förbundet blivit invigt utan blod.
Ty sedan alla buden, såsom de lyda i lagen, hade blivit av Moses kungjorda för allt folket, tog han blod av kalvar och bockar, tillika med vatten och röd ull och isop, och bestänkte såväl själva boken som allt folket
och sade: »Detta är förbundets blod, det förbunds som Gud har stadgat för eder.»
Likaledes stänkte han ock blod på tabernaklet och på alla de ting som hörde till gudstjänsten.
Så renas enligt lagen nästan allting med blod, och utan att blod utgjutes gives ingen förlåtelse.
Alltså var det nödvändigt att avbilderna av de himmelska tingen renades genom sådana medel; men de himmelska tingen själva måste renas genom bättre offer än dessa.
Ty Kristus har icke gått in i ett allraheligaste som är gjort med händer, och som allenast är en efterbildning av det sannskyldiga, utan han har gått in i själva himmelen, för att nu träda fram inför Guds ansikte, oss till godo.
Ej heller har han gått ditin, för att många gånger offra sig själv, såsom översteprästen år efter år går in i det allraheligaste, med blod som icke är hans eget.
Han hade annars måst lida många gånger allt ifrån världens begynnelse.
I stället har han uppenbarats en enda gång, nu vid tidernas ände, för att genom offret av sig själv utplåna synden.
Och såsom det är människorna förelagt att en gång dö och sedan dömas,
så skall Kristus, sedan han en gång har blivit offrad för att bära mångas synder, för andra gången, utan synd, låta sig ses av dem som bida efter honom, till frälsning.
Ty lagen innehåller en skugga av det tillkommande goda, men framställer icke tingen i deras verkliga gestalt; därför kan den aldrig genom de offer som ständigt frambäras, år efter år på samma sätt, fullkomna dem som framträda med sådana.
Annars skulle man väl hava upphört att offra, då ju de som så förrättade sin gudstjänst icke mer kunde veta med sig någon synd, sedan de en gång hade blivit renade.
Men just i offren ligger en årlig påminnelse om synd.
Ty omöjligt är att tjurars och bockars blod skulle kunna borttaga synder.
Därför säger han vid sitt inträde i världen: »Slaktoffer och spisoffer begärde du icke, men en kropp beredde du åt mig;
i brännoffer och syndoffer fann du icke behag.
Då sade jag: 'Se, jag kommer -- i bokrullen är skrivet om mig -- för att göra din vilja, o Gud.'»
Sedan han först har sagt: »Slaktoffer och spisoffer, brännoffer och syndoffer begärde du icke, och i sådana fann du icke behag» -- och dock frambäras de efter lagen --
säger han vidare: »Se, jag kommer för att göra din vilja.»
Så tager han bort det förra, för att sätta det andra i stället.
Och i kraft av denna »vilja» hava vi blivit helgade, därigenom att Jesu Kristi »kropp» en gång för alla har blivit offrad.
Och alla andra präster stå dag efter dag i sin tjänst och frambära gång på gång enahanda offer, som dock aldrig kunna borttaga synder;
men sedan denne har framburit ett enda offer för synderna, sitter han för beständigt på Guds högra sida
och väntar nu allenast på att »hans fiender skola bliva lagda honom till en fotapall».
Ty med ett enda offer har han för beständigt fullkomnat dem som bliva helgade.
Härom vittnar jämväl den helige Ande för oss.
Ty sedan Herren hade sagt:
»Detta är det förbund som jag skall sluta med dem i kommande dagar», säger han: »Jag skall lägga mina lagar i deras hjärtan, och i deras sinnen skall jag skriva dem»;
och vidare: »Deras synder och deras orättfärdiga gärningar skall jag aldrig mer komma ihåg.»
Men där förlåtelse för dessa är given, där behöves icke mer något offer för synd.
Eftersom vi nu, mina bröder, hava en fast tillförsikt att få gå in i det allraheligaste i och genom Jesu blod,
i det att han åt oss har invigt en ny och levande väg ditin genom förlåten -- det är genom sitt kött --
och eftersom vi hava en stor överstepräst över Guds hus,
så låtom oss med uppriktiga hjärtan gå fram i full trosvisshet, bestänkta till våra hjärtan och därigenom renade från ett ont samvete, och till kroppen tvagna med rent vatten.
Låtom oss oryggligt hålla fast vid hoppets bekännelse, ty den som har givit oss löftet, han är trofast.
Och låtom oss akta på varandra för att uppliva varandra till kärlek och goda gärningar;
låtom oss icke övergiva vår församlingsgemenskap, såsom somliga hava för sed, utan må vi förmana varandra -- detta så mycket mer som I sen huru »dagen» nalkas.
Ty om vi med berått mod synda, sedan vi hava undfått kunskapen om sanningen, så återstår icke mer något offer för våra synder,
utan allenast en förskräcklig väntan på dom och glöden av en eld som skall förtära motståndarna.
Den som föraktar Moses' lag, han skall »efter två eller tre vittnens utsago» dödas utan barmhärtighet;
huru mycket svårare straff tron I icke då att den skall anses värd, som förtrampar Guds Son och aktar förbundets blod för orent -- det i vilket han har blivit helgad -- och som smädar nådens Ande!
Vi veta ju vem han är som sade: »Min är hämnden; jag skall vedergälla det», och åter: »Herren skall döma sitt folk.»
Det är förskräckligt att falla i den levande Gudens händer.
Men kommen ihåg den förgångna tiden, då I, sedan ljuset hade kommit till eder, ståndaktigt uthärdaden mången lidandets kamp
och dels själva genom smälek och misshandling bleven gjorda till ett skådespel för världen, dels leden med andra som fingo genomgå sådant.
Ty I haven delat de fångnas lidanden och med glädje underkastat eder att bliva berövade edra ägodelar.
I vissten nämligen att I haven en egendom som är bättre och bliver beståndande.
Så kasten nu icke bort eder frimodighet, som ju har med sig stor lön.
I behöven nämligen ståndaktighet för att kunna göra Guds vilja och få vad utlovat är.
Ty »ännu en helt liten tid, så kommer den som skall komma, och han skall icke dröja;
och min rättfärdige skall leva av tro.
Men om någon drager sig undan, så finner min själ icke behag i honom».
Dock, vi höra icke till dem som draga sig undan, sig själva till fördärv; vi höra till dem som tro och så vinna sina själar.
Men tron är en fast tillförsikt om det som man hoppas, en övertygelse om ting som man icke ser.
På grund av den fingo ju de gamle sitt vittnesbörd.
Genom tron förstå vi att världen har blivit fullbordad genom ett ord av Gud, så att det man ser icke har blivit till av något synligt.
Genom tron frambar Abel åt Gud ett bättre offer än Kain, och genom den fick han det vittnesbördet att han var rättfärdig, i det Gud själv gav vittnesbörd om hans offergåvor; och genom tron talar han ännu, fastän han är död.
Genom tron togs Enok bort, för att han icke skulle se döden; och »man såg honom icke mer, ty Gud tog honom bort».
Förrän han togs bort, fick han nämligen det vittnesbördet att han hade täckts Gud;
men utan tro är det omöjligt att täckas Gud.
Ty den som vill komma till Gud måste tro att han är till, och att han lönar dem som söka honom.
Genom tron var det som Noa, sedan han hade fått uppenbarelse om något som man ännu icke såg, i from förtröstan byggde en ark för att rädda sitt hus; och genom den blev han världen till dom och fick till arvedel den rättfärdighet som hör tron till.
Genom tron var Abraham lydig, när han blev kallad, och han drog så ut till det land som han skulle få till arvedel; han drog ut, fastän han icke visste vart han skulle komma.
Genom tron bosatte han sig såsom främling i det utlovade landet, likasom i ett främmande land, och bodde i tält med Isak och Jakob, som voro hans medarvingar till samma löfte.
Ty han väntade på »staden med de fasta grundvalarna», vars byggmästare och skapare är Gud.
Genom tron fick jämväl Sara, fastän överårig, kraft att bliva stammoder för en avkomma, i det hon höll den för trovärdig, som hade givit löftet.
Därför föddes ock av en och samme man, en som var så gott som död, avkomlingar »så talrika som stjärnorna på himmelen och som sanden på havets strand, som man icke kan räkna».
I tron dogo alla dessa, innan de ännu hade fått vad utlovat var; de hade allenast sett det i fjärran och hade hälsat det och bekänt sig vara »gäster och främlingar» på jorden.
De som så tala giva ju därmed till känna att de söka efter ett fädernesland.
Och om de hade menat det land som de hade gått ut ifrån, så hade de haft tillfälle att vända tillbaka dit.
Men nu stod deras håg till ett bättre, nämligen det himmelska.
Därför blyges icke Gud för att kallas deras Gud; ty han har berett åt dem en stad.
Genom tron var det som Abraham frambar Isak såsom offer, när han blev satt på prov; ja, sin ende son frambar han såsom offer, han som hade mottagit löftena,
han till vilken det hade blivit sagt: »Genom Isak är det som säd skall uppkallas efter dig.»
Ty han tänkte på att Gud var mäktig att till och med uppväcka från de döda; från de döda fick han honom ock tillbaka, liknelsevis talat.
Genom tron gav jämväl Isak sin välsignelse åt Jakob och Esau för kommande tider.
Genom tron välsignade den döende Jakob Josefs båda söner och tillbad, lutad mot ändan av sin stav.
Genom tron talade Josef, när han låg för döden, om Israels barns uttåg och gav befallning om vad som skulle göras med hans ben.
Genom tron blev Moses vid sin födelse dold av sina föräldrar och hölls av dem gömd i tre månader, eftersom de sågo att »det var ett vackert barn»; och de läto icke förskräcka sig av konungens påbud.
Genom tron försmådde Moses, sedan han hade blivit stor, att kallas Faraos dotterson.
Han ville hellre utstå lidande med Guds folk än för en kort tid leva i syndig njutning;
han höll nämligen Kristi smälek för en större rikedom än Egyptens skatter, ty han hade sin blick riktad på lönen.
Genom tron övergav han Egypten, utan att låta förskräcka sig av konungens vrede; ty därigenom att han likasom såg den Osynlige kunde han härda ut.
Genom tron har han ock förordnat om påsken och blodbestrykningen, på det att »Fördärvaren», som förgjorde allt förstfött, icke skulle komma vid dem.
Genom tron drogo de fram genom Röda havet likasom på torra landet; men när egyptierna försökte gå samma väg, dränktes de.
Genom tron föllo Jerikos murar, sedan man i sju dagar hade gått runt omkring dem.
Genom tron undgick skökan Rahab att förgås tillsammans med de ohörsamma, eftersom hon hade tagit emot spejarna såsom vänner.
Och vad skall jag nu vidare säga?
Tiden bleve mig ju för kort, ifall jag skulle förtälja om Gideon, Barak, Simson och Jefta, om David och Samuel och profeterna,
om dessa som genom tron besegrade konungariken, övade rättfärdighet, fingo löften uppfyllda, tillstoppade lejons gap,
dämpade eldens kraft, undkommo svärdets egg, blevo starka från att hava varit svaga, blevo väldiga i krig och drevo främmande härar på flykten.
Kvinnor funnos som fingo igen sina döda genom deras uppståndelse.
Andra läto sig läggas på sträckbänk och ville icke taga emot någon befrielse, i hopp om en så mycket bättre uppståndelse.
Andra åter underkastade sig begabberi och gisselslag, därtill ock bojor och fängelse;
de blevo stenade, marterade, söndersågade, dödade med svärd.
De gingo omkring höljda i fårskinn och gethudar, nödställda, misshandlade, plågade,
dessa människor som världen icke var värdig att hysa; de irrade omkring i öknar och bergstrakter och levde i hålor och jordkulor.
Och fastän alla dessa genom tron hava fått sitt vittnesbörd, undfingo de ändå icke vad utlovat var;
ty Gud hade åt oss utsett något bättre, på det att de icke oss förutan skulle bliva fullkomnade.
Alltså, då vi nu hava omkring oss en så stor hop av vittnen, må ock vi lägga av allt som är oss till hinder, och särskilt synden, som så hårt omsnärjer oss, och med uthållighet löpa framåt i den tävlingskamp som är oss förelagd.
Och må vi därvid se på Jesus, trons hövding och fullkomnare, på honom, som i stället för att taga den glädje som låg framför honom, utstod korsets lidande och aktade smäleken för intet, och som nu sitter på högra sidan om Guds tron.
Ja, på honom, som har utstått så mycken gensägelse av syndare, på honom mån I tänka, så att I icke tröttnen och uppgivens i edra själar.
Ännu haven I icke stått emot ända till blods, i eder kamp mot synden.
Och I haven alldeles förgätit den förmaningens röst som talar med eder, såsom man talar med söner: »Min son, förkasta icke Herrens aga, och giv dig icke över, när du tuktas av honom.
Ty den Herren älskar, den agar han, och han straffar med riset var son som han har kär.»
Det är till eder fostran som I fån utstå lidande; Gud handlar med eder såsom med söner.
Ty var finnes den son som icke bliver agad av sin fader?
Om I lämnadens utan aga, medan alla andra finge sin del därav, så voren I oäkta söner och icke äkta.
Vidare: vi hava haft köttsliga fäder, som agade oss, och vi visade försyn för dem; skola vi då icke mycket mer vara underdåniga andarnas Fader, så att vi få leva?
De förra agade oss ju för en kort tid, såsom det syntes dem gott, men denne agar oss för vårt verkliga gagn, för att vi skola få del av hans helighet.
Väl synes alla aga för tillfället vara icke till glädje, utan till sorg; men efteråt bär den, för dem som hava blivit fostrade därmed, en fridsfrukt som är rättfärdighet.
Alltså: »stärken maktlösa händer och vacklande knän»,
och »gören räta stigar för edra fötter», så att den fot som haltar icke vrides ur led, utan fastmer bliver botad.
Faren efter frid med alla och efter helgelse; ty utan helgelse får ingen se Herren.
Och sen till, att ingen går miste om Guds nåd, och att ingen giftig rot skjuter skott och bliver till fördärv, så att menigheten därigenom bliver besmittad;
sen till, att ingen är en otuktig människa eller ohelig såsom Esau, han som för en enda maträtt sålde sin förstfödslorätt.
I veten ju att han ock sedermera blev avvisad, när han på grund av arvsrätt ville få välsignelsen; han kunde nämligen icke vinna någon ändring, fastän han med tårar sökte därefter.
Ty I haven icke kommit till ett berg som man kan taga på, ett som »brann i eld», icke till »töcken och mörker» och storm,
icke till »basunljud» och till en »röst» som talade så, att de som hörde den bådo att intet ytterligare skulle talas till dem.
Ty de kunde icke härda ut med det påbud som gavs dem: »Också om det är ett djur som kommer vid berget, skall det stenas.»
Och så förskräcklig var den syn man såg, att Moses sade: »Jag är förskräckt och bävar.»
Nej, I haven kommit till Sions berg och den levande Gudens stad, det himmelska Jerusalem, och till änglar i mångtusental,
till en högtidsskara och församling av förstfödda söner som äro uppskrivna i himmelen, och till en domare som är allas Gud, och till fullkomnade rättfärdigas andar,
och till ett nytt förbunds medlare, Jesus, och till ett stänkelseblod som talar bättre än Abels blod.
Sen till, att I icke visen ifrån eder honom som talar.
Ty om dessa icke kunde undfly, när de visade ifrån sig honom som här på jorden kungjorde Guds vilja, huru mycket mindre skola då vi kunna det, om vi vända oss ifrån honom som kungör sin vilja från himmelen?
Hans röst kom då jorden att bäva; men nu har han lovat och sagt: »Ännu en gång skall jag komma icke allenast jorden, utan ock himmelen att bäva.»
Dessa ord »ännu en gång» giva till känna att de ting, som kunna bäva, skola, eftersom de äro skapade, bliva förvandlade, för att de ting, som icke kunna bäva, skola bliva beståndande.
Därför, då vi nu skola undfå ett rike som icke kan bäva, så låtom oss vara tacksamma.
På det sättet tjäna vi Gud, honom till behag, med helig fruktan och räddhåga.
Ty »vår Gud är en förtärande eld».
Förbliven fasta i broderlig kärlek.
Förgäten icke att bevisa gästvänlighet; ty genom gästvänlighet hava några, utan att veta det, fått änglar till gäster.
Tänken på dem som äro fångna, likasom voren I deras medfångar, och tänken på dem som utstå misshandling, eftersom också I själva haven en kropp.
Äktenskapet må hållas i ära bland alla, och äkta säng bevaras obesmittad; ty otuktiga människor och äktenskapsbrytare skall Gud döma.
Varen i eder handel och vandel fria ifrån penningbegär; låten eder nöja med vad I haven.
Ty han har själv sagt: »Jag skall icke lämna dig eller övergiva dig.»
Alltså kunna vi dristigt säga: »Herren är min hjälpare, jag skall icke frukta; vad kunna människor göra mig?»
Tänken på edra lärare, som hava talat Guds ord till eder; sen huru de slutade sin levnad, och efterföljen deras tro.
Jesus Kristus är densamme i går och i dag, så ock i evighet.
Låten eder icke vilseföras av allahanda främmande läror.
Ty det är gott att bliva styrkt i sitt hjärta genom nåd och icke genom offermåltider; de som hava befattat sig med sådant hava icke haft något gagn därav.
Vi hava ett altare, från vilket de som göra tjänst vid tabernaklet icke hava rätt att få något att äta.
Det är ju så, att kropparna av de djur, vilkas blod översteprästen bär in i det allraheligaste till försoning för synd, »brännas upp utanför lägret».
Därför var det ock utanför stadsporten som Jesus utstod sitt lidande, för att han genom sitt eget blod skulle helga folket.
Låtom oss alltså gå ut till honom »utanför lägret» och bära hans smälek.
Ty vi hava här ingen varaktig stad, utan söka efter den tillkommande staden.
Så låtom oss då genom honom alltid till Gud »frambära ett lovets offer», det är »en frukt ifrån läppar» som prisa hans namn.
Men förgäten icke att göra gott och dela med eder, ty sådana offer har Gud behag till.
Varen edra lärare hörsamma, och böjen eder för dem; ty de vaka över edra själar, eftersom de skola avlägga räkenskap.
Må de då kunna göra det med glädje, och icke med suckan, ty detta vore eder icke nyttigt.
Bedjen för oss; ty vi tro oss hava ett gott samvete, eftersom vi söka att i alla stycken föra en god vandel.
Och jag uppmanar eder att göra detta, så mycket mer som jag hoppas att därigenom dess snarare bliva återgiven åt eder.
Men fridens Gud, som från de döda har återfört vår Herre Jesus, vilken genom ett evigt förbunds blod är den store herden för fåren,
han fullkomne eder i allt vad gott är, så att I gören hans vilja; och han verke i oss vad som är välbehagligt inför honom, genom Jesus Kristus.
Honom tillhör äran i evigheternas evigheter.
Amen.
Jag beder eder, mina bröder: tagen icke illa upp dessa förmaningens ord; jag har ju ock skrivit till eder helt kort.
Veten att vår broder Timoteus har blivit lösgiven.
Om han snart kommer hit, vill jag tillsammans med honom besöka eder.
Hälsen alla edra lärare och alla de heliga.
De italiska bröderna hälsa eder.
Nåd vare med eder alla.
Jakob, Guds och Herrens, Jesu Kristi, tjänare, hälsar de tolv stammar som bo kringspridda bland folken.
Mina bröder, hållen det för idel glädje, när I kommen i allahanda frestelser,
och veten, att om eder tro håller provet, så verkar detta ståndaktighet.
Och låten ståndaktigheten hava med sig fullkomlighet i gärning, så att I ären fullkomliga, utan fel och utan brist i något stycke.
Men om någon av eder brister i vishet, så må han utbedja sig sådan från Gud, som giver åt alla villigt och utan hårda ord, och den skall bliva honom given.
Men han bedje i tro, utan att tvivla; ty den som tvivlar är lik havets våg, som drives omkring av vinden och kastas hit och dit.
En sådan människa må icke tänka att hon skall få något från Herren --
en människa med delad håg, en som går ostadigt fram på alla sina vägar.
Den broder som lever i ringhet berömme sig av sin höghet.
Den åter som är rik berömme sig av sin ringhet, ty såsom gräsets blomster skall han förgås.
Solen går upp med sin brännande hetta och förtorkar gräset, och dess blomster faller av, och dess fägring förgår; så skall ock den rike förvissna mitt i sin ävlan.
Salig är den man som är ståndaktig i frestelsen; ty när han har bestått sitt prov, skall han få livets krona, vilken Gud har lovat åt dem som älska honom.
Ingen säge, när han bliver frestad, att det är från Gud som hans frestelse kommer; ty såsom Gud icke kan frestas av något ont, så frestar han icke heller någon.
Nej, närhelst någon frestas, så är det av sin egen begärelse som han drages och lockas.
Sedan, när begärelsen har blivit havande, föder hon synd, och när synden har blivit fullmogen, framföder hon död.
Faren icke vilse, mina älskade bröder.
Idel goda gåvor och idel fullkomliga skänker komma ned ovanifrån, från himlaljusens Fader, hos vilken ingen förändring äger rum och ingen växling av ljus och mörker.
Efter sitt eget beslut födde han oss till liv genom sanningens ord, för att vi skulle vara en förstling av de varelser han har skapat.
Det veten I, mina älskade bröder.
Men var människa vare snar till att höra och sen till att tala och sen till vrede.
Ty en mans vrede kommer icke åstad vad rätt är inför Gud.
Skaffen därför bort all orenhet och all ondska som finnes kvar, och mottagen med saktmod det ord som är plantat i eder, och som kan frälsa edra själar.
Men varen ordets görare, och icke allenast dess hörare, eljest bedragen I eder själva.
Ty om någon är ordets hörare, men icke dess görare, så är han lik en man som betraktar sitt ansikte i en spegel:
när han har betraktat sig däri, går han sin väg och förgäter strax hurudan han var.
Men den som skådar in i den fullkomliga lagen, frihetens lag, och förbliver därvid och icke är en glömsk hörare, utan en verklig görare, han varder salig i sin gärning.
Om någon menar sig tjäna Gud och icke tyglar sin tunga, utan bedrager sitt hjärta, så är hans gudstjänst intet värd.
En gudstjänst, som är ren och obesmittad inför Gud och Fadern, är det att vårda sig om fader- och moderlösa barn och änkor i deras bedrövelse, och att hålla sig obefläckad av världen.
Mina bröder, menen icke att tron på vår Herre Jesus Kristus, den förhärligade, kan stå tillsammans med att hava anseende till personen.
Om till exempel i eder församling inträder en man med guldring på fingret och i präktiga kläder, och jämte honom inträder en fattig man i smutsiga kläder,
och I då vänden edra blickar till den som bär de präktiga kläderna och sägen till honom: »Sitt du här på denna goda plats», men däremot sägen till den fattige: »Stå du där», eller: »Sätt dig därnere vid min fotapall» --
haven I icke då kommit i strid med eder själva och blivit domare som döma efter orätta grunder?
Hören, mina älskade bröder: Har icke Gud utvald just dem som i världens ögon äro fattiga till att bliva rika i tro, och att få till arvedel det rike han har lovat åt dem som älska honom?
I åter haven visat förakt för den fattige.
Är det då icke de rika som förtrycka eder, och är det icke just de, som draga eder inför domstolarna?
Är det icke de, som smäda det goda namn som är nämnt över eder?
Om I, såsom skriften bjuder, fullgören den konungsliga lagen: »Du skall älska din nästa såsom dig själv», då gören I visserligen väl.
Men om I haven anseende till personen, så begån I synd och bliven av lagen överbevisade om att vara överträdare.
Ty om någon håller hela lagen i övrigt, men felar i ett, så är han skyldig till allt.
Densamme som sade: »Du skall icke begå äktenskapsbrott», han sade ju ock: »Du skall icke dräpa.»
Om du nu visserligen icke begår äktenskapsbrott, men dräper, så är du dock en lagöverträdare.
Talen och handlen så, som det höves människor vilka skola dömas genom frihetens lag.
Ty domen skall utan barmhärtighet drabba den som icke har visat barmhärtighet; barmhärtighet åter kan frimodigt träda fram inför domen.
Mina bröder, vartill gagnar det, om någon säger sig hava tro, men icke har gärningar?
Icke kan väl tron frälsa honom?
Om någon, vare sig en broder eller en syster, saknade kläder och vore utan mat för dagen
och någon av eder då sade till denne: »Gå i frid, kläd dig varmt, och ät dig mätt» -- vartill gagnade detta, såframt han icke därjämte gåve honom vad hans kropp behövde?
Så är ock tron i sig själv död, om den icke har med sig gärningar.
Nu torde någon säga: »Du har ju tro?» -- »Ja, och jag har också gärningar; visa mig du din tro utan gärningar, så vill jag genom mina gärningar visa dig min tro.»
Du tror att Gud är en.
Däri gör du rätt; också de onda andarna tro det och bäva.
Men vill du då förstå, du fåkunniga människa, att tron utan gärningar är till intet gagn!
Blev icke Abraham, vår fader, rättfärdig av gärningar, när han frambar sin son Isak på altaret?
Du ser alltså att tron samverkade med hans gärningar, och av gärningarna blev tron fullkomnad,
och så fullbordades det skriftens ord som säger: »Abraham trodde Gud, och det räknades honom till rättfärdighet»; och han blev kallad »Guds vän».
I sen alltså att det är av gärningar som en människa bliver rättfärdig, och icke av tro allenast.
Och var det icke på samma sätt med skökan Rahab?
Blev icke hon rättfärdig av gärningar, när hon tog emot sändebuden och sedan på en annan väg släppte ut dem?
Ja, såsom kroppen utan ande är död, så är ock tron utan gärningar död.
Mina bröder, icke många av eder må träda upp såsom lärare; I bören veta att vi skola få en dess strängare dom.
I många stycken fela vi ju alla; om någon icke felar i sitt tal, så är denne en fullkomlig man, som förmår tygla hela sin kropp.
När vi lägga betsel i hästarnas mun, för att de skola lyda oss, då kunna vi därmed styra också hela deras övriga kropp.
Ja, till och med skeppen, som äro så stora, och som drivas av starka vindar, styras av ett helt litet roder åt det håll dit styrmannen vill.
Så är ock tungan en liten lem och kan likväl berömma sig av stora ting.
Betänken huru en liten eld kan antända en stor skog.
Också tungan är en eld; såsom en värld av orättfärdighet framstår den bland våra lemmar, tungan som befläckar hela kroppen och sätter »tillvarons hjul» i brand, likasom den själv är antänd av Gehenna.
Ty väl är det så, att alla varelsers natur, både fyrfotadjurs och fåglars och kräldjurs och vattendjurs, låter tämja sig, och verkligen har blivit tamd, genom människors natur.
Men tungan kan ingen människa tämja; ett oroligt och ont ting är den, och full av dödande gift.
Med den välsigna vi Herren och Fadern, och med den förbanna vi människorna, som äro skapade till att vara Gud lika.
Ja, från en och samma mun utgå välsignelse och förbannelse.
Så bör det icke vara, mina bröder.
Icke giver väl en källa från en och samma åder både sött och bittert vatten?
Mina bröder, icke kan väl ett fikonträd bära oliver eller ett vinträd fikon?
Lika litet kan en salt källa giva sött vatten.
Finnes bland eder någon vis och förståndig man, så må han, i visligt saktmod, genom sin goda vandel låta se de gärningar som hövas en sådan man.
Om I åter i edra hjärtan hysen bitter avund och ären genstridiga, då mån I icke förhäva eder och ljuga, i strid mot sanningen.
Sådan »vishet» kommer icke ned ovanifrån, utan är av jorden och tillhör de »själiska» människorna, ja, de onda andarna.
Ty där avund och genstridighet råda, där råder oordning och allt vad ont är.
Men den vishet som kommer ovanifrån är först och främst ren, vidare fridsam, foglig och mild, full av barmhärtighet och andra goda frukter, fri ifrån tvivel, fri ifrån skrymtan.
Och rättfärdighetens frukt kommer av en sådd i frid, dem till del som hålla frid.
Varav uppkomma strider, och varav tvister bland eder?
Månne icke av de lustar som föra krig i eder lemmar?
I ären fulla av begärelser, men haven dock intet; I dräpen och hysen avund, men kunnen dock intet vinna; och så tvisten och striden I. I haven intet, därför att I icke bedjen.
Dock, I bedjen, men I fån intet, ty I bedjen illa, nämligen för att kunna i edra lustar förslösa vad I fån.
I trolösa avfällingar, veten I då icke att världens vänskap är Guds ovänskap?
Den som vill vara världens vän, han bliver alltså Guds ovän.
Eller menen I att detta är ett tomt ord i skriften: »Med svartsjuk kärlek trängtar den Ande som han har låtit taga sin boning i oss»?
Men så mycket större är den nåd han giver; därför heter det: »Gud står emot de högmodiga, men de ödmjuka giver han nåd.»
Så varen nu Gud underdåniga, men stån emot djävulen, så skall han fly bort ifrån eder.
Nalkens Gud, så skall han nalkas eder.
Renen edra händer, I syndare, och gören edra hjärtan rena, I människor med delad håg.
Kännen edert elände och sörjen och gråten.
Edert löje vände sig i sorg och eder glädje i bedrövelse.
Ödmjuken eder inför Herren, så skall han upphöja eder.
Förtalen icke varandra, mina bröder.
Den som förtalar en broder eller dömer sin broder, han förtalar lagen och dömer lagen.
Men dömer du lagen, så är du icke en lagens görare, utan dess domare.
En är lagstiftaren och domaren, han som kan frälsa och kan förgöra.
Vem är då du som dömer din nästa?
Hören nu, I som sägen: »I dag eller i morgon vilja vi begiva oss till den och den staden, och där vilja vi uppehålla oss ett år och driva handel och skaffa oss vinning» --
I veten ju icke vad som kan ske i morgon.
Ty vad är edert liv?
En rök ären I, som synes en liten stund, men sedan försvinner.
I borden fastmera säga: »Om Herren vill, och vi får leva, skola vi göra det, eller det.»
Men nu talen I stora ord i eder förmätenhet.
All sådan stortalighet är ond.
Alltså, den som förstår att göra vad gott är, men icke gör det, för honom bliver detta till synd.
Hören nu, I rike: Gråten och jämren eder över det elände som skall komma över eder.
Eder rikedom multnar bort, och edra kläder frätas sönder av mal;
edert guld och silver förrostar, och rosten därpå skall vara eder till ett vittnesbörd och skall såsom en eld förtära edert kött.
I haven samlat eder skatter i de yttersta dagarna.
Se, den lön I haven förhållit arbetarna som hava avbärgat edra åkrar, den ropar över eder, och skördemännens rop hava kommit fram till Herren Sebaots öron.
I haven levat i kräslighet på jorden och gjort eder goda dagar; I haven gött eder av hjärtans lust »på eder slaktedag».
I haven dömt den rättfärdige skyldig och haven dräpt honom; han står eder icke emot.
Så biden nu tåligt, mina bröder, intill Herrens tillkommelse.
I sen huru åkermannen väntar på jordens dyrbara frukt och tåligt bidar efter den, till dess att den har fått höstregn och vårregn.
Ja, biden ock I tåligt, och styrken edra hjärtan; ty Herrens tillkommelse är nära.
Sucken icke mot varandra, mina bröder, på det att I icke mån bliva dömda.
Se, domaren står för dörren.
Mina bröder, tagen profeterna, som talade i Herrens namn, till edert föredöme i att uthärda lidande och visa tålamod.
Vi prisa ju dem saliga, som hava varit ståndaktiga.
Om Jobs ståndaktighet haven I hört, och I haven sett vilken utgång Herren beredde; ty Herren är nåderik och barmhärtig.
Men framför allt, mina bröder, svärjen icke, varken vid himmelen eller vid jorden, ej heller vid något annat, utan låten edert »ja» vara »ja», och edert »nej» vara »nej», så att I icke hemfallen under dom.
Får någon bland eder utstå lidande, så må han bedja.
Är någon glad, så må han sjunga lovsånger.
Är någon bland eder sjuk, må han då kalla till sig församlingens äldste; och dessa må bedja över honom och i Herrens namn smörja honom med olja.
Och trons bön skall hjälpa den sjuke, och Herren skall låta honom stå upp igen; och om han har begått synder, skall detta bliva honom förlåtet.
Bekännen alltså edra synder för varandra, och bedjen för varandra, på det att I mån bliva botade.
Mycket förmår en rättfärdig mans bön, när den bedes med kraft.
Elias var en människa, med samma natur som vi.
Han bad en bön att det icke skulle regna, och det regnade icke på jorden under tre år och sex månader;
åter bad han, och då gav himmelen regn, och jorden bar sin frukt.
Mina bröder, om någon bland eder har farit vilse från sanningen, och någon omvänder honom,
så mån I veta att den som omvänder en syndare från hans villoväg, han frälsar hans själ från döden och överskyler en myckenhet av synder.
Petrus, Jesu Kristi apostel, hälsar de utvalda främlingar som bo kringspridda i Pontus, Galatien, Kappadocien, provinsen Asien och Bitynien,
utvalda enligt Guds, Faderns, försyn, i helgelse i Anden, till lydnad och till bestänkelse med Jesu Kristi blod.
Nåd och frid föröke sig hos eder.
Lovad vare vår Herres, Jesu Kristi, Gud och Fader, som efter sin stora barmhärtighet har genom Jesu Kristi uppståndelse från de döda fött oss på nytt till ett levande hopp,
till ett oförgängligt, obesmittat och ovanskligt arv, som i himmelen är förvarat åt eder,
I som med Guds makt bliven genom tro bevarade till en frälsning som är beredd för att uppenbaras i den yttersta tiden.
Därför mån I fröjda eder, om I ock nu en liten tid, där så måste ske, liden bedrövelse under allahanda prövningar,
för att, om eder tro håller provet -- vilket är mycket mer värt än guldet, som förgås, men som dock genom eld bliver beprövat -- detta må befinnas lända eder till pris, härlighet och ära vid Jesu Kristi uppenbarelse.
Honom älsken I utan att hava sett honom; och fastän I ännu icke sen honom, tron I dock på honom och fröjden eder över honom med outsäglig och härlig glädje,
då I nu ären på väg att vinna det som är målet för eder tro, nämligen edra själars frälsning.
Angående denna frälsning hava profeter ivrigt forskat och rannsakat, de som profeterade om den nåd som skulle vederfaras eder.
De hava rannsakat för att finna vilken och hurudan tid det var som Kristi Ande i dem hänvisade till, när han förebådade de lidanden som skulle vederfaras Kristus, och den härlighet som därefter skulle följa.
Och det blev uppenbarat för dem att det icke var sig själva, utan eder, som de tjänade härmed.
Om samma ting har nu en förkunnelse kommit till eder genom de män som i helig ande, nedsänd från himmelen, hava för eder predikat evangelium; och i de tingen åstunda jämväl änglar att skåda in.
Omgjorden därför edert sinnes länder och varen nyktra; och sätten med full tillit edert hopp till den nåd som bjudes eder i och med Jesu Kristi uppenbarelse.
Då I nu haven kommit till lydnad, så följen icke de begärelser som I förut, under eder okunnighets tid, levden i,
utan bliven heliga i all eder vandel, såsom han som har kallat eder är helig.
Det är ju skrivet: »I skolen vara heliga, ty jag är helig.»
Och om I såsom Fader åkallen honom som utan anseende till personen dömer var och en efter hans gärningar, så vandren ock i fruktan under denna edert främlingsskaps tid.
I veten ju att det icke är med förgängliga ting, med silver eller guld, som I haven blivit »lösköpta» från den vandel I förden i fåfänglighet, efter fädernas sätt,
utan med Kristi dyra blod, såsom med blodet av ett felfritt lamm utan fläck.
Så var förutsett om honom före världens begynnelse; men först nu i de yttersta tiderna har han blivit uppenbarad för eder skull,
I som genom honom tron på Gud, vilken uppväckte honom från de döda och gav honom härlighet, så att eder tro nu ock kan vara ett hopp till Gud.
Renen edra själar, i lydnad för sanningen, till oskrymtad broderlig kärlek, och älsken varandra av hjärtat med uthållig kärlek,
I som ären födda på nytt, icke av någon förgänglig säd, utan av en oförgänglig: genom Guds levande ord, som förbliver.
Ty »allt kött är såsom gräs och all dess härlighet såsom gräsets blomster; gräset torkar bort, och blomstret faller av,
men Herrens ord förbliver evinnerligen».
Och det är detta ord som har blivit förkunnat för eder såsom ett glatt budskap.
Så läggen då bort all ondska och allt svek så ock skrymteri och avund och allt förtal.
Och då I nu ären nyfödda barn, så längten efter att få den andliga oförfalskade mjölken, på det att I genom den mån växa upp till frälsning,
om I annars haven »smakat att Herren är god».
Och kommen till honom, den levande stenen, som väl av människor är förkastad, men inför Gud är »utvald och dyrbar»;
och låten eder själva såsom levande stenar uppbyggas till ett andligt hus, så att I bliven ett »heligt prästerskap», som skall frambära andliga offer, vilka genom Jesus Kristus äro välbehagliga för Gud.
Det heter nämligen på ett ställe i skriften: »Se, jag lägger i Sion en utvald, dyrbar hörnsten, och den som tror på den skall icke komma på skam.»
För eder, I som tron, är stenen alltså dyrbar, men för sådana som icke tro »har den sten som byggningsmännen förkastade blivit en hörnsten»,
som är »en stötesten och en klippa till fall».
Eftersom de icke hörsamma ordet, stöta de sig; så var det ock bestämt om dem.
I åter ären »ett utvalt släkte, ett konungsligt prästerskap, ett heligt folk, ett egendomsfolk», för att I skolen förkunna hans härliga gärningar, hans som har kallat eder från mörkret till sitt underbara ljus.
I som förut »icke voren ett folk», men nu ären »ett Guds folk», I som »icke haden fått någon barmhärtighet», men nu »haven fått barmhärtighet».
Mina älskade, jag förmanar eder såsom »gäster och främlingar» att taga eder till vara för de köttsliga begärelserna, vilka föra krig mot själen.
Och fören en god vandel bland hedningarna, på det att dessa, om de i någon sak förtala eder såsom illgärningsmän, nu i stället, när de skåda edra goda gärningar, må för dessas skull prisa Gud på den dag då han söker dem.
Varen underdåniga all mänsklig ordning för Herrens skull, vare sig det är konungen, såsom den överste härskaren,
eller det är landshövdingarna, som ju äro sända av honom för att straffa dem som göra vad ont är och för att prisa dem som göra vad gott är.
Ty så är Guds vilja, att I med goda gärningar skolen stoppa munnen till på oförståndiga och fåkunniga människor.
I ären ju fria, dock icke som om I haden friheten för att därmed överskyla ondskan, utan såsom Guds tjänare.
Bevisen var man ära, älsken bröderna, »frukten Gud, ären konungen».
I tjänare, underordnen eder edra herrar med all fruktan, icke allenast de goda och milda, utan också de obilliga.
Ty det är välbehagligt för Gud, om någon, med honom för ögonen, tåligt uthärdar sina vedervärdigheter, när han får lida oförskylt.
Ty vad berömligt är däri att I bevisen tålamod, när I för edra synders skull fån uppbära hugg och slag?
Men om I bevisen tålamod, när I fån lida för goda gärningars skull, då är detta välbehaglig för Gud.
Ty därtill ären I kallade, då ju Kristus själv led för eder och efterlämnade åt eder en förebild, på det att I skullen följa honom och vandra i hans fotspår.
»Han hade ingen synd gjort, och intet svek fanns i hans mun.
När han blev smädad, smädade han icke igen, och när han led, hotade han icke, utan överlämnade sin sak åt honom som dömer rättvist.
Och »våra synder bar han» i sin kropp upp på korsets trä, för att vi skulle dö bort ifrån synderna och leva för rättfärdigheten; och »genom hans sår haven I blivit helade».
Ty I »gingen vilse såsom får», men nu haven I vänt om till edra själars herde och vårdare.
Sammalunda, i hustrur, underordnen eder edra män, för att också de män, som till äventyrs icke hörsamma ordet; må genom sina hustrurs vandel bliva vunna utan ord,
när de skåda den rena vandel som I fören i fruktan.
Eder prydnad vare icke den utvärtes prydnaden, den som består i hårflätningar och påhängda gyllene smycken eller i eder klädedräkt.
Den vare fastmer hjärtats fördolda människa, smyckad med den saktmodiga och stilla andens oförgängliga väsende; ty detta är dyrbart inför Gud.
På sådant sätt prydde sig ju ock fordom de heliga kvinnorna, de som satte sitt hopp till Gud och underordnade sig sina män.
Så var Sara lydig mot Abraham och kallade honom »herre»; och hennes barn haven I blivit, om I gören vad gott är, och icke låten eder förskräckas av något.
Sammalunda skolen I ock, I män, på förståndigt sätt leva tillsammans med edra hustrur, då ju hustrun är det svagare kärlet; och eftersom de äro edra medarvingar till livets nåd, skolen I bevisa dem all ära, på det att edra böner icke må bliva förhindrade.
Varen slutligen alla endräktiga, medlidsamma, kärleksfulla mot bröderna, barmhärtiga, ödmjuka.
Vedergällen icke ont med ont, icke smädelse med smädelse, utan tvärtom välsignen; därtill ären I ju ock kallade, att I skolen få välsignelse till arvedel.
Ty »den som vill älska livet och se goda dagar, han avhålle sin tunga från det som är ont och sina läppar från att tala svek;
han vände sig bort ifrån det som är ont, och göre vad gott är, han söke friden, och trakte därefter
Ty Herrens ögon äro vända till de rättfärdiga, och hans öron till deras bön.
Men Herrens ansikte är emot dem som göra det onda».
Och vem är den som kan göra eder något ont, om I nitälsken för det som är gott?
Skullen I än få lida för rättfärdighets skull, så ären I dock saliga. »Hysen ingen fruktan för dem, och låten eder icke förskräckas;
nej, Herren, Kristus, skolen I hålla helig i edra hjärtan.»
Och I skolen alltid vara redo att svara var och en som av eder begär skäl för det hopp som är i eder, dock med saktmod och i fruktan
och med ett gott samvete, så att de som smäda eder goda vandel i Kristus komma på skam, i fråga om det som de förtala eder för.
Ty det är bättre att lida för goda gärningar, om så skulle vara Guds vilja, än att lida för onda.
Kristus själv led ju en gång döden för synder; rättfärdig led han för orättfärdiga, på det att han skulle föra oss till Gud.
Ja, han blev dödad till köttet, men till anden blev han gjord levande.
I anden gick han gick han ock åstad och predikade för de andar som höllos i fängelse,
för sådana som fordom voro ohörsamma, när Guds långmodighet gav dem anstånd i Noas tid, då när en ark byggdes, i vilken några få -- allenast åtta personer -- blevo frälsta genom vatten.
Efter denna förebild bliven nu och I frälsta genom vatten -- nämligen genom ett dop som icke betyder att man avtvår kroppslig orenhet, utan betyder att man anropar Gud om ett gott samvete -- i kraft av Jesu Kristi uppståndelse,
hans som har farit upp till himmelen, och som nu sitter på Guds högra sida, sedan änglar och väldige och makter i andevärlden hava blivit honom underlagda.
Då nu Kristus har lidit till köttet, så väpnen ock I eder med samma sinne; ty den som har lidit till köttet har icke längre något att skaffa med synd.
Och leven sedan, under den tid som återstår eder här i köttet, icke mer efter människors onda begärelser, utan efter Guds vilja.
Ty det är nog, att I under den framfarna tiden haven gjort hedningarnas vilja och levat i lösaktighet och onda begärelser, i fylleri, vilt leverne och dryckenskap och i allahanda skamlig avgudadyrkan,
varför de ock förundra sig och smäda eder, då I nu icke löpen med till samma liderlighetens pöl.
Men de skola göra räkenskap inför honom som är redo att döma levande och döda.
Ty att evangelium blev förkunnat jämväl för döda, det skedde, för att dessa, om de än till köttet blevo dömda, såsom alla människor dömas, likväl till anden skulle få leva, så som Gud lever
Men änden på allting är nu nära.
Varen alltså besinningsfulla och nyktra, så att I kunnen bedja.
Och varen framför allt uthålliga i eder kärlek till varandra, ty »kärleken överskyler en myckenhet av synder».
Varen gästvänliga mot varandra utan knot,
och tjänen varandra, var och en med den nådegåva han har undfått, såsom goda förvaltare av Guds mångfaldiga nåd.
Om någon talar, så vare hans tal i enlighet med Guds ord, om någon har en tjänst, så sköte han den efter måttet av den kraft som Gud förlänar, så att Gud i allt bliver ärad genom Jesus Kristus.
Honom tillhör äran och väldet i evigheternas evigheter, amen.
Mina älskade, förundren eder icke över den luttringseld som är tänd bland eder, och som I till eder prövning måsten genomgå, och menen icke att därmed något förunderligt vederfares eder;
utan ju mer I fån dela Kristi lidanden, dess mer mån I glädja eder, för att I ock mån kunna glädjas och fröjda eder vid hans härlighets uppenbarelse.
Saliga ären I, om I för Kristi namns skull bliven smädade, ty härlighetens Ande, Guds Ande, vilar då över eder.
Det må nämligen icke ske, att någon av eder får lida såsom dråpare eller tjuv eller illgärningsman, eller därför att han blandar sig i vad honom icke vidkommer.
Men om någon får lida för att han är en kristen, då må han icke blygas, utan prisa Gud för detta namns skull.
Ty tiden är inne att domen skall begynna, och det på Guds hus; men om begynnelsen sker med oss, vad bliver då änden för dem som icke hörsamma Guds evangelium?
Och om den rättfärdige med knapp nöd bliver frälst, »huru skall det då gå den ogudaktige och syndaren?»
Alltså, de som efter Guds vilja få lida, de må anbefalla sina själar åt sin trofaste Skapare, allt under det att de göra vad gott är.
Till de äldste bland eder ställer jag nu denna förmaning, jag som själv är en av de äldste och en som vittnar om Kristi lidanden, och som jämväl har del i den härlighet som kommer att uppenbaras:
Varen herdar för Guds hjord, som I haven i eder vård, varen det icke av tvång, utan av fri vilja, icke för slem vinnings skull, utan med villigt hjärta.
Uppträden icke såsom herrar över edra församlingar, utan bliven föredömen för hjorden.
Då skolen I, när Överherden uppenbaras, undfå härlighetens oförvissneliga segerkrans.
Så skolen I ock, I yngre, å eder sida underordna eder de äldre.
Ikläden eder alla, i umgängelsen med varandra, ödmjukheten såsom en tjänardräkt.
Ty »Gud står emot de högmodiga, men de ödmjuka giver han nåd».
Ödmjuken eder alltså under Guds mäktiga hand, för att han må upphöja eder i sinom tid.
Och »kasten alla edra bekymmer på honom», ty han har omsorg om eder.
Varen nyktra och vaken.
Eder vedersakare, djävulen, går omkring såsom ett rytande lejon och söker vem han må uppsluka.
Stån honom emot, fasta i tron, och veten att samma lidanden vederfaras edra bröder här i världen.
Men all nåds Gud, som har kallat eder till sin eviga härlighet i Kristus, sedan I en liten tid haven lidit, han skall fullkomna, stödja, styrka och stadfästa eder.
Honom tillhör väldet i evigheternas evigheter.
Amen.
Genom Silvanus, eder trogne broder -- för en sådan håller jag honom nämligen -- har jag nu i korthet skrivit detta, för att förmana eder, och för att betyga att den nåd I stån i är Guds rätta nåd.
Församlingen i Babylon, utvald likasom eder församling, hälsar eder.
Så gör ock min son Markus.
Hälsen varandra med en kärlekens kyss.
Frid vare med eder alla som ären i Kristus.
Simon Petrus, Jesu Kristi tjänare och apostel, hälsar dem som i och genom vår Guds och Frälsarens, Jesu Kristi, rättfärdighet hava fått sig beskärd en lika dyrbar tro som vi.
Nåd och frid föröke sig hos eder, i kunskap om Gud och vår Herre Jesus Kristus.
Allt det som leder till liv och gudsfruktan har hans gudomliga makt skänkt oss, genom kunskapen om honom som har kallat oss medelst sin härlighet och underkraft.
Genom dem har han ock skänkt oss sina dyrbara och mycket stora löften, för att I skolen, i kraft av dem, bliva delaktiga av gudomlig natur och undkomma den förgängelse som i följd av den onda begärelsen råder i världen.
Vinnläggen eder just därför på allt sätt om att i eder tro bevisa dygd, i dygden kunskap,
i kunskapen återhållsamhet, i återhållsamheten ståndaktighet, i ståndaktigheten gudsfruktan,
i gudsfruktan broderlig kärlek, i den broderliga kärleken allmännelig kärlek.
Ty om detta finnes hos eder och mer och mer förökas, så tillstädjer det eder icke att vara overksamma eller utan frukt i fråga om kunskapen om vår Herre Jesus Kristus.
Den åter som icke har detta, han är blind och kan icke se; han har förgätit att han har blivit renad från sina förra synder,
Vinnläggen eder därför, mina bröder, så mycket mer om att göra eder kallelse och utkorelse fast.
Ty om I det gören, skolen I aldrig någonsin komma på fall.
Så skall inträdet i vår Herres och Frälsares, Jesu Kristi, eviga rike förlänas eder i rikligt mått.
Därför kommer jag alltid att påminna eder om detta, fastän I visserligen redan kännen det och ären befästa i den sanning som har kommit till eder.
Och jag håller det för rätt och tillbörligt, att så länge jag ännu är i denna kroppshydda, genom mina påminnelser väcka eder.
Ty jag vet att jag snart skall lämna min kroppshydda; detta har vår Herre Jesus Kristus givit till känna för mig.
Men jag vill härmed sörja för, att I också efter min bortgång städse kunnen draga eder detta till minnes.
Ty det var icke några slugt uttänkta fabler vi följde, när vi kungjorde för eder vår Herres, Jesu Kristi, makt och hans tillkommelse utan vi hade själva skådat hans härlighet.
Ty han fick ifrån Gud, fadern, ära och pris, när från det högsta Majestätet en röst kom till honom och sade: »Denne är min älskade Son, i vilken jag har funnit behag.»
Den rösten hörde vi själva komma från himmelen, när vi voro med honom på det heliga berget.
Så mycket fastare står nu också för oss det profetiska ordet; och I gören väl, om I akten därpå, såsom på ett ljus som lyser i en dyster vildmark, till dess att dagen gryr, och morgonstjärnan går upp i edra hjärtan.
Men det mån I framför allt veta, att ingen profetia i något skriftens ord kan av någon människas egen kraft utläggas.
Ty ingen profetia har någonsin framkommit av en människas vilja, utan därigenom att människor, drivna av den helige Ande, talade vad som gavs dem från Gud.
Men också falska profeter uppstodo bland folket, likasom jämväl bland eder falska lärare skola komma att finnas, vilka på smygvägar skola införa fördärvliga partimeningar och draga över sig själva plötsligt fördärv, i det att de till och med förneka den Herre som har köpt dem.
De skola få många efterföljare i sin lösaktighet, och för deras skull skall sanningens väg bliva smädad.
I sin girighet skola de ock med bedrägliga ord bereda sig vinning av eder.
Men sedan länge är deras dom i annalkande, den dröjer icke, och deras fördärv sover icke.
Ty Gud skonade ju icke de änglar som syndade, utan störtade dem ned i avgrunden och överlämnade dem åt mörkrets hålor, för att där förvaras till domen.
Ej heller skonade han den forntida världen, om han ock, när han lät floden komma över de ogudaktigas värld, bevarade Noa såsom rättfärdighetens förkunnare, jämte sju andra.
Och städerna Sodom och Gomorra lade han i aska och dömde dem till att omstörtas; han gjorde dem så till ett varnande exempel för kommande tiders ogudaktiga människor.
Men han frälste den rättfärdige Lot, som svårt pinades av de gudlösa människornas lösaktiga vandel.
Ty genom de ogärningar som han, den rättfärdige mannen, måste se och höra, där han bodde ibland dem, plågades han dag efter dag i sin rättfärdiga själ.
Så förstår Herren att frälsa de gudfruktiga ur prövningen, men ock att under straff förvara de orättfärdiga till domens dag.
Och detta gör han först och främst med dem som i oren begärelse stå efter köttslig lust och förakta andevärldens herrar.
I sitt trots och sin självgodhet bäva dessa människor icke för att smäda andevärldens härlige,
under det att änglar som stå ännu högre i starkhet och makt icke om dem uttala någon smädande dom inför Herren.
Men på samma sätt som oskäliga djur förgås, varelser som av naturen äro födda till att fångas och förgås, på samma sätt skola ock dessa förgås, eftersom de smäda vad de icke känna till;
och de skola så bliva bedragna på den lön som de vilja vinna genom orättfärdighet.
De hava sin lust i kräsligt leverne mitt på ljusa dagen.
De äro skamfläckar och styggelser, där de vid gästabuden, som de få hålla med eder, frossa i sina njutningar.
Deras ögon äro fulla av otuktigt begär och kunna icke få nog av synd.
De locka till sig obefästa själar.
De hava hjärtan övade i girighet.
Förbannade äro de.
De hava övergivit den raka vägen och kommit vilse genom att efterfölja Balaam, Beors son, på hans väg.
Denne åtrådde ju att vinna lön genom orättfärdighet;
men han blev tillrättavisad för sin överträdelse: en stum arbetsåsninna begynte tala med människoröst och hindrade profeten i hans galenskap.
Dessa människor äro källor utan vatten, skyar som drivas av stormvinden, och det svarta mörkret är förvarat åt dem.
Ty de tala stora ord som äro idel fåfänglighet; och då de nu själva leva i köttsliga begärelser, locka de genom sin lösaktighet till sig människor som med knapp nöd rädda sig undan sådana som vandra i villfarelse.
De lova dem frihet, fastän de själva äro förgängelsens trälar; ty den som har låtit sig övervinnas av någon, han har blivit dennes träl.
Och då de genom kunskapen om Herren och Frälsaren, Jesus Kristus, hava undkommit världens besmittelser, men sedan åter låta sig insnärjas och övervinnas av dem, så har det sista för dem blivit värre än det första.
Ty det hade varit bättre för dem att icke hava lärt känna rättfärdighetens väg, än att nu, sedan de hava lärt känna den, vända tillbaka, bort ifrån det heliga bud som har blivit dem meddelat.
Det har gått med dem såsom det riktigt heter i ordspråket: »En hund vänder åter till sina spyor», och: »Ett tvaget svin vältrar sig åter i smutsen.»
Detta är nu redan det andra brevet som jag skriver till eder, mina älskade; och i båda har jag genom mina påminnelser velat uppväcka edert rena sinne,
så att I kommen ihåg vad som har blivit förutsagt av de heliga profeterna, så ock det bud som av edra apostlar har blivit eder givet från Herren och Frälsaren.
Och det mån I framför allt veta, att i de yttersta dagarna bespottare skola komma med bespottande ord, människor som vandra efter sina egna begärelser.
De skola säga: »Huru går det med löftet om hans tillkommelse?
Från den dag då våra fäder avsomnade har ju allt förblivit sig likt, ända ifrån världens begynnelse.»
Ty när de vilja påstå detta, förgäta de att i kraft av Guds ord himlar funnos till från uråldrig tid, så ock en jord som hade kommit till av vatten och genom vatten;
och genom översvämning av vatten från dem förgicks också den värld som då fanns.
Men de himlar och den jord som nu finnas, de hava i kraft av samma ord blivit sparade åt eld, och de förvaras nu till domens dag, då de ogudaktiga människorna skola förgås.
Men ett vare icke fördolt för eder, mina älskade, detta, att »en dag är för Herren såsom tusen år, och tusen år såsom en dag».
Herren fördröjer icke uppfyllelsen av sitt löfte, såsom somliga mena att han fördröjer sig.
Men han är långmodig mot eder, eftersom han icke vill att någon skall förgås, utan att alla skola vända sig till bättring.
Men Herrens dag skall komma såsom en tjuv, och då skola himlarna med dånande hast förgås, och himlakropparna upplösas av hetta, och jorden och de verk som äro därpå brännas upp.
Eftersom nu allt detta sålunda går till sin upplösning, hurudana bören icke I då vara i helig vandel och gudsfruktan,
medan I förbiden och påskynden Guds dags tillkommelse, varigenom himlar skola upplösas av eld, och himlakroppar smälta av hetta!
Men »nya himlar och en ny jord», där rättfärdighet bor, förbida vi efter hans löfte.
Därför, mina älskade, eftersom I förbiden detta, skolen I med all flit sörja för, att I mån för honom befinnas vara obefläckade och ostraffliga, i frid.
Och I skolen hålla före, att vår Herres långmodighet länder till frälsning; såsom ock vår älskade broder Paulus har skrivit till eder efter den vishet som har blivit honom given.
Så gör han i alla sina brev, när han i dem talar om sådant, fastän visserligen i dem finnes ett och annat som är svårt att förstå, och som okunniga och obefästa människor vrångt uttyda, såsom de ock göra med de övriga skrifterna, sig själva till fördärv.
Då I nu således, mina älskade, haven fått veta detta i förväg, så tagen eder till vara för att bliva indragna i de gudlösas villfarelse och därigenom förlora edert fäste.
Växen i stället till i nåd och i kunskap om vår Herre och Frälsare, Jesus Kristus.
Honom tillhör äran, nu och till evighetens dag.
Amen.
Det som var från begynnelsen, det vi hava hört, det vi med egna ögon hava sett, det vi skådade och med egna händer togo på, det förkunna vi: om livets Ord tala vi.
Ty livet uppenbarades, och vi hava sett det; och vi vittna därom och förkunna för eder livet, det eviga, som var hos Fadern och uppenbarades för oss.
Ja, det vi hava sett och hört, det förkunna vi ock för eder, på det att också I mån hava gemenskap med oss; och vi hava vår gemenskap med Fadern och med hans Son, Jesus Kristus.
Och vi skriva nu detta, för att vår glädje skall bliva fullkomlig.
Och detta är det budskap som vi hava hört från honom, och som vi förkunna för eder, att Gud är ljus, och att intet mörker finnes i honom.
Om vi säga oss hava gemenskap med honom, och vi vandra i mörkret, så ljuga vi och göra icke sanningen.
Men om vi vandra i ljuset, såsom han är i ljuset, så hava vi gemenskap med varandra, och Jesu, hans Sons, blod renar oss från all synd.
Om vi säga att vi icke hava någon synd, så bedraga vi oss själva, och sanningen är icke i oss.
Om vi bekänna våra synder, så är han trofast och rättfärdig, så att han förlåter oss våra synder och renar oss från all orättfärdighet.
Om vi säga att vi icke hava syndat, så göra vi honom till en ljugare, och hans ord är icke i oss.
Mina kära barn, detta skriver jag till eder, för att I icke skolen synda.
Men om någon syndar, så hava vi en förespråkare hos Fadern, Jesus Kristus, som är rättfärdig;
och han är försoningen för våra synder, ja, icke allenast för våra, utan ock för hela världens.
Därav veta vi att vi hava lärt känna honom, därav att vi hålla hans bud.
Den som säger sig hava lärt känna honom och icke håller hans bud, han är en lögnare och i honom är icke sanningen.
Men den som håller hans ord, i honom är förvisso Guds kärlek fullkomnad.
Därav veta vi att vi äro i honom.
Den som säger sig förbliva i honom, han är ock pliktig att själv så vandra som Han vandrade.
Mina älskade, det är icke ett nytt bud jag skriver till eder, utan ett gammalt bud, som I haven haft från begynnelsen.
Detta gamla bud är ordet som I haven fått höra.
På samma gång är det dock ett nytt bud som jag skriver till eder.
Och detta är sant både i fråga om honom och i fråga om eder; ty mörkret förgår, och det sanna ljuset lyser redan.
Den som säger sig vara i ljuset och hatar sin broder, han är ännu alltjämt i mörkret.
Den som älskar sin broder, han förbliver i ljuset, och i honom är intet som länder till fall.
Men den som hatar sin broder, han är i mörkret och vandrar i mörkret, och han vet icke vart han går; ty mörkret har förblindat hans ögon.
Jag skriver till eder, kära barn, ty synderna äro eder förlåtna för hans namns skull.
Jag skriver till eder, I fäder, ty I haven lärt känna honom som är från begynnelsen.
Jag skriver till eder, I ynglingar, ty I haven övervunnit den onde.
Jag har skrivit till eder, mina barn, ty I haven lärt känna Fadern.
Jag har skrivit till eder, I fäder, ty I haven lärt känna honom som är från begynnelsen.
Jag har skrivit till eder, I ynglingar, ty I ären starka, och Guds ord förbliver i eder, och I haven övervunnit den onde.
Älsken icke världen, ej heller vad som är i världen.
Om någon älskar världen, så är Faderns kärlek icke i honom.
Ty allt som är i världen, köttets begärelse och ögonens begärelse och högfärd över detta livets goda, det är icke av Fadern, utan av världen.
Och världen förgår och dess begärelse, men den som gör Guds vilja, han förbliver evinnerligen.
Mina barn, nu är den yttersta tiden.
I haven ju hört att en antikrist skall komma, och redan hava många antikrister uppstått; därav förstå vi att den yttersta tiden är inne.
Från oss hava de utgått, men de hörde icke till oss, ty hade de hört till oss, så hade de förblivit hos oss.
Men det skulle bliva uppenbart att icke alla höra till oss.
I åter haven mottagit smörjelse från den Helige, och I haven all kunskap.
Jag har skrivit till eder, icke därför att I icke kännen sanningen, utan därför att I kännen den och veten att ingen lögn kommer av sanningen.
Vilken är »Lögnaren», om icke den som förnekar att Jesus är Kristus?
Denne är Antikrist, denne som förnekar Fadern och Sonen.
Var och en som förnekar Sonen, han har icke heller Fadern; den som bekänner Sonen, han har ock Fadern.
I åter skolen låta det som I haven hört från begynnelsen förbliva i eder.
Om det som I haven hört från begynnelsen förbliver i eder så skolen ock I själva förbliva i Sonen och i Fadern.
Och detta är vad han själv har lovat oss: det eviga livet.
Detta har jag skrivit till eder med tanke på dem som söka förvilla eder.
Men vad eder angår, så förbliver i eder den smörjelse I haven undfått från honom, och det behöves icke att någon undervisar eder; ty vad hans smörjelse lär eder om allting, det är sant och är icke lögn.
Förbliven alltså i honom, såsom den har lärt eder.
Ja, kära barn, förbliven nu i honom, så att vi, när han en gång uppenbaras, kunna frimodigt träda fram, och icke med skam nödgas gå bort ifrån honom vid hans tillkommelse.
Om I veten att han är rättfärdig, så kunnen I förstå att också var och en som gör vad rättfärdigt är, han är född av honom.
Se vilken kärlek Fadern har bevisat oss därmed att vi få kallas Guds barn, vilket vi ock äro.
Därför känner världen oss icke, eftersom den icke har lärt känna honom.
Mina älskade, vi äro nu Guds barn, och vad vi skola bliva, det är ännu icke uppenbart.
Men det veta vi, att när han en gång uppenbaras, skola vi bliva honom lika; ty då skola vi få se honom sådan han är.
Och var och en som har detta hopp till honom, han renar sig, likasom Han är ren.
Var och en som gör synd, han överträder ock lagen, ty synd är överträdelse av lagen.
Och i veten att Han uppenbarades, för att han skulle borttaga synderna; och synd finnes icke i honom.
Var och en som förbliver i honom, han syndar icke; var och en som syndar, han har icke sett honom och icke lärt känna honom.
Kära barn, låten ingen förvilla eder.
Den som gör vad rättfärdigt är, han är rättfärdig, likasom Han är rättfärdig.
Den som gör synd, han är av djävulen, ty djävulen har syndat från begynnelsen.
Och just därför uppenbarades Guds Son, att han skulle göra om intet djävulens gärningar.
Var och en som är född av Gud, han gör icke synd, ty Guds säd förbliver i honom; han kan icke synda, eftersom han är född av Gud.
Därav är uppenbart vilka som äro Guds barn, och vilka som äro djävulens barn, därav att var och en som icke gör vad rättfärdigt är, han är icke av Gud, ej heller den som icke älskar sin broder.
Ty detta är det budskap som I haven hört från begynnelsen, att vi skola älska varandra
och icke likna Kain, som var av den onde och slog ihjäl sin broder.
Och varför slog han ihjäl honom?
Därför att hans egna gärningar voro onda och hans broders gärningar rättfärdiga.
Förundren eder icke, mina bröder, om världen hatar eder.
Vi veta att vi hava övergått från döden till livet, ty vi älska bröderna.
Den som icke älskar, han förbliver i döden.
Var och en som hatar sin broder, han är en mandråpare; och I veten att ingen mandråpare har evigt liv förblivande i sig.
Därav att Han gav sitt liv för oss hava vi lärt känna kärleken; så äro ock vi pliktiga att giva våra liv för bröderna.
Men om någon har denna världens goda och tillsluter sitt hjärta för sin broder, när han ser honom lida nöd, huru kan då Guds kärlek förbliva i honom?
Kära barn, låtom oss älska icke med ord eller med tungan, utan i gärning och i sanning.
Därav skola vi veta att vi äro av sanningen; och så kunna vi inför honom övertyga vårt hjärta därom,
att om vårt hjärta fördömer oss, så är Gud större än vårt hjärta och vet allt.
Mina älskade, om vårt hjärta icke fördömer oss, så hava vi frimodighet inför Gud,
och vadhelst vi bedja om, det få vi av honom, eftersom vi hålla hans bud och göra vad som är välbehagligt för honom.
Och detta är hans bud, att vi skola tro på hans Sons, Jesu Kristi, namn och älska varandra, enligt det bud han har givit oss.
Och den som håller hans bud, han förbliver i Gud, och Gud förbliver i honom.
Och att han förbliver i oss, det veta vi av Anden, som han har givit oss.
Mina älskade, tron icke var och en ande, utan pröven andarna, huruvida de äro av Gud; ty många falska profeter hava gått ut i världen.
Därpå skolen I känna igen Guds Ande: var och en ande som bekänner att Jesus är Kristus, kommen i köttet, han är av Gud;
men var och en ande som icke så bekänner Jesus, han är icke av Gud.
Den anden är Antikrists ande, om vilken I haven hört att den skulle komma, och som redan nu är i världen.
I, kära barn, I ären av Gud och haven övervunnit dessa; ty han som är i eder är större än den som är i världen.
De äro av världen; därför tala de vad som är av världen, och världen lyssnar till dem.
Vi åter äro av Gud.
Den som känner Gud, han lyssnar till oss; den som icke är av Gud, han lyssnar icke till oss.
Härpå känna vi igen sanningens Ande och villfarelsens ande.
Mina älskade, låtom oss älska varandra; ty kärleken är av Gud, och var och en som älskar, han är född av Gud och känner Gud.
Den som icke älskar, han har icke lärt känna Gud, ty Gud är kärleken.
Därigenom har Guds kärlek blivit uppenbarad bland oss, att Gud har sänt sin enfödde Son i världen, för att vi skola leva genom honom.
Icke däri består kärleken, att vi hava älskat Gud, utan däri, att han har älskat oss och sänt sin Son till försoning för våra synder.
Mina älskade, om Gud så har älskat oss, då äro ock vi pliktiga att älska varandra.
Ingen har någonsin sett Gud.
Om vi älska varandra, så förbliver Gud i oss, och hans kärlek är fullkomnad i oss.
Därav att han har givit oss av sin Ande veta vi att vi förbliva i honom, och att han förbliver i oss.
Och vi hava själva sett, och vi vittna om att Fadern har sänt sin Son till att vara världens Frälsare.
Den som bekänner att Jesus är Guds Son, i honom förbliver Gud, och han själv förbliver i Gud.
Och vi hava lärt känna den kärlek som Gud har i oss, och vi hava kommit till tro på den.
Gud är kärleken, och den som förbliver i kärleken, han förbliver i Gud, och Gud förbliver i honom.
Därigenom är kärleken fullkomnad hos oss, att vi hava frimodighet i fråga om domens dag; ty sådan Han är, sådana äro ock vi i denna världen.
Räddhåga finnes icke i kärleken, utan fullkomlig kärlek driver ut räddhågan, ty i räddhågan ligger tanke på straff, och den som rädes är icke fullkomnad i kärleken.
Vi älska, därför att han först har älskat oss.
Om någon säger sig älska Gud och hatar sin broder, så är han en lögnare.
Ty den som icke älskar sin broder, som han har sett, han kan icke älska Gud, som han icke har sett.
Och det budet hava vi från honom, att den som älskar Gud, han skall ock älska sin broder.
Var och en som tror att Jesus är Kristus, han är född av Gud; och var och en som älskar honom som födde, han älskar ock den som är född av honom.
Därför, när vi älska Gud och hålla hans bud, då veta vi att vi älska Guds barn.
Ty däri består kärleken till Gud, att vi hålla hans bud; och hans bud äro icke tunga.
Ty allt som är fött av Gud, det övervinner världen; och detta är den seger som har övervunnit världen: vår tro.
Vilken annan kan övervinna världen, än den som tror att Jesus är Guds Son?
Han är den som kom genom vatten och blod, Jesus Kristus, icke med vattnet allenast, utan med vattnet och blodet.
Och Anden är den som vittnar, eftersom Anden är sanningen.
Ty tre äro de som vittna:
Anden, vattnet och blodet; och de tre vittna ett och detsamma.
Om vi taga människors vittnesbörd för gott, så må väl Guds vittnesbörd vara förmer.
Detta är ju Guds vittnesbörd, att han har vittnat om sin Son.
Den som tror på Guds Son, han har vittnesbördet inom sig själv; den som icke tror Gud, han har gjort honom till en ljugare, eftersom han icke har trott på Guds vittnesbörd om sin Son.
Och detta är vittnesbördet: att Gud har givit oss evigt liv; och det livet är i hans Son.
Den som har Sonen, han har livet; den som icke har Guds Son, han har icke livet.
Detta har jag skrivit till eder, för att I skolen veta att I haven evigt liv, I som tron på Guds Sons namn.
Och detta är den fasta tillförsikt vi hava till honom, att om vi bedja om något efter hans vilja, så hör han oss.
Och om vi veta att han hör oss, vadhelst vi bedja om, så veta vi ock att vi redan hava det som vi hava bett honom om i vår bön.
Om någon ser sin broder begå en synd som icke är en synd till döds, då må han bedja, och så skall han giva honom liv, om nämligen synden icke är till döds.
Det finnes synd till döds; för sådan säger jag icke att man skall bedja.
All orättfärdighet är synd; dock finnes det synd som icke är till döds.
Vi veta om var och en som är född av Gud att han icke syndar, ty den som har blivit född av Gud, han tager sig till vara, och den onde kommer icke vid honom.
Vi veta att vi äro av Gud, och att hela världen är i den ondes våld.
Och vi veta att Guds Son har kommit och givit oss förstånd, så att vi kunna känna den Sanne; och vi äro i den Sanne, i hans Son, Jesus Kristus.
Denne är den sanne Guden och evigt liv.
Kära barn, tagen eder till vara för avgudarna.
Den äldste hälsar den utvalda frun och hennes barn, vilka jag i sanning älskar, och icke jag allenast, utan ock alla andra som hava lärt känna sanningen.
Vi älska dem för sanningens skull, som förbliver i oss, och som skall vara med oss till evig tid.
Nåd, barmhärtighet och frid ifrån Gud, Fadern, och ifrån Jesus Kristus, Faderns Son, skall vara med oss i sanning och i kärlek.
Det har gjort mig stor glädje att jag har funnit flera av dina barn vandra i sanningen, efter det bud som vi hava fått ifrån Fadern.
Och nu har jag en bön till dig, kära fru.
Icke som om jag skreve för att giva dig ett nytt bud; det gäller allenast det bud som vi hava haft från begynnelsen: att vi skola älska varandra.
Och däri består kärleken, att vi vandra efter de bud han har givit.
Ja, detta är budet, att I skolen vandra i kärleken, enligt vad I haven hört från begynnelsen.
Ty många villolärare hava gått ut i världen, vilka icke bekänna att Jesus är Kristus, som skulle komma i köttet; en sådan är Villoläraren och Antikrist.
Tagen eder till vara, så att I icke förloren det som vi med vårt arbete hava kommit åstad, utan fån full lön.
Var och en som så går framåt, att han icke förbliver i Kristi lära, han har icke Gud; den som förbliver i den läran, han har både Fadern och Sonen.
Om någon kommer till eder och icke har den läran med sig, så tagen icke emot honom i edra hus, och hälsen honom icke.
Ty den som hälsar honom, han gör sig delaktig i hans onda gärningar.
Jag hade väl mycket annat att skriva till eder, men jag vill icke göra det med papper och bläck.
Jag hoppas att i stället få komma till eder och muntligen tala med eder, för att vår glädje skall bliva fullkomlig.
Din utvalda systers barn hälsa dig.
Den äldste hälsar Gajus, den älskade brodern, som jag i sanning älskar.
Min älskade, jag önskar att det i allt må stå väl till med dig, och att du må vara vid god hälsa, såsom det ock står väl till med din själ.
Ty det gjorde mig stor glädje, då några av bröderna kommo och vittnade om den sanning som bor i dig, eftersom du ju vandrar i sanningen.
Jag har ingen större glädje än den att få höra att mina barn vandra i sanningen.
Min älskade, du handlar såsom en trofast man i allt vad du gör mot bröderna, och detta jämväl när de komma såsom främlingar.
Dessa hava nu inför församlingen vittnat om din kärlek.
Och du gör väl, om du på ett sätt som är värdigt Gud utrustar dem också för fortsättningen av deras resa.
Ty för hans namns skull hava de dragit åstad, utan att hava tagit emot något av hedningarna.
Därför äro vi å vår sida pliktiga att taga oss an sådana män, så att vi bliva deras medarbetare till att främja sanningen.
Jag har skrivit till församlingen, men Diotrefes, som önskar att vara den främste bland dem, vill icke göra något för oss.
Om jag kommer, skall jag därför påvisa huru illa han gör, då han skvallrar om oss med elaka ord.
Och han nöjer sig icke härmed; utom det att han själv intet vill göra för bröderna, hindrar han också andra som vore villiga att göra något, ja, han driver dem ut ur församlingen.
Mina älskade, följ icke onda föredömen, utan goda.
Den som gör vad gott är, han är av Gud; den som gör vad ont är, han har icke sett Gud.
Demetrius har fått gott vittnesbörd om sig av alla, ja, av sanningen själv.
Också vi giva honom vårt vittnesbörd; och du vet att vårt vittnesbörd är sant.
Jag hade väl mycket annat att skriva till dig, men jag vill icke skriva till dig med bläck och penna.
Ty jag hoppas att rätt snart få se dig, och då skola vi muntligen tala med varandra.
Frid vare med dig.
Vännerna hälsa dig.
Hälsa vännerna, var och en särskilt.
Judas, Jesu Kristi tjänare och Jakobs broder, hälsar de kallade, dem som äro upptagna i Guds, Faderns, kärlek och bevarade åt Jesus Kristus.
Barmhärtighet och frid och kärlek föröke sig hos eder.
Mina älskade, då jag nu med all iver har tagit mig för att skriva till eder om vår gemensamma frälsning, finner jag det nödigt att i min skrivelse förmana eder att kämpa för den tro som en gång för alla har blivit meddelad åt de heliga.
Några människor hava nämligen innästlat sig hos eder -- några om vilka det för länge sedan blev skrivet att de skulle hemfalla under den domen -- ogudaktiga människor, som missbruka vår Guds nåd till lösaktighet och förneka vår ende härskare och herre, Jesus Kristus.
Men fastän I redan en gång haven fått kunskap om alltsammans, vill jag påminna eder därom, att Herren, sedan han hade frälst sitt folk ur Egyptens land, efteråt förgjorde dem som icke trodde,
så ock därom, att de änglar som icke behöllo sin furstehöghet, utan övergåvo sin boning, hava av honom med eviga bojor blivit förvarade i mörker till den stora dagens dom.
Likaså hava ock Sodom och Gomorra med kringliggande städer, vilka på samma sätt som de förra bedrevo otukt och stodo efter annat umgänge än det naturliga, blivit satta till ett varnande exempel, i det att de få lida straff i evig eld.
Dock göra nu också dessa människor på samma sätt, förblindade av sina drömmar: köttet besmitta de, men andevärldens herrar förakta de, och dess härlige smäda de.
Icke så Mikael, överängeln; när denne tvistade med djävulen angående Moses' kropp, dristade han sig icke att över honom uttala någon smädande dom, utan sade allenast: »Herren näpse dig.»
Dessa åter smäda vad de icke känna till; och vad de, likasom de oskäliga djuren, med sina naturliga sinnen kunna fatta, det bruka de till sitt fördärv.
Ve dem!
De hava trätt in på Kains väg, de hava för löns skull störtat sig i Balaams villfarelse och hava gått förlorade till följd av en gensträvighet lik Koras.
Det är dessa som få hålla gästabud med eder, där de sitta såsom skamfläckar vid edra kärleksmåltider och oförsynt se sig själva till godo.
De äro skyar utan vatten, skyar som drivas bort av vindarna.
De äro träd som stå nakna på senhösten, ofruktbara, i dubbel måtto döda, uppryckta med rötterna.
De äro vilda havsvågor som uppkasta sina egna skändligheters skum.
De äro irrande stjärnor, åt vilka det svarta mörkret är förvarat till evig tid.
Om dessa var det ock som Enok, den sjunde från Adam, profeterade och sade: »Se, Herren kommer med sina mångtusen heliga,
för att hålla dom över alla och bestraffa alla de ogudaktiga för alla de ogudaktiga gärningar som de hava övat, och för alla de förmätna ord som de i sin syndiga ogudaktighet hava talat mot honom.»
De äro människor som alltid knorra och knota över sin lott, medan de likväl vandra efter sina egna begärelser.
Och deras mun talar stora ord, under det att de dock av egennytta söka vara människor till behag.
Men kommen ihåg, I mina älskade, vad som har blivit förutsagt av vår Herres, Jesu Kristi, apostlar,
huru de sade till eder: »I den yttersta tiden skola bespottare uppstå, som vandra efter sina egna ogudaktiga begärelser.»
Det är dessa människor som vålla söndringar, dessa som äro »själiska» och icke hava ande.
Men I, mina älskade, uppbyggen eder på eder allraheligaste tro, bedjen i den helige Ande,
och bevaren eder så i Guds kärlek, under det att I vänten på vår Herres, Jesu Kristi, barmhärtighet, till evigt liv.
Mot somliga av dem, sådana som äro tvivlande, mån I vara barmhärtiga
och frälsa dem genom att rycka dem ur elden; mot de andra mån I också vara barmhärtiga, dock med fruktan, så att I avskyn till och med deras livklädnad, den av köttet befläckade.
Men honom som förmår bevara eder ifrån fall och ställa eder inför sin härlighet ostraffliga, i fröjd,
honom som allena är Gud, och som är vår Frälsare genom Jesus Kristus, vår Herre, honom tillhör ära, majestät, välde och makt, såsom före all tid, så ock nu och i alla evigheter.
Amen.
Detta är en uppenbarelse från Jesus Kristus, en som Gud gav honom för att visa sina tjänare, vad som snart skall ske.
Och medelst ett budskap genom sin ängel gav han det till känna för sin tjänare Johannes,
som här vittnar och frambär Guds ord och Jesu Kristi vittnesbörd, allt vad han själv har sett.
Salig är den som får uppläsa denna profetias ord, och saliga äro de som få höra dem och som taga vara på, vad däri är skrivet; ty tiden är nära.
Johannes hälsar de sju församlingarna i provinsen Asien.
Nåd vare med eder och frid från honom som är, och som var, och som skall komma, så ock från de sju andar, som stå inför hans tron,
och från Jesus Kristus, det trovärdiga vittnet, den förstfödde bland de döda, den som är härskaren över konungarna på jorden.
Honom som älskar oss, och som har löst oss från våra synder med sitt blod
och gjort oss till ett konungadöme, till präster åt sin Gud och Fader, honom tillhör äran och väldet i evigheternas evigheter, amen.
Se, han kommer med skyarna, och allas ögon skola se honom, ja ock deras som hava stungit honom; och alla släkter på jorden skola jämra sig vid hans åsyn.
Ja, amen.
Jag är A och O, säger Herren Gud, han som är, och som var, och som skall komma, den Allsmäktige.
Jag, Johannes, eder broder, som med eder har del i bedrövelsen och riket och ståndaktigheten i Jesus, jag befann mig på den ö som heter Patmos, för Guds ords och Jesu vittnesbörds skull.
Jag kom i andehänryckning på Herrens dag och fick då bakom mig höra en stark röst, lik ljudet av en basun,
och den sade: »Skriv upp i en bok vad du får se, och sänd den till de sju församlingarna i Efesus och Smyrna och Pergamus och Tyatira och Sardes och Filadelfia och Laodicea.»
Och jag vände mig om för att se vad det var för en röst som talade till mig; och när jag vände mig om, fick jag se sju gyllene ljusstakar
och mitt i bland ljusstakarna någon som liknade en människoson, klädd i en fotsid klädnad och omgjordad kring bröstet med ett gyllene bälte.
Hans huvud och hår var vitt såsom vit ull, såsom snö, och hans ögon voro såsom eldslågor.
Hans fötter liknade glänsande malm, när den har blivit glödgad i en ugn.
Och hans röst var såsom bruset av stora vatten.
I sin högra hand hade han sju stjärnor, och från hans mun utgick ett skarpt tveeggat svärd, och hans ansikte var såsom solen, när den skiner i sin fulla kraft.
När jag såg honom, föll jag ned för hans fötter, såsom hade jag varit död.
Men han lade sin högra hand på mig och sade: »Frukta icke.
Jag är den förste och den siste
och den levande; jag var död, men se, jag lever i evigheternas evigheter och jag har nycklarna till döden och dödsriket.
Så skriv nu upp, vad du har sett, och skriv upp både vad som nu är, och vad som härefter skall ske.
Vad angår hemligheten med de sju stjärnorna, som du har sett i min högra hand, och de sju gyllene ljusstakarna, så må du veta att de sju stjärnorna äro de sju församlingarnas änglar, och att de sju ljusstakarna äro de sju församlingarna.»
Skriv till Efesus' församlings ängel: »Så säger han som håller de sju stjärnorna i sin högra hand, han som går omkring bland de sju gyllene ljusstakarna:
Jag känner dina gärningar och ditt arbete och din ståndaktighet, och jag vet att du icke kan lida onda människor; du har prövat dem som säga sig vara apostlar, men icke äro det, och har funnit dem vara lögnare.
Och du är ståndaktig och har burit mycket för mitt namns skull och har icke förtröttats.
Men jag har det emot dig, att du har övergivit din första kärlek.
Betänk då varifrån du har fallit, och bättra dig, och gör åter sådana gärningar som du gjorde under din första tid.
Varom icke, så skall jag komma över dig och skall flytta din ljusstake från dess plats, såframt du icke gör bättring.
Men den berömmelsen har du, att du hatar nikolaiternas gärningar, som också jag hatar. --
Den som har öra, han höre vad Anden säger till församlingarna.
Den som vinner seger, åt honom skall jag giva att äta av livets träd, som står i Guds paradis.»
Och skriv till Smyrnas församlings ängel: »Så säger den förste och den siste, han som var död och åter har blivit levande:
Jag känner din bedrövelse och din fattigdom -- dock, du är rik! -- och jag vet vilken försmädelse du utstår av dem som säga sig vara judar, men icke äro detta, utan äro en Satans synagoga.
Frukta icke för det som du skall få lida.
Se, djävulen skall kasta somliga av eder i fängelse, för att I skolen sättas på prov; och I skolen få utstå bedrövelse i tio dagar.
Var trogen intill döden, så skall jag giva dig livets krona,
Den som har öra, han höre vad Anden säger till församlingarna.
Den som vinner seger, han skall förvisso icke lida någon skada av den andra döden.»
Och skriv till Pergamus' församlings ängel: »Så säger han som har det skarpa tveeggade svärdet:
Jag vet var du bor: där varest Satan har sin tron.
Och dock håller du fast vid mitt namn; och tron på mig förnekade du icke ens på den tid då Antipas, mitt vittne, min trogne tjänare, blev dräpt hos eder -- där varest Satan bor.
Men jag har något litet emot dig: du har hos dig några som hålla fast vid Balaams lära, hans som lärde Balak huru han skulle lägga en stötesten för Israels barn, så att de skulle äta kött från avgudaoffer och bedriva otukt.
Så har också du några som på lika sätt hålla sig till nikolaiternas lära.
Gör då bättring; varom icke, så skall jag snart komma över dig och skall strida mot dem med min muns svärd.
Den som har öra, han höre vad Anden säger till församlingarna.
Den som vinner seger, åt honom skall jag giva av det fördolda mannat; och jag skall giva honom en vit sten och ett nytt namn skrivet på den stenen, ett namn som ingen känner, utom den som får det.»
Och skriv till Tyatiras församlings ängel: »Så säger Guds Son, han som har ögon såsom eldslågor, han vilkens fötter likna glänsande malm:
Jag känner dina gärningar och din kärlek och din tro, och jag vet huru du har tjänat och varit ståndaktig, och huru dina sista gärningar äro flera än dina första.
Men jag har det emot dig att du är så efterlåten mot kvinnan Jesabel -- hon som säger sig vara en profetissa och uppträder såsom lärare och förleder mina tjänare till att bedriva otukt och till att äta kött från avgudaoffer.
Jag har givit henne tid till bättring, men hon vill icke göra bättring och upphöra med sin otukt.
Se, jag vill lägga henne ned på sjuksängen; och över dem som med henne begå äktenskapsbrott vill jag sända stor vedermöda, såframt de icke bättra sig och upphöra med att göra hennes gärningar.
Och hennes barn skall jag dräpa.
Och alla församlingarna skola förnimma, att jag är den som rannsakar njurar och hjärtan; och jag skall giva var och en av eder efter hans gärningar.
Men till eder, I andra som bon i Tyatira, till eder alla som icke haven denna lära, då I ju icke »haven lärt känna djupheterna», såsom de säga -- ja, Satans djupheter! -- till eder säger jag: Jag lägger icke på eder någon ny börda;
hållen allenast fast vid det som I haven, till dess jag kommer.
Den som vinner seger och intill änden troget gör mina gärningar, åt honom skall jag giva makt över hedningarna.
och han skall styra dem med järnspira, likasom när man krossar lerkärl,
såsom ock jag har fått den makten av min Fader; och jag skall giva honom morgonstjärnan.
Den som har öra, han höre vad Anden säger till församlingarna.»
Och skriv till Sardes' församlings ängel: »Så säger han som har Guds sju andar och de sju stjärnorna: Jag känner dina gärningar; du har det namnet om dig, att du lever, men du är död.
Vakna upp och håll dig vaken, och styrk det som ännu är kvar, det som har varit nära att dö.
Ty jag har icke funnit dina gärningar vara fullkomliga inför min Gud.
Tänk nu på huru du undfick ordet och hörde det, och tag vara på därpå och gör bättring.
Om du icke håller dig vaken, så skall jag komma såsom en tjuv, och du skall förvisso icke veta vilken stund jag kommer över dig.
Dock kunna hos dig i Sardes nämnas några få som icke hava fläckat sina kläder; och dessa skola vandra med mig i vita kläder, ty de äro värdiga därtill.
Den som vinner seger, han skall så bliva klädd i vita kläder, och jag skall aldrig utplåna hans namn ur livets bok, utan kännas vid hans namn inför min Fader och inför hans änglar.
Den som har öra, han höre vad Anden säger till församlingarna.»
Och skriv till Filadelfias församlings ängel: »Så säger den Helige, den Sannfärdige, han som har 'Davids nyckel', han som 'upplåter, och ingen kan tillsluta', han som 'tillsluter, och ingen upplåter':
Jag känner dina gärningar.
Se, jag har låtit dig finna en öppen dörr, som ingen kan tillsluta.
Ty väl är din kraft ringa, men du har tagit vara på mitt ord och icke förnekat mitt namn.
Se, jag vill överlämna åt dig några från Satans synagoga, några av dem som säga sig vara judar, men icke äro det, utan ljuga; ja, jag vill göra så, att de komma ock falla ned för dina fötter, och de skola förstå, att jag har fått dig kär.
Eftersom du har tagit vara på mitt bud om ståndaktighet, skall ock jag taga vara på dig och frälsa dig ut ur den prövningens stund som skall komma över hela världen, för att sätta jordens inbyggare på prov.
Jag kommer snart; håll fast det du har, så att ingen tager din krona.
Den som vinner seger, honom skall jag göra till en pelare i min Guds tempel, och han skall aldrig mer lämna det; och jag skall skriva på honom min Guds namn och namnet på min Guds stad, det nya Jerusalem, som kommer ned från himmelen, från min Gud, så ock mitt eget nya namn.
Den som har öra, han höre vad Anden säger till församlingarna.
Och skriv till Laodiceas församlings ängel: »Så säger han som är Amen, den trovärdiga och sannfärdiga vittnet, begynnelsen till Guds skapelse:
Jag känner dina gärningar: du är varken kall eller varm.
Jag skulle önska att du vore antingen kall eller varm.
Men nu, då du är ljum och varken varm eller kall, skall jag utspy dig ur min mun.
Du säger ju: 'Jag är rik, ja, jag har vunnit rikedomar och behöver intet'; och du vet icke att du just är eländig och ömkansvärd och fattig och blind och naken.
Så råder jag dig då att du köper av mig guld som är luttrat i eld, för att du skall bliva rik, och att du köper vita kläder till att kläda dig i, för att din nakenhets skam icke skall bliva uppenbar, och att du köper ögonsalva till att smörja dina ögon med, för att du skall kunna se.
'Alla som jag älskar, dem tuktar och agar jag.'
Så gör nu bättring med all flit.
Se, jag står för dörren och klappar; om någon lyssnar till min röst och upplåter dörren, så skall jag gå in till honom och hålla måltid med honom och han med mig.
Den som vinner seger, honom skall jag låta sitta med mig på min tron, likasom jag själv har vunnit seger och satt mig med min Fader på hans tron.
Den som har öra, han höre vad Anden säger till församlingarna.
Sedan fick jag se en dörr vara öppnad i himmelen; och den röst, lik ljudet av en basun, som jag förut hade hört tala till mig, sade: »Kom hit upp, så skall jag visa dig, vad som skall ske härefter.»
I detsamma kom jag i andehänryckning.
Och jag fick se en tron vara framsatt i himmelen, och någon satt på den tronen;
och han som satt därpå var till utseendet såsom jaspissten och karneol.
Och runt omkring tronen gick en regnbåge, som till utseendet var såsom en smaragd.
Och jag såg tjugufyra andra troner runt omkring tronen, och på de tronerna sutto tjugufyra äldste, klädda i vita kläder, med gyllene kransar på sina huvuden.
Och från tronen utgingo ljungeldar och dunder och tordön; och framför tronen brunno sju eldbloss, det är Guds sju andar.
Framför tronen syntes ock likasom ett glashav, likt kristall; och runt omkring tronen stodo fyra väsenden, ett mitt för var sida av tronen och de voro fullsatta med ögon framtill och baktill.
Och det första väsendet liknade ett lejon, det andra väsendet liknade en ung tjur, det tredje väsendet hade ett ansikte såsom en människa, det fjärde väsendet liknade en flygande örn.
Och vart och ett av de fyra väsendena hade sex vingar; runt omkring, jämväl under vingarna voro de fullsatta med ögon.
Och dag och natt sade de utan uppehåll: »Helig, helig, helig är Herren Gud den Allsmäktige, han som var, och som är, och som skall komma.»
Och när väsendena hembära pris och ära och tack åt honom som sitter på tronen och tillbedja honom som lever i evigheternas evigheter,
då falla de tjugufyra äldste ned inför honom som sitter på tronen, och tillbedja honom som lever i evigheternas evigheter, och lägga sina kransar ned inför tronen och säga;
»Du, vår Herre och Gud, är värdig att mottaga pris och ära och makt, ty du har skapat allting, och därför att så var din vilja, kom det till och blev skapat.»
Och i högra handen på honom som satt på tronen såg jag en bokrulle, med skrift både på insidan och på utsidan, och förseglad med sju insegel.
Och jag såg en väldig ängel som utropade med hög röst: »Vem är värdig att öppna bokrullen och bryta dess insegel?»
Men ingen, vare sig i himmelen eller på jorden eller under jorden, kunde öppna bokrullen eller se vad som stod däri.
Och jag grät bittert över att ingen befanns vara värdig att öppna bokrullen eller se, vad som stod däri.
Men en av de äldste sade till mig: »Gråt icke.
Se, lejonet av Juda stam, telningen från Davids rot, har vunnit seger, så att han kan öppna bokrullen och och bryta dess sju insegel.»
Då fick jag se att mellan tronen och de fyra väsendena och de äldste stod ett lamm, som såg ut såsom hade det varit slaktat.
Det hade sju horn och sju ögon, det är Guds sju andar, vilka äro utsända över hela jorden.
Och det trädde fram och tog bokrullen ur högra handen på honom som satt på tronen.
Och när han tog bokrullen, föllo de fyra väsendena och de tjugufyra äldste ned inför Lammet; och de hade var och en sin harpa och hade gyllene skålar, fulla med rökelse, det är de heligas böner.
Och de sjöngo en ny sång som lydde så: »Du är värdig att taga bokrullen och att bryta dess insegel, ty du har blivit slaktad, och med ditt blod har du åt Gud köpt människor, av alla stammar och tungomål och folk och folkslag,
och gjort dem åt vår Gud till ett konungadöme och till präster, och de skola regera på jorden»
Och i min syn fick jag höra röster av många änglar runt omkring tronen och omkring väsendena och de äldste; och deras antal var tio tusen gånger tio tusen och tusen gånger tusen.
Och de sade med hög röst: »Lammet som blev slaktat, är värdigt att mottaga makten, så ock rikedom och vishet och starkhet och ära, och pris och lov.»
Och allt skapat, både i himmelen och på jorden och under jorden och på havet, och allt vad i dem var, hörde jag säga: »Honom, som sitter på tronen, och Lammet tillhör lovet och äran och priset och väldet i evigheternas evigheter.»
Och de fyra väsendena sade »amen», och de äldste föllo ned och tillbådo.
Och jag såg Lammet bryta det första av de sju inseglen; och jag hörde ett av de fyra väsendena säga såsom med tordönsröst: »Kom.»
Då fick jag se en vit häst; och mannen som satt på den hade en båge, och en segerkrans blev honom given, och han drog ut såsom segrare och för att segra.
Och när det bröt det andra inseglet, hörde jag det andra väsendet säga »Kom.»
Då kom en annan häst fram, en som var röd; och åt mannen som satt på den blev givet att taga friden bort från jorden, så att människorna skulle slakta varandra.
Och ett stort svärd blev honom givet.
Och när det bröt det tredje inseglet, hörde jag det tredje väsendet säga »Kom.»
Då fick jag se en svart häst; och mannen som satt på den hade en vågskål i sin hand.
Och jag hörde likasom en röst mitt ibland de fyra väsendena säga: »Ett mått vete för en silverpenning och tre mått korn för en silverpenning!
Och oljan och vinet må du icke skada.»
Och när det bröt det fjärde inseglet, hörde jag det fjärde väsendets röst säga: »Kom.»
Då fick jag se en blekgul häst; och mannen som satt på den, hans namn var Döden, och Dödsriket följde med honom.
Och åt dem gavs makt över fjärdedelen av jorden, så att de skulle få dräpa med svärd och genom hungersnöd och pest och genom vilddjuren på jorden.
Och när det bröt det femte inseglet, såg jag under altaret de människors själar, som hade blivit slaktade för Guds ords skull och för det vittnesbörds skull, som de hade.
Och de ropade med hög röst och sade: »Huru länge, du helige och sannfärdige Herre, skall du dröja att hålla dom och att utkräva vårt blod av jordens inbyggare?»
Och åt var och en av dem gavs en vit, fotsid klädnad, och åt dem blev tillsagt att de ännu en liten tid skulle giva sig till ro, till dess jämväl skaran av deras medtjänare och bröder, som skulle bliva dräpta likasom de själva, hade blivit fulltalig.
Och jag såg Lammet bryta det sjätte inseglet.
Då blev det en stor jordbävning, och solen blev svart som en sorgdräkt, och månen blev hel och hållen såsom blod;
och himmelens stjärnor föllo ned på jorden, såsom när ett fikonträd fäller sina omogna frukter, då det skakas av en stark vind.
Och himmelen vek undan, såsom när en bokrulle rullas tillhopa; och alla berg och öar flyttades bort ifrån sin plats.
Och konungarna på jorden och stormännen och krigsöverstarna och alla de rika och de väldiga, ja, alla, både trälar och fria, dolde sig i hålor och bland bergsklippor.
Och de sade till bergen och klipporna: »Fallen över oss och döljen oss för dens ansikte, som sitter på tronen, och för Lammets vrede.
Ty deras vredes stora dag är kommen, och vem kan bestå?»
Sedan såg jag fyra änglar stå vid jordens fyra hörn och hålla tillbaka jordens fyra vindar, för att ingen vind skulle blåsa över jorden eller över havet eller mot något träd.
Och jag såg en annan ängel träda fram ifrån öster med den levande Gudens signet.
Och han ropade med hög röst till de fyra änglar som hade fått sig givet att skada jorden och havet,
och sade: »Gören icke jorden eller havet eller träden någon skada, förrän vi hava tecknat vår Guds tjänare med insegel på deras pannor.»
Och jag fick höra antalet av dem som voro tecknade med insegel, ett hundra fyrtiofyra tusen tecknade, av alla Israels barns stammar;
av Juda stam tolv tusen tecknade, av Rubens stam tolv tusen, av Gads stam tolv tusen,
av Asers stam tolv tusen, av Neftalims stam tolv tusen, av Manasses' stam tolv tusen,
av Simeons stam tolv tusen, av Levi stam tolv tusen, av Isaskars stam tolv tusen,
av Sabulons stam tolv tusen, av Josefs stam tolv tusen, av Benjamins stam tolv tusen tecknade.
Sedan fick jag se en stor skara, som ingen kunde räkna, en skara ur alla folkslag och stammar och folk och tungomål stå inför tronen och inför Lammet; och de voro klädda i vita, fotsida kläder och hade palmer i sina händer.
Och de ropade med hög röst och sade: »Frälsningen tillhör vår Gud, honom som sitter på tronen, och Lammet.»
Och alla änglar, som stodo runt omkring tronen och omkring de äldste och de fyra väsendena, föllo ned på sina ansikten inför tronen och tillbådo Gud
och sade: »Amen.
Lovet och priset och visheten och tacksägelsen och äran och makten och starkheten tillhöra vår Gud i evigheternas evigheter.
Amen.»
Och en av de äldste tog till orda och sade till mig: »Dessa som äro klädda i de vita, fotsida kläderna, vilka äro de, och varifrån hava de kommit?»
Jag svarade honom: »Min herre, du vet själv det.»
Då sade han till mig: »Dessa äro de som komma ur den stora bedrövelsen, och som hava tvagit sina kläder och gjort dem vita i Lammets blod.
Därför stå de inför Guds tron och tjäna honom, dag och natt, i hans tempel.
Och han som sitter på tronen skall slå upp sitt tabernakel över dem.
'De skola icke mer hungra och icke mer törsta, och solens hetta skall icke träffa dem, ej heller eljest någon brännande hetta.
Ty Lammet, som står mitt för tronen, skall vara deras herde och leda dem till livets vattenkällor, och 'Gud skall avtorka alla tårar från deras ögon'.»
Och när Lammet bröt det sjunde inseglet, uppstod i himmelen en tystnad, som varade vid pass en halv timme.
Och jag fick se de sju änglar, som stå inför Gud; åt dem gåvos sju basuner.
Och en annan ängel kom och ställde sig vid altaret, och han hade ett gyllene rökelsekar; och mycken rökelse var given åt honom, för att han skulle lägga den till alla de heligas böner på det gyllene altare som stod framför tronen.
Och ur ängelns hand steg röken av rökelsen med de heligas böner upp inför Gud.
Och ängeln tog rökelsekaret och fyllde det med eld från altaret och kastade elden ned på jorden.
Då kommo tordön och dunder och ljungeldar och jordbävning.
Och de sju änglarna, som hade de sju basunerna, gjorde sig redo att stöta i sina basuner.
Och den förste stötte i sin basun.
Då kom hagel och eld, blandat med blod, och det kastades ned på jorden; och tredjedelen av jorden brändes upp, och tredjedelen av träden brändes upp, och allt grönt gräs brändes upp.
Och den andre ängeln stötte i sin basun.
Då var det som om ett stort brinnande berg hade blivit kastat i havet; och tredjedelen av havet blev blod.
Och tredjedelen av de levande varelser som funnos i havet omkom; och tredjedelen av skeppen förgicks.
Och den tredje ängeln stötte i sin basun.
Då föll från himmelen en stor stjärna, brinnande såsom ett bloss; och den föll ned över tredjedelen av strömmarna och över vattenkällorna.
Och stjärnans namn var Malört.
Och tredjedelen av vattnet blev bitter malört; och många människor omkommo genom vattnet, därför att det hade blivit så bittert.
Och den fjärde ängeln stötte i sin basun.
Då drabbade hemsökelsen tredjedelen av solen och tredjedelen av månen och tredjedelen av stjärnorna, så att tredjedelen av dem förmörkades och dagen miste tredjedelen av sitt ljus, sammalunda ock natten.
Sedan fick jag i min syn höra en örn, som flög fram uppe i himlarymden, ropa med hög röst: »Ve, ve, ve över jordens inbyggare, när de tre övriga änglar, som skola stöta i basun, låta sina basuner ljuda!»
Och den femte ängeln stötte i sin basun.
Då såg jag en stjärna vara fallen ifrån himmelen ned på jorden; och åt henne gavs nyckeln till avgrundens brunn.
Och hon öppnade avgrundens brunn.
Då steg en rök upp ur brunnen, lik röken från en stor ugn, och solen och luften förmörkades av röken från brunnen.
Och ur röken kommo gräshoppor ut över jorden; och åt dem gavs samma makt som skorpionerna på jorden hava.
Och dem blev tillsagt, att de icke skulle skada gräset på jorden eller något annat grönt eller något träd, utan allenast de människor som icke hade Guds insegel på sina pannor.
Och åt dem blev givet att, icke att döda dem, men att plåga dem i fem månader; och plågan, som de vållade var såsom den plåga en skorpion åstadkommer, när den stinger en människa.
På den tiden skola människorna söka döden, men icke kunna finna den; de skola åstunda att dö, men döden skall fly undan ifrån dem.
Och gräshopporna tedde sig såsom hästar, rustade till strid.
På sina huvuden hade de likasom kransar, som syntes vara av guld.
Deras ansikten voro såsom människors ansikten.
De hade hår såsom kvinnors hår, och deras tänder voro såsom lejons.
De hade bröst, som liknade järnpansar; och rasslet av deras vingar var såsom vagnsrasslet, när många hästar med sina vagnar störta fram till strid.
De hade stjärtar med gaddar, såsom skorpioner hava; och i deras stjärtar låg den makt de hade fått att i fem månader skada människorna.
Till konung över sig hade de avgrundens ängel, vilkens namn på hebreiska är Abaddon och som på grekiska har namnet Apollyon.
Det första ve har gått till ända; se, efter detta komma ännu två andra ve.
Och den sjätte ängeln stötte i sin basun.
Då hörde jag en röst från de fyra hornen på det gyllene altare, som stod inför Guds ansikte,
säga till den sjätte ängeln, den som hade basunen: »Lös de fyra änglar, som hållas bundna invid den stora floden Eufrat.»
Och de fyra änglarna löstes, de som just för den timmen, på den dagen, i den månaden, under det året hade hållits redo att dräpa tredjedelen av människorna.
Och antalet ryttare i de ridande skarorna var två gånger tio tusen gånger tio tusen; jag fick höra att de voro så många.
Och hästarna och männen som sutto på dem tedde sig för min syn på detta sätt: männen hade eldröda och mörkblå och svavelgula pansar; och hästarna hade huvuden såsom lejon, och ur deras gap gick ut eld och rök och svavel.
Av dessa tre plågor -- av elden och röken och svavlet som gick ut ur deras gap -- dödades tredjedelen av människorna.
Ty hästarnas makt låg i deras gap och i deras svansar.
Deras svansar liknade nämligen ormar, och hade huvuden, och med dem var det, som de gjorde skada.
Men de återstående människorna, de som icke hade blivit dödade genom dessa plågor, gjorde icke bättring; de vände sig icke ifrån belätena, som de hade gjort med egna händer, och upphörde icke att tillbedja onda andar och avgudar av guld och silver och koppar och sten och trä, som varken kunna se eller höra eller gå.
De gjorde icke bättring och upphörde icke med sina mordgärningar och trolldomskonster, sin otukt och sitt tjuveri.
Och jag såg en annan väldig ängel komma ned från himmelen.
Han var klädd i en sky och hade regnbågen över sitt huvud, och hans ansikte var såsom solen, och hans ben voro såsom eldpelare;
och i sin hand hade han en öppen liten bokrulle.
Och han satte sin högra fot på havet och sin vänstra på jorden.
Och han ropade med hög röst, såsom när ett lejon ryter.
Och när han hade ropat, läto de sju tordönen höra sina röster.
Och sedan de sju tordönen hade talat, tänkte jag skriva, men jag fick då höra en röst från himmelen säga: »Göm såsom under insegel vad de sju tordönen hava talat, och skriv icke upp det.»
Och ängeln, som jag såg stå på havet och på jorden, lyfte sin högra hand upp mot himmelen
och svor vid honom som lever i evigheternas evigheter, vid honom som har skapat himmelen och vad däri är, och jorden och vad därpå är, och havet och vad däri är, och sade: »Ingen tid skall mer givas,
utan i de dagar, då den sjunde ängelns röst höres, när det sker att han stöter i sin basun, då är Guds hemliga rådslut fullbordat, i enlighet med det glada budskap som han har förkunnat för sina tjänare profeterna.»
Och den röst som jag hade hört från himmelen hörde jag nu åter tala till mig; den sade: »Gå och tag den öppna bokrulle som ängeln har i sin hand, han som står på havet och på jorden.»
Då gick jag bort till ängeln och bad honom att han skulle giva mig bokrullen.
Och han sade till mig: »Tag den och ät upp den; den skall vålla dig bitter plåga i din buk, men i din mun skall den vara söt såsom honung.»
Då tog jag bokrullen ur ängelns hand och åt upp den; och den var i min mun söt såsom honung, men när jag hade ätit upp den, kände jag bitter plåga i min buk.
Och mig blev sagt: »Du måste än ytterligare profetera om många folk och folkslag och tungomål och konungar.
Och ett rör, likt en mätstång, gavs åt mig, och mig blev sagt: »Stå upp och mät Guds tempel och altaret tillika med dem som tillbedja därinne.
Men lämna å sido templets yttre förgård och mät den icke; ty den är prisgiven åt hedningarna, och de skola under fyrtiotvå månader förtrampa den heliga staden.
Och jag skall låta mina två vittnen under ett tusen två hundra sextio dagar profetera, höljda i säcktyg.
Dessa vittnen äro de två olivträd och de två ljusstakar som stå inför jordens Herre.
Och om någon vill göra dem skada, så går eld ut ur deras mun och förtär deras ovänner; ja, om någon vill göra dem skada, så skall han bliva dödad på det sättet.
De hava makt att tillsluta himmelen, så att intet regn faller under den tid de profetera; de hava ock makt över vattnet, att förvandla det till blod, och makt att slå jorden med alla slags plågor, så ofta de vilja.
Och när de hava till fullo framburit sitt vittnesbörd, skall vilddjuret, det som skall stiga upp ur avgrunden, giva sig i strid med dem och skall övervinna dem och döda dem.
Och deras döda kroppar skola bliva liggande på gatan i den stora staden som, andligen talat, heter Sodom och Egypten, den stad där också deras Herre blev korsfäst.
Och människor av allahanda folk och stammar och tungomål och folkslag skola i tre och en halv dagar se deras döda kroppar ligga där, och de skola icke tillstädja att kropparna läggas i någon grav.
Och jordens inbyggare skola glädjas över vad som har vederfarits dem och skola fröjda sig och sända varandra gåvor; ty dessa två profeter hade varit en plåga för jordens inbyggare.»
Men efter tre och en halv dagar kom livets ande från Gud in i dem, och de reste sig upp på sina fötter; och en stor fruktan föll över dem som sågo dem.
Och de hörde en stark röst från himmelen, som sade till dem: »Kommen hit upp.»
Då stego de i en sky upp till himmelen, i sina ovänners åsyn.
Och i samma stund blev det en stor jordbävning, och tiondedelen av staden störtade samman, och genom jordbävningen omkommo sju tusen människor; och de övriga blevo förskräckta och gåvo ära åt Gud i himmelen.
Det andra ve har gått till ända; se, det tredje ve kommer snart.
Och den sjunde ängeln stötte i sin basun.
Då ljödo i himmelen starka röster som sade: »Väldet över världen har blivit vår Herres och hans Smordes, och han skall vara konung i evigheternas evigheter.»
Och de tjugufyra äldste, som sutto på sina troner inför Gud, föllo ned på sina ansikten och tillbådo Gud
och sade: »Vi tacka dig, Herre Gud, du Allsmäktige, du som är, och som var, för att du har tagit i besittning din stora makt och trätt fram såsom konung.
Folken vredgades, men din vredes dag har nu kommit, och den tid då de döda skola få sin dom, och då du skall löna dina tjänare profeterna och de heliga och dem som frukta ditt namn, både små och stora, och då du skall fördärva dem som fördärva jorden.»
Och Guds tempel i himmelen öppnades, och hans förbundsark blev synlig i hans tempel.
Då kommo ljungeldar och dunder och tordön och jordbävning och starkt hagel.
Och ett stort tecken visade sig i himmelen: där syntes en kvinna, som hade solen till sin klädnad och månen under sina fötter, och en krans av tolv stjärnor på sitt huvud.
Hon var havande och ropade i barnsnöd och födslovånda.
Ännu ett annat tecken visade sig i himmelen: där syntes en stor röd drake, som hade sju huvuden och tio horn, och på sina huvuden sju kronor.
Och hans stjärt drog med sig tredjedelen av himmelens stjärnor och kastade den ned på jorden.
Och draken stod framför kvinnan som skulle föda, ty han ville uppsluka hennes barn, när hon hade fött det.
Och hon födde ett barn gossebarn, som en gång skall styra alla folk med järnspira.
Men hennes barn blev uppryckt till Gud och till hans tron;
Och kvinnan flydde ut i öknen, där hon har en plats sig beredd av Gud, och där hon skulle få sitt uppehälle under ett tusen två hundra sextio dagar.
Och en strid uppstod i himmelen: Mikael och hans änglar gåvo sig i strid med draken; och draken och hans änglar stridde mot dem,
men de förmådde intet mot dem, och i himmelen fanns nu icke mer någon plats för dem.
Och den store draken, den gamle ormen, blev nedkastad, han som kallas Djävul och Satan, och som förvillar hela världen; han blev nedkastad till jorden, och hans änglar kastades ned jämte honom.
Och jag hörde en stark röst i himmelen säga: »Nu har frälsningen och makten och riket blivit vår Guds, och väldet hans Smordes; ty våra bröders åklagare är nedkastad, han som dag och natt anklagade dem inför vår Gud.
De övervunno honom i kraft av Lammets blod och i kraft av sitt vittnesbörds ord: de älskade icke så sitt liv, att de drogo sig undan döden.
Glädjens fördenskull, I himlar och I som bon i dem.
Men ve dig, du jord, och dig, du hav!
Ty djävulen har kommit ned till eder i stor vrede, eftersom han vet att den tid han har kvar är kort.»
Och när draken såg att han var nedkastad på jorden, förföljde han kvinnan, som hade fött gossebarnet.
Men åt kvinnan gåvos den stora örnens två vingar, för att hon skulle flyga ut i öknen till den plats där hon skulle få sitt uppehälle under en tid och tider och en halv tid, fjärran ifrån ormens åsyn.
Då sprutade ormen ur sitt gap vatten efter kvinnan såsom en ström, för att strömmen skulle bortföra henne.
Men jorden kom kvinnan till hjälp; jorden öppnade sin mun och drack upp strömmen, som draken hade sprutat ut ur sitt gap.
Och draken vredgades än mer på kvinnan och gick åstad för att föra krig mot de övriga av hennes säd, mot dem som hålla Guds bud och hava Jesu vittnesbörd.
Och han ställde sig på sanden invid havet.
Då såg jag ett vilddjur stiga upp ur havet; det hade tio horn och sju huvuden, och på sina horn hade det tio kronor och på sina huvuden hädiska namn.
Och vilddjuret, som jag såg, liknade en panter, men det hade fötter såsom en björn och gap såsom ett lejon.
Och draken gav det sin makt och sin tron och gav det stor myndighet.
Och jag såg ett av dess huvuden vara likasom sårat till döds, men dess dödssår blev läkt.
Och hela jorden såg med förundran efter vilddjuret.
Och de tillbådo draken, därför att han hade givit vilddjuret sådan myndighet; de tillbådo och vilddjuret och sade »Vem är lik vilddjuret, och vem kan strida mot det?»
Och det fick en mun sig given, som talade stora ord och vad hädiskt var, och det fick makt att så göra under fyrtiotvå månader.
Och den öppnade sin mun till att föra hädiskt tal mot Gud, till att häda hans namn och hans tabernakel och dem som bo i himmelen.
Och det fick makt att föra krig mot de heliga och att övervinna dem; och det fick makt över alla stammar och folk och tungomål och folkslag.
Och alla jordens inbyggare skola tillbedja det, ja, envar som icke har sitt namn från världens begynnelse skrivet i livets bok, det slaktade Lammets bok.
Den som har öra, han höre.
Den som för andra bort i fångenskap, han skall själv bliva bortförd i fångenskap; den som dräper andra med svärd, han skall själv bliva dräpt med svärd.
Här gäller det för de heliga att hava ståndaktighet och tro.
Och jag såg ett annat vilddjur stiga upp ur jorden; det hade två horn, lika ett lamms, och det talade såsom en drake.
Och det utövar det första vilddjurets hela myndighet, i dess åsyn.
Och det kommer jorden och dem som bo därpå att tillbedja det första vilddjuret, det vars dödssår blev läkt.
Och det gör stora tecken, så att det till och med låter eld i människornas åsyn falla ned från himmelen på jorden.
Och genom de tecken, som det har fått makt att göra i vilddjurets åsyn, förvillar det jordens inbyggare; det förmår genom sitt tal jordens inbyggare att göra en bild åt vilddjuret, det som var sårat med svärd, men åter kom till liv.
Och det fick makt att giva ande åt vilddjurets bild, så att vilddjurets bild till och med kunde tala och kunde låta döda alla som icke tillbådo vilddjurets bild.
Och det förmår alla, både små och stora, både rika och fattiga, både fria och trälar, att låta giva sig ett märke på högra handen eller på pannan,
så att ingen får vare sig köpa eller sälja något, utom den som är märkt med vilddjurets namn eller dess namns tal.
Här gäller det att vara vis; den som har förstånd, han räkne ut betydelsen av vilddjurets tal, ty det är en människas tal.
Och dess tal är sex hundra sextiosex.
Och jag fick se Lammet stå på Sions berg jämte det ett hundra fyrtiofyra tusen som hade dess namn och dess Faders namn skrivna på sina pannor.
Och jag hörde ett ljud från himmelen, likt bruset av stora vatten och dånet av ett starkt tordön; och ljudet som jag hörde var såsom när harpospelare spela på sina harpor.
Och de sjöngo inför tronen och inför de fyra väsendena och de äldste vad som tycktes vara en ny sång; och ingen kunde lära sig den sången, utom de ett hundra fyrtiofyra tusen som voro friköpta ifrån jorden.
Dessa äro de som icke hava orenat sig med kvinnor; ty de äro såsom jungfrur.
Dessa äro de som följa Lammet varthelst det går.
De hava blivit friköpta ifrån människorna till en förstling åt Gud och Lammet.
Och i deras mun har ingen lögn blivit funnen; de äro ostraffliga.
Och jag såg en annan ängel flyga fram uppe i himlarymden; han hade ett evigt evangelium, som han skulle förkunna för dem som bo på jorden, för alla folkslag och stammar och tungomål och folk.
Och han sade med hög röst: »Frukten Gud och given honom ära; ty stunden är kommen, då han skall hålla dom.
Ja, tillbedjen honom som har skapat himmel och jord och hav och vattenkällor.
Och ännu en annan ängel följde honom; denne sade: »Fallet, fallet är det stora Babylon, som har givit alla folk att dricka av sin otukts vredesvin.»
Och ännu en tredje ängel följde dem; denne sade med hög röst: »Om någon tillbeder vilddjuret och dess bild och tager dess märke på sin panna eller på sin hand,
så skall ock han få dricka av Guds vredesvin, det som är iskänkt i hans vredes kalk, obemängt; och han skall bliva plågad med eld och svavel, i heliga änglars och i Lammets åsyn.
Och när de så plågas, uppstiger röken därav i evigheters evigheter, och de hava ingen ro, vaken dag eller natt, de som tillbedja vilddjuret och dess bild, eller som låta märka sig med dess namn.
Här gäller det för de heliga att hava ståndaktighet, för dem som hålla Guds bud och bevara tron på Jesus.»
Och jag hörde en röst från himmelen säga: »Skriv: Saliga äro de döda som dö i Herren härefter.
Ja, säger Anden, de skola få vila sig från sitt arbete, ty deras gärningar följa dem.»
Och jag fick se en vit sky, och på skyn satt en som liknade en människoson; och han hade på sitt huvud en gyllene krans, och i sin hand en vass lie.
Och en annan ängel kom ut ur templet och ropade med hög röst till den som satt på skyn: »Låt din lie gå, och inbärga skörden; ty skördetiden är kommen, och säden på jorden är fullt mogen till skörd.»
Den som satt på skyn högg då till med sin lie på jorden, och jorden blev avbärgad.
Och en annan ängel kom ut ur templet i himmelen, och jämväl han hade en vass lie.
Och ännu en ängel kom fram ifrån altaret, den som hade makt över elden.
Denne ropade med hög röst till den som hade den vassa lien; han sade »Låt din vassa lie gå, och skär av druvklasarna från vinträden på jorden, ty deras druvor äro fullmogna.»
Och ängeln högg till med sin lie på jorden och skar av frukten ifrån vinträden på jorden och kastade den i Guds vredes stora vinpress.
Och vinpressen trampade utanför staden, och blod gick ut från pressen och steg ända upp till betslen på hästarna, på en sträcka av ett tusen sex hundra stadier.
Och jag såg ett annat tecken i himmelen, stort och underbart; sju änglar med de sju plågor som bliva de sista, ty med dem är Guds vredesdom fullbordad.
Och jag fick se något som såg ut såsom ett glashav, blandat med eld.
Och jag såg dem som hade vunnit seger över vilddjuret, med dess bild och dess namns tal, stå vid glashavet, med Guds harpor i sina händer.
Och de sjöngo Moses', Guds tjänares, sång och Lammets sång: de sjöngo: »Stora och underbara äro dina verk, Herre Gud, du Allsmäktige; rättfärdiga och rätta äro dina vägar, du folkens konung.
Vem skulle icke frukta dig, Herre, och prisa ditt namn?
Du allena är helig, och alla folk skola komma och tillbedja inför dig.
Ty dina domar hava blivit uppenbara.»
Sedan såg jag att vittnesbördets tabernakels tempel i himmelen öppnades.
Och de sju änglarna med de sju plågorna kommo ut ur templet, klädda i rent, skinande linne, och omgjordade kring bröstet med gyllene bälten.
Och ett av de fyra väsendena gav de sju änglarna sju gyllene skålar, fulla av Guds vrede, hans som lever i evigheternas evigheter.
Och templet blev uppfyllt av rök från Guds härlighet och från hans makt, och ingen kunde gå in i templet, förrän de sju änglarnas sju plågor hade fått sin fullbordan.
Och jag hörde en stark röst från templet säga till de sju änglarna: »Gån åstad och gjuten ut Guds sju vredesskålar på jorden.»
Och den förste gick åstad och göt ut sin skål på jorden.
Då kommo onda och svåra sårnader på de människor som buro vilddjurets märke och tillbådo dess bild.
Och den andre göt ut sin skål i havet.
Då förvandlades det till blod, likt blodet av en död människa, och alla levande varelser i havet dogo.
Och den tredje göt ut sin skål i strömmarna och vattenkällorna.
Då förvandlades dessa till blod.
Och jag hörde vattnens ängel säga: »Rättfärdig är du, du som är och som var, du helige, som har dömt så.
De hava utgjutit heliga mäns och profeters blod.
Därför har ock du givit dem blod att dricka; de äro det värda.»
Och jag hörde altaret säga: »Ja, Herre Gud, du Allsmäktige, rätta och rättfärdiga äro dina domar.»
Och den fjärde göt ut sin skål över solen.
Då fick denna makt att bränna människorna såsom med eld.
Och när nu människorna blevo brända av stark hetta, hädade de Guds namn, hans som hade makten över dessa plågor; de gjorde icke bättring och gåvo honom icke ära.
Och den femte göt ut sin skål över vilddjurets tron.
Då blev dess rike förmörkat, och människorna beto sönder sina tungor i sin vånda.
Och de hädade himmelens Gud för sin våndas och sina sårnaders skull; de gjorde icke bättring och upphörde icke med sina gärningar.
Och den sjätte göt ut sin skål över den stora floden Eufrat.
Då torkade dess vatten ut, för att väg skulle beredas åt konungarna från östern.
Och ur drakens gap och ur vilddjurets gap och ur den falske profetens mun såg jag tre orena andar utgå, lika paddor.
De äro nämligen onda andar som göra tecken, och som gå ut till konungarna i hela världen, för att samla dem till striden på Guds, den Allsmäktiges, stora dag.
(»Se, jag kommer såsom en tjuv; salig är den som vakar och bevarar sina kläder, så att han icke måste gå naken, och man får se hans skam.»)
Och de församlade dem till den plats som på hebreiska heter Harmagedon.
Och den sjunde göt ut sin skål i luften.
Då gick en stark röst ut från tronen i templet och sade »Det är gjort.»
Och nu kommo ljungeldar och dunder och tordön, och det blev en stor jordbävning, en jordbävning så våldsam och så stor, att dess like icke hade förekommit, alltsedan människor blevo till på jorden.
Och den stora staden rämnade söder i tre delar, och folkens städer störtade samman; och Gud kom ihåg det stora Babylon, så att han räckte det kalken med sin stränga vredes vin.
Och alla öar flydde, och inga berg funnos mer.
Och stora hagel, centnertunga, föllo ned från himmelen på människorna; och människorna hädade Gud för den plåga som haglen vållade, ty den plågan var mycket stor.
Och en av de sju änglarna med de sju skålarna kom och talade med mig och sade: »Kom hit, så skall jag visa dig, huru den stora skökan får sin dom, hon som tronar vid stora vatten,
hon som jordens konungar hava bedrivit otukt med och av vilkens otukts vin jordens inbyggare hava druckit sig druckna.»
Sedan förde han mig i anden bort till en öken.
Där såg jag en kvinna som satt på ett scharlakansrött vilddjur, fulltecknat med hädiska namn; och det hade sju huvuden och tio horn.
Och kvinnan var klädd i purpur och scharlakan och glänste av guld och ädla stenar och pärlor; och i sin hand hade hon en gyllene kalk, full av styggelser och av hennes otukts orenlighet.
Och på hennes panna var skrivet ett namn med hemlig betydelse: »Det stora Babylon, hon som är moder till skökorna och till styggelserna på jorden.»
Och jag såg kvinnan vara drucken av de heligas blod och av Jesu vittnens blod.
Och jag förundrade mig storligen, när jag såg henne.
Och ängeln sade till mig: »Varför förundrar du dig?
Jag skall säga dig hemligheten om kvinnan, och om vilddjuret som bär henne, och som har de sju huvudena och de tio hornen.
Vilddjuret som du har sett, det har varit, och är icke mer; men det skall stiga upp ur avgrunden, och det går sedan i fördärvet.
Och de av jordens inbyggare, vilkas namn icke från världens begynnelse äro skrivna i livets bok, skola förundra sig, när de få se vilddjuret som har varit, och icke mer är, men dock skall komma. --
Här gäller det att äga ett förstånd med vishet.
De sju huvudena äro sju berg, som kvinnan tronar på.
De äro ock sju konungar;
fem av dem hava fallit, en är, och den återstående har ännu icke kommit, och när han kommer, skall han bliva kvar en liten tid.
Och vilddjuret som har varit, och icke mer är, det är självt den åttonde, och dock en av de sju, och det går i fördärvet.
Och de tio horn som du har sett, de äro tio konungar, som ännu icke hava kommit till konungavälde, men som för en kort tid, tillika med vilddjuret, få makt såsom konungar.
Dessa hava ett och samma sinne, och de giva sin makt och myndighet åt vilddjuret.
De skola giva sig i strid med Lammet; men Lammet jämte de kallade och utvalda och trogna som följa det, skall övervinna dem, ty Lammet är herrarnas herre och konungarnas konung.»
Och han sade ytterligare till mig: »Vattnen som du har sett, där varest skökan tronar, äro folk och människoskaror och folkslag och tungomål.
Och de tio horn, som du har sett, och vilddjuret, de skola hata skökan och göra henne utblottad och naken, och skola äta hennes kött och bränna upp henne i eld.
Ty Gud har ingivit dem i hjärtat att de skola utföra vad han har i sinnet, och att de alla skola handla i ett och samma sinne, och att de skola giva sitt välde åt vilddjuret, till dess Guds utsagor hava fullbordats.
Och kvinnan som du har sett är den stora staden, som har konungsligt välde över jordens konungar.»
Därefter såg jag en annan ängel komma ned från himmelen; han hade stor makt, och jorden upplystes av hans härlighet.
Och han ropade med stark röst och sade: »Fallet, fallet är det stora Babylon; det har blivit en boning för onda andar, ett tillhåll för alla slags orena andar och ett tillhåll för alla slags orena och vederstyggliga fåglar.
Ty av hennes otukts vredesvin hava alla folk druckit; konungarna på jorden hava bedrivit otukt med henne, och köpmännen på jorden hava skaffat sig rikedom genom hennes omåttliga vällust.»
Och jag hörde en annan röst från himmelen säga: »Dragen ut ifrån henne, I mitt folk, så att I icke gören eder delaktiga i hennes synder och fån eder del av hennes plågor.
Ty hennes synder räcka ända upp till himmelen, och Gud har kommit ihåg hennes orättfärdiga gärningar.
Vedergällen henne vad hon har gjort, ja, given henne dubbelt igen för hennes gärningar; iskänken dubbelt åt henne i den kalk vari hon har iskänkt.
Så mycken ära och vällust som hon har berett sig, så mycken pina och sorg mån I bereda henne.
Eftersom hon säger i sitt hjärta: 'Jag tronar såsom drottning och och sitter icke såsom änka, och aldrig skall jag veta av någon sorg',
därför skola på en och samma dag hennes plågor komma över henne: död och sorg och hungersnöd; och hon skall brännas upp i eld.
Ty stark är Herren Gud, han som har dömt henne.
Och jordens konungar, som hava bedrivit otukt och levat i vällust med henne, skola gråta och jämra sig över henne, när de se röken av hennes brand.
De skola stå långt ifrån, av förfäran över hennes pina, och skola säga: 'Ve, ve dig, Babylon, du stora stad, du starka stad!
Plötsligt har nu din dom kommit.'
Och köpmännen på jorden gråta och sörja över henne, då nu ingen mer köper de varor som de frakta:
guld och silver, ädla stenar och pärlor, fint linne och purpur, siden och scharlakan, allt slags välluktande trä, alla slags arbeten av elfenben och dyrbaraste trä, av koppar och järn och marmor,
därtill kanel och kostbar salva, rökverk, smörjelse och välluktande harts, vin och olja, fint mjöl och vete, fäkreatur och får, hästar och vagnar, livegna och trälar.
De frukter som din själ hade begär till hava försvunnit ifrån dig; allt vad kräsligt och präktigt du hade har gått förlorat för dig och skall aldrig mer bliva funnet.
De som handlade med sådant, de som skaffade sig rikedom genom henne, de skola stå långt ifrån, av förfäran över hennes pina; de skola gråta och sörja
och skola säga: 'Ve, ve dig, du stora stad, du som var klädd i fint linne och purpur och scharlakan, du som glänste av guld och ädla stenar och pärlor!
I ett ögonblick har nu denna stora rikedom blivit förödd.'
Och alla skeppare och alla kustfarare och sjömän och alla andra som hava sitt arbete på havet stå långt ifrån;
och när de ser röken av hennes brand, ropa de och säga: 'Var fanns den stora stadens like?'
Och de strö stoft på sina huvuden och ropa under gråt och sorg och säga: 'Ve, ve dig, du stora stad, genom vars skatter alla de därinne, som hade skepp på havet, blevo rika!
I ett ögonblick har den nu blivit förödd.
Gläd dig över vad som har vederfarits henne, du himmel och I helige och I apostlar och profeter, då nu Gud har hållit dom över henne och utkrävt vedergällning för eder!»
Och en väldig ängel tog upp en sten, lik en stor kvarnsten, och kastade den i havet och sade: »Så skall Babylon, den stora staden, med fart störtas ned och aldrig mer bliva funnen.
Av harpospelare och sångare, av flöjtblåsare och basunblåsare skall aldrig mer något ljud bliva hört i dig; aldrig mer skall någon konstförfaren man av något slags yrke finnas i dig; bullret av en kvarn skall aldrig mer höras i dig;
en lampas sken skall aldrig mer lysa i dig; rop för brudgum och brud skall aldrig mer höras i dig -- du vars köpmän voro stormän på jorden, du genom vars trolldom alla folk blevo förvillade,
och i vilken man såg profeters och heliga mäns blod, ja, alla de människors blod, som hade blivit slaktade på jorden.»
Sedan hörde jag likasom starka röster av en stor skara i himmelen, som sade »Halleluja!
Frälsningen och äran och makten tillhöra vår Gud.
Ty rätta och rättfärdiga äro hans domar; han har dömt den stora skökan, som fördärvade jorden genom sin otukt, och han har utkrävt sina tjänares blod av hennes hand.»
Och åter sade de: »Halleluja!»
Och röken från henne stiger upp i evigheternas evigheter!
Och de tjugufyra äldste och de fyra väsendena föllo ned och tillbådo Gud, som satt på tronen; de sade: »Amen!
Halleluja!»
Och från tronen utgick en röst, som sade: »Loven vår Gud, alla I hans tjänare, I som frukten honom, både små och stora.»
Och jag hörde likasom röster av en stor skara, lika bruset av stora vatten och dånet av starka tordön; de sade: »Halleluja!
Herren, vår Gud, den Allsmäktige, har nu trätt fram såsom konung.
Låtom oss glädjas och fröjda oss och giva honom äran; ty tiden är inne för Lammets bröllop, och dess brud har gjort sig redo.
Och åt henne har blivit givet att kläda sig i fint linne, skinande och rent.»
Det fina linnet är de heligas rättfärdighet.
Och han sade till mig: »Skriv: Saliga äro de som äro bjudna till Lammets bröllopsmåltid.»
Ytterligare sade han till mig: »Dessa ord äro sanna Guds ord.»
Och jag föll ned för hans fötter för att tillbedja honom, men han sade till mig: »Gör icke så.
Jag är din medtjänare och dina bröders, deras som hava Jesu vittnesbörd.
Gud skall du tillbedja.
Ty Jesu vittnesbörd är profetians ande.»
Och jag såg himmelen öppen och fick där se en vit häst; och mannen som satt på den heter »Trofast och sannfärdig», och han dömer och strider i rättfärdighet.
Hans ögon voro såsom eldslågor, och på sitt huvud bar han många kronor och hade ett namn där skrivet, som ingen känner utom han själv.
Och han var klädd i en mantel som var doppad i blod; och det namn han har fått är »Guds Ord».
Och honom följde, på vita hästar, de himmelska härskarorna, klädda i fint linne, vitt och rent.
Och från hans mun utgick ett skarpt svärd, varmed han skulle slå folken.
Och han skall styra dem med järnspira; och han trampar Guds, den Allsmäktiges, stränga vredes vinpress.
Och på sin mantel, över sin länd, har han detta namn skrivet: »Konungarnas konung och herrarnas herre.»
Och jag såg en ängel stå i solen, och denne ropade med hög röst och sade till alla fåglar som flögo fram uppe i himlarymden: »Kommen hit, församlen eder till Guds stora gästabud,
för att äta kött av konungar och krigsöverstar och hjältar, kött av hästar och deras ryttare, ja, kött av alla, både fria och trälar, både små och stora.»
Och jag såg vilddjuret och konungarna på jorden med sina härskaror, samlade för att utkämpa sin strid mot honom som satt på hästen och mot hans härskara.
Och vilddjuret blev gripet, därjämte ock den falske profeten, som i dess åsyn hade gjort de tecken med vilka han hade förvillat dem som hade tagit vilddjurets märke, och dem som hade tillbett dess bild.
Båda blevo de levande kastade i eldsjön, som brann med svavel.
Och de andra blevo dräpta med ryttarens svärd, det som utgick från hans mun; och alla fåglar blevo mättade av deras kött.
Och jag såg en ängel komma ned från himmelen; han hade nyckeln till avgrunden och hade en stor kedja i sin hand.
Och han grep draken, den gamle ormen, det är djävulen och Satan, och fängslade honom för tusen år
och kastade honom i avgrunden och stängde igen och satte dit ett insegel över honom på det att han icke mer skulle förvilla folken, förrän de tusen åren hade gått till ända.
Därefter skall han åter komma lös för en liten tid.
Och jag såg troner stå där, och de satte sig på dem, de åt vilka gavs makt att hålla dom.
Och jag såg de människors själar, som hade blivit halshuggna för Jesu vittnesbörds och Guds Ords skull, och som icke hade tillbett vilddjuret eller dess bild, och icke heller tagit dess märke på sina pannor och sina händer; dessa blevo nu åter levande och fingo regera med Kristus i tusen år.
(De övriga döda blevo icke levande, förrän de tusen åren hade gått till ända.)
Detta är den första uppståndelsen.
Salig och helig är den som har del i den första uppståndelsen; över dem har den andra döden ingen makt, utan de skola vara Guds och Kristi präster och skola få regera med honom de tusen åren.
Men när de tusen åren hava gått till ända, skall Satan komma lös ur sitt fängelse.
Han skall då gå ut för att förvilla de folk som bo vid jordens fyra hörn, Gog och Magog, och samla dem till den stundande striden; och de äro till antalet såsom sanden i havet.
Och de draga fram över jordens hela vidd och omringa de heligas läger och »den älskade staden»; men eld faller ned från himmelen och förtär dem.
Och djävulen, som förvillade dem, bliver kastad i samma sjö av eld och svavel, dit vilddjuret och den falske profeten hade blivit kastade; och de skola där plågas dag och natt i evigheternas evigheter.
Och jag såg en stor vit tron och honom som satt därpå; och för hans ansikte flydde jord och himmel, och ingen plats blev funnen för dem.
Och jag såg de döda, både stora och små, stå inför tronen, och böcker blevo upplåtna.
Och jämväl en annan bok blev upplåten; det var livets bok.
Och de döda blevo dömda efter sina gärningar, på grund av det som var upptecknat i böckerna.
Och havet gav igen de döda som voro däri, och döden och dödsriket gåvo igen de döda som voro i dem; och dessa blev dömda, var och en efter sina gärningar.
Och döden och dödsriket blevo kastade i den brinnande sjön; detta, den brinnande sjön, är den andra döden.
Och om någon icke fanns skriven i livets bok, så blev han kastad i den brinnande sjön.
Och jag såg en ny himmel och en ny jord; ty den förra himmelen och den förra jorden voro förgångna, och havet fanns icke mer.
Och jag såg den heliga staden, ett nytt Jerusalem, komma ned från himmelen, från Gud, färdigsmyckad såsom en brud som är prydd för sin brudgum.
Och jag hörde en stark röst från tronen säga: »Se, nu står Guds tabernakel bland människorna, och han skall bo ibland dem, och de skola vara hans folk; ja, Gud själv skall vara hos dem
och skall avtorka alla tårar från deras ögon.
Och döden skall icke mer vara till, och ingen sorg eller klagan eller plåga skall vara mer; ty det som förr var är nu förgånget.»
Och han som satt på tronen sade: »Se, jag gör allting nytt.»
Ytterligare sade han: »Skriv: ty dessa ord äro visa och sanna.»
Han sade vidare till mig: »Det är gjort.
Jag är A och O, begynnelsen och änden.
Åt den som törstar skall jag giva att dricka för intet ur källan med livets vatten.
Den som vinner seger, han skall få detta till arvedel, och jag skall vara hans Gud, och han skall vara min son.
Men de fega och de otrogna, och de som hava gjort vad styggeligt är, och dråpare och otuktiga människor och trollkarlar och avgudadyrkare och alla lögnare skola få sin del i den sjö som brinner med eld och svavel; detta är den andra döden.»
Och en av de sju änglarna med de sju skålar, som voro fulla med de sju sista plågorna, kom och talade till mig och sade: »Kom hit, så skall jag visa dig bruden, Lammets hustru.»
Och han förde mig i anden åstad upp på ett stort och högt berg och visade mig den heliga staden Jerusalem, som kom ned från himmelen, från Gud,
med Guds härlighet.
Den glänste likt den dyrbaraste ädelsten, den var såsom kristallklar jaspis.
Den hade en stor och hög mur med tolv portar, och vid portarna stodo tolv änglar, och över portarna voro skrivna namn: namnen på Israels barns tolv stammar.
I öster voro tre portar, i norr tre portar, i söder tre portar och i väster tre portar.
Och stadsmuren hade tolv grundstenar, och på dem stodo tolv namn: namnen på Lammets tolv apostlar.
Och han som talade till mig hade en gyllene mätstång för att därmed mäta staden och dess portar och dess mur.
Och staden utgjorde en fyrkant, och dess längd var lika stor som dess bredd.
Och med stången mätte han staden: dess mått var tolv tusen stadier, dess längd och bredd och höjd voro lika.
Och han mätte dess mur: den var ett hundra fyrtiofyra alnar efter människors mått, som ock är änglars.
Och stadsmuren var byggd av jaspis, men staden själv var av rent guld, likt rent glas.
Stadsmurens grundstenar voro skönt lagda och utgjordes av alla slags ädelstenar.
Den första grundstenen var en jaspis, den andra en safir, den tredje en kalcedon, den fjärde en smaragd,
den femte en sardonyx, den sjätte en karneol, den sjunde en krysolit, den åttonde den beryll, den nionde en topas, den tionde en krysopras, den elfte en hyacint, den tolfte en ametist.
Och de tolv portarna utgjordes av tolv pärlor; var särskild port utgjordes av en enda pärla.
Och stadens gata var av rent guld, likt genomskinligt glas.
Och jag såg i den intet tempel, ty Herren Gud, den Allsmäktige, är dess tempel, han och Lammet.
Och staden behöver icke sol eller måne till att lysa där, ty Guds härlighet upplyser den och dess ljus är Lammet.
Och folken skola vandra i dess ljus, och jordens konungar föra ditin, vad härligt de hava.
Dess portar skola aldrig stängas om dagen -- natt skall icke finnas där
och vad härligt och dyrbart folken hava skall man föra ditin.
Men intet orent skall någonsin komma ditin, och ingen som gör vad styggeligt är och lögn, utan allenast de som äro skrivna i livets bok, Lammets bok.
Och han visade mig en ström med vatten, klar som kristall.
Den gick ut från Guds och Lammets tron
och flöt fram mitt igenom stadens gata.
Och på båda sidor om strömmen stodo livsträd, som gåvo tolv skördar, ty de buro frukt var månad; och trädens löv tjänade till läkedom för folken.
Och ingen förbannelse skall vara mer.
Och Guds och Lammets tron skall stå där inne, och hans tjänare skall tjäna honom
och skola se hans ansikte; och hans namn skall stå tecknat på deras pannor.
Och ingen natt skall vara mer; och de behöva icke någon lampas ljus, ej heller solens ljus, ty Herren Gud skall lysa över dem, och de skola regera i evigheternas evigheter.
Och han sade till mig: »Dessa ord äro vissa och sanna; och Herren, profeternas andars Gud, har sänt sin ängel för att visa sina tjänare, vad som snart skall ske.
Och se, jag kommer snart.
Salig är den som tager vara på de profetians ord som stå i denna bok.»
Och jag, Johannes, var den som hörde och såg detta.
Och när jag hade hört och sett det, föll jag ned för att tillbedja inför ängelns fötter, hans som visade mig detta.
Men han sade till mig: »Gör icke så.
Jag är din medtjänare och dina bröders, profeternas, och deras som taga vara på denna boks ord.
Gud skall du tillbedja.»
Och han sade till mig: »Göm icke under något insegel de profetians ord som stå i denna bok; ty tiden är nära.
Må den som är orättfärdig fortfara att öva sin orättfärdighet och den som är oren att orena sig.
Så ock den som är rättfärdig, han fortfare att öva sin rättfärdighet, och den som är helig att helga sig.
Se, jag kommer snart och har med mig min lön, för att vedergälla var och en efter som hans gärningar äro.
Jag är A och O, den förste och den siste, begynnelsen och änden.
Saliga äro de som två sina kläder för att få rätt att äta av livets träd och att gå in i staden genom dess portar.
Men de som äro hundar och trollkarlar och otuktiga och dråpare och avgudadyrkare och alla som älska och göra lögn, de måste alla stanna därutanför.»
Jag, Jesus, har sänt min ängel för att i församlingarna vittna om detta för eder.
Jag är telningen från Davids rot och kommen av hans släkt, jag är den klara morgonstjärnan.
Och Anden och bruden säga: »Kom.»
Och den som hör det, han säge »Kom.»
Och den som törstar, han komme; ja den som vill, han tage livets vatten för intet.
För var och en som hör de profetians ord, som stå i denna bok betygar jag detta: »Om någon lägger något till dem, så skall Gud på honom lägga de plågor om vilka är skrivet i denna bok.
Och om någon tager bort något från de ord som stå i denna profetias bok, så skall Gud taga ifrån honom hans del i livets träd och i den heliga staden, om vilka är skrivet i denna bok.»
Han som betygar detta säger: »Ja, jag kommer snart.»
Amen.
Kom Herre Jesus!
Herren Jesu nåd vare med alla.