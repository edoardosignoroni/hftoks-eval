Josua, Nuns son, som hade varit Moses tjänare allt ifrån sin ungdom, tog då till orda och sade: »Mose, min herre, förbjud dem det.»
Men Mose sade till honom: »Skall du så nitälska för mig?
Ack att fastmer allt HERRENS folk bleve profeter, därigenom att HERREN läte sin Ande komma över dem!»
Sedan gick Mose tillbaka till lägret med de äldste i Israel.
Och en stormvind for ut ifrån HERREN, och den förde med sig vaktlar från havet och drev dem över lägret, en dagsresa vitt på vardera sidan, runt omkring lägret, och vid pass två alnar högt över marken.
Då stod folket upp och gick hela den dagen och sedan hela natten och hela den följande dagen och samlade ihop vaktlar; det minsta någon samlade var tio homer.
Och de bredde ut dem runt omkring lägret.
Men under det att de ännu hade köttet mellan tänderna, innan det var förtärt, upptändes HERRENS vrede mot folket, och HERREN anställde ett mycket stort nederlag bland folket.
Och detta ställe fick namnet Kibrot-Hattaava, ty där begrov man dem av folket, som hade gripits av lystnad.
Från Kibrot-Hattaava bröt folket upp och tågade till Haserot; och i Haserot stannade de.
Och Mirjam jämte Aron talade illa om Mose för den etiopiska kvinnans skull som han hade tagit till hustru; han hade nämligen tagit en etiopisk kvinna till hustru.
Och de sade: »Är då Mose den ende som HERREN talar med?
Talar han icke också med oss?»
Och HERREN hörde detta.
Men mannen Mose var mycket saktmodig, mer än någon annan människa på jorden.
Och strax sade HERREN till Mose, Aron och Mirjam: »Gån ut, I tre, till uppenbarelsetältet.»
Och de gingo ditut, alla tre.
Då steg HERREN ned i en molnstod och blev stående vid ingången till tältet; och han kallade på Aron och Mirjam, och de gingo båda ditut.
Och han sade: »Hören nu mina ord.
Eljest om någon är en profet bland eder, giver jag, HERREN, mig till känna för honom i syner och talar med honom i drömmar.
Men så gör jag icke med min tjänare Mose; i hela mitt hus är han betrodd.
Muntligen talar jag med honom, öppet och icke i förtäckta ord, och han får skåda HERRENS gestalt.
Varför haven I då icke haft försyn för att tala illa om min tjänare Mose?»
Och HERRENS vrede upptändes mot dem, och han övergav dem.
När så molnskyn drog sig tillbaka från tältet, se, då var Mirjam vit såsom snö av spetälska; när Aron vände sig till Mirjam, fick han se att hon var spetälsk.
Då sade Aron till Mose: »Ack, min herre, lägg icke på oss bördan av en synd som vi i vår dårskap hava begått.
Låt henne icke bliva lik ett dödfött foster, vars kropp är till hälften förstörd, när det kommer ut ur sin moders liv.»
Då ropade Mose till HERREN och sade: »O Gud, gör henne åter frisk.»
HERREN svarade Mose: »Om hennes fader hade spottat henne i ansiktet, skulle hon ju hava fått sitta med skam i sju dagar.
Må hon alltså nu hållas innestängd i sju dagar utanför lägret; sedan får hon komma tillbaka dit igen.»
Så hölls då Mirjam innestängd i sju dagar utanför lägret, och folket bröt icke upp, förrän Mirjam hade kommit tillbaka.
Därefter bröt folket upp från Haserot och lägrade sig i öknen Paran.
Och HERREN talade till Mose och sade:
»Sänd åstad några män för att bespeja Kanaans land, som jag vill giva åt Israels barn.
En man ur var fädernestam skolen I sända, men allenast sådana som äro hövdingar bland dem.»
Och Mose sände från öknen Paran åstad sådana män, efter HERRENS befallning; allasammans hörde de till huvudmännen bland Israels barn.
Och dessa voro namnen på dem: Av Rubens stam: Sammua, Sackurs son;
av Simeons stam: Safat, Horis son;
av Juda stam: Kaleb, Jefunnes son;
av Isaskars stam: Jigeal, Josefs son;
av Efraims stam: Hosea, Nuns son;
av Benjamins stam: Palti, Rafus son;
av Sebulons stam: Gaddiel, Sodis son;
av Josefs stam: av Manasse stam: Gaddi, Susis son;
av Dans stam: Ammiel, Gemallis son;
av Asers stam: Setur, Mikaels son;
av Naftali stam: Nahebi, Vofsis son;
av Gads stam; Geuel, Makis son.
Dessa voro namnen på de män som Mose sände åstad för att bespeja landet.
Men Mose gav Hosea, Nuns son, namnet Josua.
Och Mose sände dessa åstad för att bespeja Kanaans land.
Och han sade till dem: »Dragen nu upp till Sydlandet, och dragen vidare upp till Bergsbygden.
Och sen efter, hurudant landet är, och om folket som bor däri är starkt eller svagt, om det är litet eller stort,
och hurudant landet är, vari de bo, om det är gott eller dåligt, och hurudana de platser äro, där de bo, om de bo i läger eller i befästa städer,
och hurudant själva landet är, om det är fett eller magert, om träd finnas där eller icke.
Varen vid gott mod, och tagen med eder hit av landets frukt.»
Det var nämligen vid den tid då de första druvorna voro mogna
Så drogo de åstad och bespejade landet från öknen Sin ända till Rehob, där vägen går till Hamat.
De drogo upp till Sydlandet och kommo till Hebron; där bodde Ahiman, Sesai och Talmai, Anaks avkomlingar.
Men Hebron byggdes sju år före Soan i Egypten.
Och de kommo till Druvdalen; där skuro de av en kvist med en ensam druvklase på, och denna bars sedan på en stång av två man.
Därtill togo de granatäpplen och fikon.
Detta ställe blev kallat Druvdalen för den druvklases skull som Israels barn där skuro av.
Och efter fyrtio dagar vände de tillbaka, sedan de hade bespejat landet.
De gingo åstad och kommo till Mose och Aron och Israels barns hela menighet i öknen Paran, i Kades, och avgåvo sin berättelse inför dem och hela menigheten och visade dem landets frukt.
De förtäljde för honom och sade: »Vi kommo till det land dit du sände oss.
Och det flyter i sanning av mjölk och honung, och här är dess frukt.
Men folket som bor i landet är starkt, och städerna äro välbefästa och mycket stora; ja, vi sågo där också avkomlingar av Anak.
Amalekiterna bo i Sydlandet, hetiterna, jebuséerna och amoréerna bo i Bergsbygden, och kananéerna bo vid havet och utmed Jordan.»
Men Kaleb sökte stilla folket, så att de icke skulle knota emot Mose; han sade: »Låt oss ändå draga ditupp och intaga det, ty förvisso skola vi bliva det övermäktiga.»
Men de män som hade varit däruppe med honom sade: »Vi kunna icke draga upp mot detta folk, ty de äro oss för starka.»
Och de talade bland Israels barn illa om landet som de hade bespejat; de sade: »Det land som vi hava genomvandrat och bespejat är ett land som förtär sina inbyggare, och alla människor, som vi där sågo, voro resligt folk.
Vi sågo där ock jättarna, Anaks barn, av jättestammen; vi tyckte då att vi själva voro såsom gräshoppor, och sammalunda tyckte de om oss.
Då begynte hela menigheten ropa och skria, och folket grät den natten.
Och alla Israels barn knorrade emot Mose och Aron, och hela menigheten sade till dem: »O att vi hade fått dö i Egyptens land, eller att vi hade fått dö här i öknen!
Varför vill då HERREN föra oss in i detta andra land, där vi måste falla för svärd, och där våra hustrur och barn skola bliva fiendens byte?
Det vore förvisso bättre för oss att vända tillbaka till Egypten.»
Och de sade till varandra: »Låt oss välja en anförare och vända tillbaka till Egypten.»
Då föllo Mose och Aron ned på sina ansikten inför Israels barns hela församlade menighet.
Och Josua, Nuns son, och Kaleb, Jefunnes son, vilka voro bland dem som hade bespejat landet, revo sönder sina kläder
och sade till Israels barns hela menighet: »Det land som vi hava genomvandrat och bespejat är ett övermåttan gott land.
Om HERREN har behag till oss, så skall han föra oss in i det landet och giva det åt oss -- ett land som flyter av mjölk och honung.
Allenast mån I icke sätta eder upp mot HERREN; och för folket i landet mån I icke frukta, ty de skola bliva såsom en munsbit för oss.
Deras beskärm har vikit ifrån dem, men med oss är HERREN; frukten icke för dem.»
Men hela menigheten ropade att man skulle stena dem.
Då visade sig HERRENS härlighet i uppenbarelsetältet för alla Israels barn.
Och HERREN sade till Mose: »Huru länge skall detta folk förakta mig, och huru länge skola de framhärda i att icke vilja tro på mig, oaktat alla de tecken jag har gjort bland dem?
Jag skall slå dem med pest och förgöra dem, men dig vill jag göra till ett folk, större och mäktigare än detta.»
Mose sade till HERREN: »Egyptierna hava ju förnummit att du med din kraft har fört detta folk ut ifrån dem hitupp,
och de hava omtalat det för inbyggarna här i landet, så att de hava fått höra att du är HERREN mitt ibland detta folk, att du, HERRE, visar dig för dem ansikte mot ansikte, att din molnsky står över dem, och att du går framför dem i en molnstod om dagen och i en eldstod om natten.
Om du nu dödade detta folk, alla tillsammans, då skulle hedningarna, som finge höra detta berättas om dig, säga så:
'Därför att HERREN icke förmådde föra detta folk in i det land som han med ed hade lovat åt dem, därför har han slaktat dem i öknen.'
Nej, må nu Herrens kraft bevisa sig stor, såsom du har talat och sagt:
'HERREN är långmodig och stor i mildhet, han förlåter missgärning och överträdelse, fastän han icke låter någon bliva ostraffad, utan hemsöker fädernas missgärning på barn och efterkommande i tredje och fjärde led.'
Så tillgiv nu detta folk dess missgärning, enligt din stora nåd, såsom du har låtit din förlåtelse följa detta folk allt ifrån Egypten och ända hit.»
Då sade HERREN: »Jag vill tillgiva dem efter din bön.
Men så sant jag lever, och så sant hela jorden skall bliva full av HERRENS härlighet:
av alla de män som hava sett min härlighet och de tecken jag har gjort i Egypten och i öknen, och som dock nu tio gånger hava frestat mig och icke velat höra min röst,
av dem skall ingen få se det land som jag med ed har lovat åt deras fäder; ingen av dem som hava föraktat mig skall få se det.
Men eftersom i min tjänare Kaleb är en annan ande, så att han i allt har efterföljt mig, därför vill jag låta honom komma in i det land där han nu har varit, och hans avkomlingar skola besitta det.
Men då nu amalekiterna och kananéerna bo i dalbygden, så vänden eder i morgon åt annat håll bryten upp och tagen vägen mot öknen, åt Röda havet till.»
Och HERREN talade till Mose och Aron och sade:
»Huru länge skall denna onda menighet fortfara att knorra mot mig?
Ty jag har hört huru Israels barn knorra mot mig.
Säg nu till dem: 'Så sant jag lever, säger HERREN, jag skall göra med eder såsom I själva haven sagt inför mig.
Här i öknen skola edra döda kroppar bliva liggande; så skall det gå eder alla, så många I ären som haren blivit inmönstrade, alla som äro tjugu år gamla eller därutöver, eftersom I haven knorrat mot mig.
Sannerligen, ingen av eder skall komma in i det land som jag med upplyft hand har lovat giva eder till boning, ingen förutom Kaleb, Jefunnes son, och Josua, Nuns son.
Men edra barn, om vilka I saden att de skulle bliva fiendens byte? dem skall jag låta komma ditin, och de skola lära känna det land som I haven föraktat.
I själva däremot -- edra döda kroppar skola bliva liggande här i öknen.
Och edra barn skola draga omkring såsom herdar i öknen i fyrtio år, och skola bära på bördan av eder trolösa avfällighet, till dess att edra döda kroppar hava förgåtts i öknen.
Såsom I under fyrtio dagar haven bespejat landet, så skolen I under fyrtio år -- ett år för var dag -- komma att bära på edra missgärningar; I skolen då förnimma vad det är att jag tager min hand ifrån eder.'
Jag, HERREN, talar; jag skall förvisso göra så med hela denna onda menighet, som har rotat sig samman mot mig; här i öknen skola de förgås, här skola de dö.»
Och de män som Mose hade sänt åstad för att bespeja landet, och som vid sin återkomst hade förlett hela menigheten att knorra mot honom, därigenom att de talade illa om landet,
dessa män som hade talat illa om landet träffades nu av döden genom en hemsökelse, inför HERRENS ansikte.
Av de män som hade gått åstad för att bespeja landet blevo dock Josua, Nuns son, och Kaleb, Jefunnes son, vid liv.
Och Mose talade detta till alla Israels barn.
Då blev folket mycket sorgset.
Och de stodo upp bittida följande morgon för att draga åstad upp mot den övre bergsbygden; och de sade: »Se, här äro vi; vi vilja nu draga upp till det land som HERREN har talat om; ty vi hava syndat.»
Men Mose sade: »Varför viljen I så överträda HERRENS befallning?
Det kan ju icke lyckas väl.
HERREN är icke med bland eder; dragen därför icke ditupp, på det att I icke mån bliva slagna av edra fiender.
Ty amalekiterna och kananéerna skola där möta eder, och I skolen falla för svärd; I haven ju vänt eder bort ifrån HERREN, och HERREN skall därför icke vara med eder.»
Likväl drogo de i sitt övermod upp mot den övre bergsbygden; men HERRENS förbundsark och Mose lämnade icke lägret.
Då kommo amalekiterna och kananéerna, som bodde där i bergsbygden, ned och slogo dem och förskingrade dem och drevo dem ända till Horma.
Och HERREN talade till Mose och sade:
Tala till Israels barn och säg till dem: Om I, när I kommen in i det land som jag vill giva eder, och där I skolen bo,
viljen offra ett eldsoffer åt HERREN, ett brännoffer eller ett slaktoffer -- vare sig det gäller att fullgöra ett löfte, eller det gäller ett frivilligt offer, eller det gäller edra högtidsoffer -- för att bereda HERREN en välbehaglig lukt, genom fäkreatur eller småboskap,
så skall den som vill offra åt HERREN ett sådant offer bära fram såsom spisoffer en tiondedels efa fint mjöl, begjutet med en fjärdedels hin olja;
och såsom drickoffer skall du offra en fjärdedels hin vin till vart lamm, vare sig det är ett brännoffer som offras, eller det är ett slaktoffer.
Men till en vädur skall du såsom spisoffer offra två tiondedels efa fint mjöl, begjutet med en tredjedels hin olja,
och såsom drickoffer skall du bära fram en tredjedels hin vin, till er välbehaglig lukt för HERREN.
Och när du offrar en ungtjur till brännoffer eller till slaktoffer, vare sig det gäller att fullgöra ett löfte eller det gäller tackoffer åt HERREN.
Så skall, jämte ungtjuren, såsom spisoffer frambäras tre tiondedels efa fint mjöl, begjutet med en halv in olja,
och såsom drickoffer skall du bära fram en halv hin vin: ett eldsoffer till en välbehaglig lukt för HERREN.
Vad här är sagt skall offras till var tjur, var vädur, vart djur av småboskapen, vare sig får eller get.
Efter antalet av de djur I offren skolen I offra till vart och ett vad här är sagt, efter deras antal.
Var inföding skall offra detta, såsom här är sagt, när han vill offra ett eldsoffer till en välbehaglig lukt för HERREN.
Och när en främling som vistas hos eder, eller som i kommande släkten bor ibland eder, vill offra ett eldsoffer till en välbehaglig lukt för HERREN, så skall han offra på samma sätt som I offren.
Inom församlingen skall en och samma stadga gälla för eder och för främlingen som bor ibland eder.
Detta skall vara en evärdlig stadga för eder från släkte till släkte: I själva och främlingen skolen förfara på samma sätt inför HERRENS ansikte.
Samma lag och samma rätt skall gälla för eder och för främlingen som bor hos eder.
Och HERREN talade till Mose och sade:
Tala till Israels barn och säg till dem: När I kommen in i det land dit jag vill föra eder,
skolen I, då I äten av landets bröd, giva åt HERREN en offergärd därav.
Såsom förstling av edert mjöl skolen I giva en kaka till offergärd; I skolen giva den, likasom I given en offergärd från eder loge.
Av förstlingen av edert mjöl skolen I giva åt HERREN en offergärd, släkte efter släkte.
Och om I begån synd ouppsåtligen, i det att I underlåten att göra efter något av dessa bud som HERREN har kungjort för Mose,
efter något av det som HERRENS har bjudit eder genom Mose, från den dag då HERREN gav sina bud och allt framgent, släkte efter släkte,
så skall, om synden har blivit begången ouppsåtligen, utan att menigheten visste det, hela menigheten offra en ungtjur såsom brännoffer, till en välbehaglig lukt för HERREN, med det spisoffer och det drickoffer som på föreskrivet sätt skall offras därtill, och tillika en bock såsom syndoffer.
Och prästen skall bringa försoning för Israels barns hela menighet, och så bliver dem förlåtet; ty det var en ouppsåtlig synd, och de hava burit fram sitt offer, ett eldsoffer åt HERREN, och sitt syndoffer inför HERRENS ansikte för sin ouppsåtliga synd.
Ja, så bliver dem förlåtet, Israels barns hela menighet och främlingen som bor ibland dem; ty hela folket var delaktigt i den ouppsåtliga synden.
Och om någon enskild syndar ouppsåtligen, skall han såsom syndoffer föra fram en årsgammal get.
Och prästen skall bringa försoning för denne som har försyndat sig genom ouppsåtlig synd, inför HERRENS ansikte; på det att honom må bliva förlåtet, när försoning bringas för honom.
För infödingen bland Israels barn och för främlingen som bor ibland dem, för eder alla skall gälla en och samma lag, när någon begår synd ouppsåtligen.
Men den som begår något med upplyft hand, evad han är inföding eller främling, han hånar HERREN, och han skall utrotas ur sitt folk.
Ty HERRENS ord har han föraktat, och mot hans bud har han brutit; utan förskoning skall han utrotas; missgärning vilar på honom.
Medan nu Israels barn voro i öknen, ertappades en man med att samla ihop ved på sabbatsdagen.
Och de som ertappade honom med att samla ihop ved förde honom fram inför Mose och Aron och hela menigheten.
Och då det icke var bestämt vad som borde göras med honom, satte de honom i förvar.
Och HERREN sade till Mose: »Mannen skall straffas med döden; hela menigheten skall stena honom utanför lägret.»
Då förde hela menigheten ut honom utanför lägret och stenade honom till döds, såsom HERREN hade bjudit Mose.
Och HERREN talade till Mose och sade:
Tala till Israels barn och säg till dem att de och deras efterkommande skola göra sig tofsar i hörnen på sina kläder och sätta ett mörkblått snöre på var hörntofs.
Och detta skolen I hava till tofsprydnad, för att I, när I sen därpå, mån tänka på alla HERRENS bud och göra efter dem, och icke sväva omkring efter edra hjärtans och ögons lustar, som I nu löpen efter i trolös avfällighet.
Ty jag vill att I skolen tänka på och göra efter alla mina bud och vara helgade åt eder Gud.
Jag är HERREN, eder Gud, som har fört eder ut ur Egyptens land, för att jag skall vara eder Gud Jag är HERREN, eder Gud.
Och Kora, son till Jishar, son till Kehat, son till Levi, samt Datan och Abiram, Eliabs söner, och On, Pelets son, av Rubens söner, dessa togo till sig folk
och gjorde uppror emot Mose; och dem följde två hundra femtio män av Israels barn, hövdingar i menigheten, ombud i folkförsamlingen, ansedda män.
Och de församlade sig emot Mose och Aron och sade till dem: »Nu må det vara nog.
Hela menigheten är ju helig, alla äro det, och HERREN är mitt ibland dem; varför upphäven I eder då över HERRENS församling?»
När Mose hörde detta, föll han ned på sitt ansikte.
Sedan talade han till Kora och hela hans hop och sade: »I morgon skall HERREN göra kunnigt vem som hör honom till, och vem som är den helige åt vilken han giver tillträde till sig.
Och den han utväljer, honom skall han giva tillträde till sig.
Gören nu på detta sätt: tagen edra fyrfat, du Kora och hela din hop,
och läggen eld i dem och strön rökelse på dem inför HERRENS ansikte i morgon; den man som HERREN då utväljer, han är den helige.
Ja, nu må det vara nog, I Levi söner.»
Ytterligare sade Mose till Kora: Hören nu, I Levi söner.
Är det eder icke nog att Israels Gud har avskilt eder från Israels menighet och givit eder tillträde till sig, så att I fån förrätta tjänsten i HERRENS tabernakel och stå inför menigheten och betjäna den?
Åt dig, och åt alla dina bröder, Levi söner, jämte dig, har han givit tillträde till sig; och nu stån I också efter prästadömet!
Därför, tagen eder till vara, du och hela din hop, I som haven rotat eder samman mot HERREN -- ty vad är Aron, att I knorren mot honom?»
Och Mose sände och lät kalla till sig Datan och Abiram, Eliabs söner.
Men de sade: »vi komma icke.
Är det icke nog att du har fört oss hitupp ur ett land som flöt av mjölk och honung, för att låta oss dö I öknen?
Vill du nu ock upphäva dig till herre över oss?
Ingalunda har du fört oss in i ett land som flyter av mjölk och honung, eller givit oss åkrar och vingårdar till arvedel.
Eller tror du att du kan sticka ut ögonen på dessa människor?
Nej, vi komma icke.»
Då blev Mose mycket vred och sade till HERREN: »Se icke till deras offergåva.
Icke så mycket som en enda åsna har jag tagit av dem, och ingen av dem har jag gjort något ont.»
Och Mose sade till Kora: »Du och hela din hop mån inställa eder inför HERRENS ansikte i morgon, du själv och de, så ock Aron.
Och var och en av eder må taga sitt fyrfat och lägga rökelse därpå, och sedan bära sitt fyrfat fram inför HERRENS ansikte, två hundra femtio fyrfat; du själv och Aron mån ock taga var sitt fyrfat.»
Och de togo var och en sitt fyrfat och lade eld därpå och strödde rökelse därpå, och ställde sig vid ingången till uppenbarelsetältet; och Mose och Aron likaså.
Och Kora församlade mot dem hela menigheten vid ingången till uppenbarelsetältet.
Då visade sig HERRENS härlighet för hela menigheten.
och HERREN talade till Mose och Aron och sade:
»Skiljen eder från denna menighet, så skall jag i ett ögonblick förgöra dem.»
Då föllo de ned på sina ansikten och sade: »O Gud, du Gud som råder över allt kötts anda, skall du förtörnas på hela menigheten, därför att en enda man syndar?»
Då talade HERREN till Mose och sade:
»Tala till menigheten och säg: Dragen eder bort ifrån platsen runt omkring Koras, Datans och Abirams lägerställe.»
Och Mose stod upp och gick till Datan och Abiram, och de äldste i Israel följde honom.
Och han talade till menigheten och sade: »Viken bort ifrån dessa ogudaktiga människors tält, och kommen icke vid något som tillhör dem, på det att I icke mån förgås genom alla deras synder.»
Då drogo de sig bort ifrån platsen runt omkring Koras, Datans och Abirams lägerställe; men Datan och Abiram hade gått ut och ställt sig vid ingången till sina tält med sina hustrur och barn, både stora och små.
Och Mose sade: »Därav skolen I förnimma att det är HERREN som har sänt mig för att göra alla dessa gärningar, och att jag icke har handlat efter eget tycke:
om dessa dö på samma sätt som andra människor dö, eller drabbas av hemsökelse på samma sätt som andra människor, så har HERREN icke sänt mig;
men om HERREN här låter något alldeles nytt ske, i det att marken öppnar sin mun och uppslukar dem med allt vad de hava, så att de levande fara ned i dödsriket, då skolen I därav veta att dessa människor hava föraktat HERREN.»
Och just som han hade slutat att tala allt detta, rämnade marken under dem,
och jorden öppnade sin mun och uppslukade dem och deras hus och allt Koras folk och alla deras ägodelar;
och de foro levande ned i dödsriket, de med allt vad de hade, och jorden övertäckte dem, och så utrotades de ur församlingen.
Och hela Israel, som stod runt omkring dem, flydde vid deras rop, ty de fruktade att bliva uppslukade av jorden.
Men eld gick ut från HERREN och förtärde de två hundra femtio männen som hade burit fram rökelse.
Och HERREN talade till Mose och sade:
»Säg till Eleasar, prästen Arons son, att han skall taga fyrfaten ut ur branden, men kasta ut elden i dem långt bort,
ty de hava blivit heliga.
Och dessa fyrfat -- de mäns som genom sin synd förverkade sina liv -- dem skall man hamra ut till plåtar för att därmed överdraga altaret; ty de hava varit framburna inför HERRENS ansikte och hava därigenom blivit heliga.
Och de skola så vara ett tecken för Israels barn.»
Då tog prästen Eleasar kopparfyrfaten som de uppbrända männen hade burit fram, och man hamrade ut dem för att därmed överdraga altaret,
till en påminnelse för Israels barn att ingen främmande, ingen som icke vore av Arons säd, måtte träda fram för att antända rökelse inför HERRENS ansikte, på det att det icke skulle gå honom såsom det gick Kora och hans hop: allt i enlighet med vad HERREN hade sagt honom genom Mose.
Men dagen därefter knorrade Israels barns hela menighet emot Mose och Aron och sade: »Det är I som haven dödat HERRENS folk.»
Då nu menigheten församlade sig emot Mose och Aron, vände dessa sig mot uppenbarelsetältet och fingo då se molnskyn övertäcka det; och HERRENS härlighet visade sig.
Då gingo Mose och Aron fram inför uppenbarelsetältet.
Och HERREN talade till Mose och sade:
»Gån bort ifrån denna menighet, så skall jag i ett ögonblick förgöra dem.»
Då föllo de ned på sina ansikten.
Och Mose sade till Aron: »Tag ditt fyrfat och lägg eld från altaret därpå och strö rökelse därpå, och bär det så med hast bort till menigheten och bringa försoning för dem; ty förtörnelse har gått ut från HERRENS ansikte, och hemsökelsen har begynt.»
Då tog Aron det som Mose hade tillsagt honom och skyndade mitt in i församlingen, och se, hemsökelsen hade redan begynt ibland folket, men han lade rökelsen på och bragte försoning för folket.
När han så stod mellan de döda och de levande, upphörde hemsökelsen.
Men de som hade omkommit genom hemsökelsen utgjorde fjorton tusen sju hundra, förutom dem som hade omkommit för Koras skull.
Sedan vände Aron tillbaka till Mose vid uppenbarelsetältets ingång; och hemsökelsen hade upphört.
Och HERREN talade till Mose och sade:
»Tala till Israels barn, och tag av dem, av alla som bland dem äro hövdingar för stamfamiljer, en stav för var stamfamilj, tillsammans tolv stavar.
Vars och ens namn skall du skriva på hans stav.
Och Arons namn skall du skriva på Levi stav; ty huvudmannen för denna stams familjer skall hava sin särskilda stav.
Sedan skall du lägga in dem i uppenbarelsetältet framför vittnesbördet, där jag uppenbarar mig för eder.
Då skall ske att den man som jag utväljer, hans stav skall grönska.
Och så skall jag göra slut på Israels barns knorrande, så att jag slipper höra huru de knorra mot eder.»
Och Mose talade till Israels barn, och hövdingarna för deras stamfamiljer gåvo honom alla var och en sin stav, tillsammans tolv stavar; och Arons stav var med bland deras stavar.
Och Mose lade stavarna inför HERRENS ansikte i vittnesbördets tält.
När nu Mose dagen därefter gick in i vittnesbördets tält, se, då grönskade Arons stav, som var där för Levi hus, den hade knoppar och utslagna blommor och mogna mandlar.
Och Mose bar alla stavarna ut från HERRENS ansikte till alla Israels barn; och de sågo på dem och togo var och en sin stav.
Och HERREN sade till Mose: »Lägg Arons stav tillbaka framför vittnesbördet, för att den där må förvaras såsom ett tecken för de gensträviga; så skall du göra en ände på deras knorrande, så att jag slipper höra det, på det att de icke må dö.»
Och Mose gjorde så; såsom HERREN hade bjudit honom, så gjorde han.
Och Israels barn ropade till Mose: »Se, vi omkomma, vi förgås, vi förgås allasammans!
Var och en som kommer därvid, som kommer vid HERRENS tabernakel, han dör.
Skola vi då verkligen alla omkomma?»
Och HERREN sade till Aron: Du och dina söner, och din faders hus jämte dig, skolen bära den missgärning som vidlåder helgedomen; och du och dina söner jämte dig skolen bära den missgärning som vidlåder edert prästämbete.
Men också dina fränder, Levi stam, din faders stam, skall du låta få tillträde dit jämte dig, och de skola hålla sig till dig och betjäna dig, under det att du och dina söner jämte dig gören tjänst inför vittnesbördets tält.
Och de skola iakttaga vad du har att iakttaga, och vad som eljest är att iakttaga vid hela tältet; men de må icke komma vid de heliga redskapen eller altaret, på det att icke både de och I mån dö.
De skola hålla sig till dig och iakttaga vad som är att iakttaga vid uppenbarelsetältet, under all tjänstgöring vid tältet; men ingen främmande får komma eder nära.
Och I skolen iakttaga vad som är att iakttaga vid helgedomen och vid altaret, på det att icke förtörnelse åter må komma över Israels barn.
Se, jag har uttagit edra bröder, leviterna, bland Israels barn; en gåva äro de åt eder, givna åt HERREN, till att förrätta tjänsten vid uppenbarelsetältet.
Men du och dina söner jämte dig skolen iakttaga vad som hör till edert prästämbete, i allt vad som angår altaret och det som är innanför förlåten, och skolen så göra tjänst.
Jag giver eder edert prästämbete såsom en gåvotjänst; men om någon främmande kommer därvid, skall han dödas.
Och HERREN talade till Aron: Se, jag giver åt dig vad som skall förvaras av det som gives mig såsom gärd.
Av Israels barns alla heliga gåvor giver jag detta till ämbetslott åt dig och dina söner, såsom en evärdlig rätt.
Detta skall tillhöra dig av det! högheliga som icke lämnas åt elden: alla deras offergåvor, så ofta de frambära spisoffer eller syndoffer, eller frambära skuldoffer till ersättning åt mig, detta skall såsom högheligt tillhöra dig och dina söner.
På en höghelig plats skall du äta detta; allt mankön må äta det, det skall vara dig heligt.
Och detta är rad som skall tillhöra dig såsom en gärd av Israels barns gåvor, så ofta de frambära viftoffer; åt dig och åt dina söner och döttrar jämte dig giver jag det till en evärdlig rätt; var och en i ditt hus som är ren må äta det:
allt det bästa av olja och allt det bästa av vin och av säd, förstlingen därav, som de giva åt HERREN, detta giver jag åt dig.
Förstlingsfrukterna av allt som växer i deras land, vilka de bära fram åt HERREN, skola tillhöra dig; var och en i ditt hus som är ren må äta därav.
Allt tillspillogivet i Israel skall tillhöra dig.
Allt det som öppnar moderlivet, vad kött det vara må, evad det är människor eller boskap som de föra fram till HERREN, det skall tillhöra dig; dock så, att du tager lösen för det som är förstfött bland människor, och likaledes tager lösen för det som är förstfött bland orena djur.
Och vad angår dem som skola lösas, skall du taga lösen för dem, när de äro en månad gamla, och detta efter det värde du har bestämt: fem siklar silver, efter helgedomssikelns vikt, denna räknad till tjugu gera.
Men för det som är förstfött bland fäkreatur eller får eller getter må du icke taga lösen; det är heligt.
Deras blod skall du stänka på altaret, och deras fett skall du förbränna såsom ett eldsoffer, till en välbehaglig lukt för HERREN.
Men deras kött skall tillhöra dig; det skall tillhöra dig likasom viftoffersbringan och det högra lårstycket.
Alla heliga gåvor som Israels barn giva åt HERREN såsom gärd, dem giver jag åt dig och åt dina söner och döttrar jämte dig, såsom en evärdlig rätt.
Ett evärdligt saltförbund inför HERRENS ansikte skall detta vara för dig och för dina avkomlingar jämte dig.
och HERREN sade till Aron: I deras land skall du icke hava någon arvedel, och du skall icke hava någon lott bland dem; jag skall vara din lott och arvedel bland Israels barn.
Och se, åt Levi barn giver jag all tionde i Israel till arvedel, såsom lön för den tjänst de förrätta, tjänsten vid uppenbarelsetältet.
Men de övriga israeliterna må hädanefter icke komma vid uppenbarelsetältet, ty de skola därigenom komma att bära på synd och så träffas av döden;
utan leviterna skola förrätta tjänsten vid uppenbarelsetältet, och de skola bära de missgärningar som begås.
Detta skall vara en evärdlig stadga för eder från släkte till släkte; bland Israels barn skola de icke hava någon arvedel.
Ty den tionde som Israels barn giva åt HERREN såsom gärd, den giver jag åt leviterna till arvedel.
Därför är det som jag säger om dem att de icke skola hava någon arvedel bland Israels barn.
Och HERREN talade till Mose och sade:
Till leviterna skall du så tala och säga: När I av Israels barn mottagen den tionde som jag har bestämt att I skolen få av dem såsom eder arvedel, då skolen I därav giva en gärd åt HERREN, en tionde av tionden.
Och denna eder gärd skall så anses, som när andra giva säd från logen och vin och olja från pressen.
På detta sätt skolen ock I av all tionde som I mottagen av Israels barn giva en gärd åt HERREN; och denna HERRENS gärd av tionden skolen I giva åt prästen Aron.
Av alla gåvor som I fån skolen giva åt HERREN hela den gärd som tillkommer honom; av allt det bästa av gåvorna skolen I giva den, sådant bland dessa som passar till heliga gåvor.
Och du skall säga till dem: När I nu given såsom gärd det bästa av dem, skall denna leviternas gåva så anses, som när andra giva vad loge och press avkasta.
I med edert husfolk mån äta det på vilken plats som helst; ty det är eder lön för eder tjänstgöring vid uppenbarelsetältet.
När I så given det bästa av dem såsom gärd, skolen I icke för deras skull komma att bära på synd; och då skolen I icke ohelga Israels barns heliga gåvor och så träffas av döden.
Och HERREN talade till Mose och Aron och sade:
Detta är den lagstadga som HERREN har påbjudit: Säg till Israels barn att de skaffa fram till dig en röd, felfri ko, en som icke har något lyte, och som icke har burit något ok.
Denna skolen I lämna åt prästen Eleasar; och man skall föra ut henne utanför lägret och slakta henne i hans åsyn.
Och prästen Eleasar skall taga något av hennes blod på sitt finger, och stänka med hennes blod sju gånger mot framsidan av uppenbarelsetältet.
Sedan skall man bränna upp kon inför hans ögon; hennes hud och kött och blod jämte hennes orenlighet skall man bränna upp.
Och prästen skall taga cederträ, isop och rosenrött garn och kasta det i elden vari kon brännes upp.
Och prästen skall två sina kläder och bada sin kropp i vatten; därefter får han gå in i lägret.
Dock skall prästen vara oren ända till aftonen.
Också den som brände upp henne skall två sina kläder i vatten och bada sin kropp i vatten, och vara oren ända till aftonen.
Och en man som är ren skall samla ihop askan efter kon och lägga den utanför lägret på en ren plats.
Den skall förvaras åt Israels barns menighet, till stänkelsevatten.
Det är ett syndoffer.
Och mannen som samlade ihop askan efter kon skall två sina kläder och vara oren ända till aftonen.
Detta skall vara en evärdlig stadga för Israels barn och för främlingen som bor ibland dem.
Den som kommer vid någon död, vid en människas lik, han skall vara oren i sju dagar.
Han skall rena sig härmed på tredje dagen och på sjunde dagen, så bliver han ren.
Men om han icke renar sig på tredje dagen och på sjunde dagen, så bliver han icke ren.
Var och en som kommer vid någon död, vid liket av en människa som har dött, och sedan icke renar sig, han orenar HERRENS tabernakel, och han skall utrotas ur Israel.
Därför att stänkelsevatten icke har blivit stänkt på honom, skall han vara oren; orenhet låder alltjämt vid honom.
Detta är lagen: När en människa dör i ett tält, skall var och en som kommer in i tältet och var och en som redan är i tältet vara oren i sju dagar.
Och alla öppna kärl, alla som icke hava stått överbundna, skola vara orena.
Och var och en som ute på marken kommer vid någon som har fallit för svärd eller på annat sätt träffats av döden, eller vid människoben eller vid en grav, han skall vara oren i sju dagar.
Och för att rena den som så har blivit oren skall man taga av askan efter det uppbrända syndoffret och gjuta friskt vatten därpå i ett kärl.
Och en man som är ren skall taga isop och doppa i vattnet och stänka på tältet och på allt bohaget, och på de personer som hava varit därinne, och på honom som har kommit vid benen eller vid den fallne eller vid den som har dött på annat sätt, eller vid graven.
Och mannen som är ren skall på tredje dagen och på sjunde dagen bestänka den som har blivit oren.
När så på sjunde dagen hans rening är avslutad, skall han två sina kläder och bada sig i vatten, så bliver han ren om aftonen.
Men om någon har blivit oren och sedan icke renar sig, skall han utrotas ur församlingen; ty han har orenat HERRENS helgedom; stänkelsevatten har icke blivit stänkt på honom, han är oren.
Och detta skall vara för dem en evärdlig stadga.
Mannen som stänkte stänkelsevattnet skall två sina kläder; och om någon annan kommer vid stänkelsevattnet, skall han vara oren ända till aftonen.
Och allt som den orene kommer vid skall vara orent, och den som kommer vid honom skall vara oren ända till aftonen.
Och Israels barn, hela menigheten, kommo in i öknen Sin i den första månaden, och folket stannade i Kades; där dog Mirjam och blev där också begraven.
Och menigheten hade intet vatten; då församlade de sig emot Mose och Aron.
Och folket begynte tvista med Mose och sade: »O att också vi hade fått förgås, när våra broder förgingos inför HERRENS ansikte!
Varför haven I fört HERRENS församling in i denna öken, så att vi och vår boskap måste dö här?
Och varför haven I fört oss upp ur Egypten och låtit oss komma till denna svåra plats, där varken säd eller fikonträd eller vinträd eller granatträd växa, och där intet vatten finnes att dricka?»
Men Mose och Aron gingo bort ifrån församlingen till uppenbarelsetältets ingång och föllo ned på sina ansikten.
Då visade sig HERRENS härlighet för dem.
Och HERREN talade till Mose och sade:
»Tag staven, och församla menigheten, du med din broder Aron, och talen till klippan inför deras ögon, så skall den giva vatten ifrån sig; så skaffar du fram vatten åt dem ur klippan och giver menigheten och dess boskap att dricka.
Då tog Mose stav en från dess plats inför HERRENS ansikte, såsom han hade bjudit honom.
Och Mose och Aron sammankallade församlingen framför klippan; där sade han till dem: »Hören nu, I gensträvige; kunna vi väl ur denna klippa skaffa fram vatten åt eder?»
Och Mose lyfte upp sin hand och slog på klippan med sin stav två gånger; då kom mycket vatten ut, så att menigheten och dess boskap fick dricka.
Men HERREN sade till Mose och Aron: »Eftersom I icke trodden på mig och icke höllen mig helig inför Israels barns ögon, därför skolen I icke få föra denna församling in i det land som jag har givit dem.»
Detta var Meribas vatten, där Israels barn tvistade med HERREN, och där han bevisade sig helig på dem.
Och Mose skickade sändebud från Kades till konungen i Edom och lät säga: »Så säger din broder Israel: Du känner alla de vedermödor som vi hava haft att utstå,
huru våra fäder drogo ned till Egypten, och huru vi bodde i Egypten i lång tid, och huru vi och våra fäder blevo illa behandlade av egyptierna.
Men vi ropade till HERREN, och han hörde vår röst och sände en ängel som förde oss ut ur Egypten; och se, vi äro nu i Kades, staden som ligger vid gränsen till ditt område.
Låt oss tåga genom ditt land.
Vi skola icke taga vägen över åkrar och vingårdar, och icke dricka vatten ur brunnarna; stora vägen skola vi gå, utan att vika av vare sig till höger eller till vänster, till dess vi hava kommit igenom ditt område.»
Men Edom svarade honom: »Du får icke tåga genom mitt land.
Om du det gör, skall jag draga ut emot dig med svärd.»
Men Israels barn sade till honom: »På den allmänna farvägen skola vi draga fram, och om jag eller min boskap dricker av ditt vatten, skall jag betala det.
Jag begär ju ingenting: allenast att få tåga vägen fram härigenom.»
Han svarade: »Nej, du får icke tåga härigenom.»
Och Edom drog ut mot honom med mycket folk och ned stor makt.
Då alltså Edom icke tillstadde Israel att tåga genom sitt område, vek Israel av och gick undan för honom.
Och de bröto upp från Kades.
Och Israels barn, hela menigheten, kommo till berget Hor.
Och HERREN talade till Aron på berget Hor, vid gränsen till Edoms land, och sade:
»Aron skall samlas till sina fäder: han skall icke komma in i det land som jag har givit åt Israels barn; ty I voren gensträviga mot min befallning vid Meribas vatten.
Tag nu Aron och hans son Eleasar med dig, och för dem upp på berget Hor,
och tag av Aron hans kläder och sätt dem på hans son Eleasar.
Så skall Aron samlas till sina fäder och I dö där.»
Och Mose gjorde såsom HERREN hade bjudit; och de stego upp på berget Hor inför hela menighetens ögon.
Och Mose tog av Aron hans kläder och satte dem på hans son Eleasar.
Och Aron dog där uppe på bergets topp; men Mose och Eleasar stego ned från berget.
Och när hela menigheten förnam att Aron hade givit upp andan, begräto de honom i trettio dagar, hela Israels hus.
Då nu konungen i Arad, kananéen, som bodde i Sydlandet, hörde att Israel var i antågande på Atarimvägen, gav han sig i strid med Israel och tog några av dem till fånga.
Då gjorde Israel ett löfte åt HERREN och sade: »Om du giver detta folk i min hand, så skall jag giva deras städer till spillo.»
Och HERREN hörde Israels röst och gav kananéerna i deras hand, och de gåvo dem och deras städer till spillo; så fick stället namnet Horma.
Och de bröto upp från berget Hor och togo vägen åt Röda havet till, för att gå omkring Edoms land.
Men under vägen blev folket otåligt.
Och folket talade emot Gud och emot Mose och sade: »Varför haven I fört oss upp ur Egypten, så att vi måste dö i öknen?
Här finnes ju varken bröd eller vatten, och vår själ vämjes vid den usla föda vi få.»
Då sände HERREN giftiga ormar bland folket, och dessa stungo folket; och mycket folk i Israel blev dödat.
Då kom folket till Mose och sade: »Vi hava syndat därmed att vi talade mot HERREN och mot dig.
Bed till HERREN att han tager bort dessa ormar ifrån oss.»
Och Mose bad för folket.
Då sade HERREN till Mose: »Gör dig en orm och sätt upp den på en stång; sedan må var och en som har blivit ormstungen se på den, så skall han bliva vid liv.»
Då gjorde Mose en orm av koppar och satte upp den på en stång; när sedan någon hade blivit stungen av en orm, såg han upp på kopparormen och blev så vid liv.
Och Israels barn bröto upp och lägrade sig i Obot;
och från Obot bröto de upp och lägrade sig vid Ije-Haabarim i öknen som ligger framför Moab, österut.
Därifrån bröto de upp och lägrade sig i Sereds dal.
Därifrån bröto de upp och lägrade sig på andra sidan Arnon, där denna bäck från amoréernas område, där den har runnit upp, flyter fram i öknen; ty Arnon är Moabs gräns och flyter fram mellan Moabs land och amoréernas.
Därför heter det i »Boken om HERRENS krig»: »Vaheb i Sufa och dalarna där Arnon går fram,
och dalarnas sluttning, som sänker sig mot Ars bygd och stöder sig mot Moabs gräns.»
Därifrån drogo de till Beeri om brunnen där var det som HERREN sade till Mose: »Församla folket, så vill jag giva dem vatten.»
Då sjöng Israel denna sång: »Flöda, du brunn!
Ja, sjungen om den,
om brunnen som furstar grävde, som folkets ypperste borrade, med spiran, med sina stavar.
Från öknen drogo de till Mattana, från Mattana till Nahaliel, från: Nahaliel till Bamot,
från Bamot till den dal som ligger: på Moabs mark uppe på Pisga, där man kan se ut över ödemarken.
Och Israel skickade sändebud till Sihon, amoréernas konung, och lät säga:
»Låt mig taga genom ditt land.
Vi skola icke vika av ifrån vägen in i åkrar eller vingårdar, och icke dricka vatten ur brunnarna.
Stora vägen skola vi gå, till dess vi hava kommit igenom ditt område.»
Men Sihon tillstadde icke Israel att tåga genom sitt område, utan församlade allt sitt folk och drog ut mot Israel i öknen, till dess han kom till Jahas; där gav han sig i strid med Israel.
Men Israel slog honom med svärdsegg och intog hans land från Arnon ända till Jabbok, ända till Ammons barns land, ty Ammons barns gräns var befäst.
Och Israel intog alla städerna där; och Israel bosatte sig i amoréernas alla städer, i Hesbon och alla underlydande orter.
Hesbon var nämligen Sihons, amoréernas konungs, stad, ty denne hade fört krig med den förre konungen i Moab och tagit ifrån honom hela hans land ända till Arnon.
Därför säga skalderna: »Kommen till Hesbon!
Byggas och befästas skall Sihons stad.
Ty eld gick ut från Hesbon, en låga från Sihons stad; den förtärde Ar i Moab, dem som bodde på Arnons höjder.
Ve dig, Moab!
Förlorat är du, Kemos' folk!
Han lät sina söner bliva slagna på flykten och sina döttrar föras bort i fångenskap, bort till amoréernas konung, Sihon.
Vi sköto ned dem -- förlorat var Hesbon, landet ända till Dibon; vi härjade ända till Nofa, Nofa, som når till Medeba.»
Så bosatte sig då Israel i amoréernas land.
Och Mose sände ut och lät bespeja Jaeser, och de intogo dess underlydande orter; och han fördrev amoréerna som bodde där.
Sedan vände de sig åt annat hål. och drogo upp åt Basan till.
Och Og, konungen i Basan, drog med allt sitt folk ut till strid mot dem, till Edrei.
Men HERREN sade till Mose: »Frukta icke för honom, ty i din hand har jag givit honom och allt hans folk och hans land.
Och du skall göra med honom på samma sätt som du gjorde med Sihon, amoréernas konung, som bodde i Hesbon.»
Och de slogo honom jämte hans söner och allt hans folk, och läto ingen av dem slippa undan.
Så intogo de hans land.
Och Israels barn bröto upp och lägrade sig på Moabs hedar, på andra sidan Jordan mitt emot Jeriko.
Och Balak, Sippors son, såg allt vad Israel hade gjort mot amoréerna.
Och Moab bävade storligen för folket, därför att det var så talrikt; Moab gruvade sig för Israels barn.
Och Moab sade till de äldste i Midjan: »Nu kommer denna hop att äta upp allt som finnes här runt omkring oss, likasom oxen äter upp vad grönt som finnes på marken.»
Och Balak, Sippors son, var på den tiden konung i Moab.
Och han skickade sändebud till Bileam, Beors son, i Petor vid floden, i hans stamfränders land, för att kalla honom till sig; han lät säga: »Se, här är ett folk som har dragit ut ur Egypten; se, det övertäcker marken, och det har lägrat sig mitt emot mig.
Så kom nu och förbanna åt mig detta folk, ty det är mig för mäktigt; kanhända skall jag då kunna slå det och förjaga det ur landet.
Ty jag vet att den du välsignar, han är välsignad, och den du förbannar, han bliver förbannad.»
Så gingo nu de äldste i Moab och de äldste i Midjan åstad och hade med sig spådomslön; och de kommo till Bileam och framförde till honom Balaks ord.
Och han sade till dem: »Stannen här över natten, så vill jag sedan giva eder svar efter vad HERREN talar till mig.»
Då stannade Moabs furstar kvar hos Bileam.
Och Gud kom till Bileam; han sade: »Vad är det för män som du har hos dig?»
Bileam svarade Gud: »Balak, Sippors son, konungen i Moab, har sänt till mig detta bud:
'Se, här är det folk som har dragit ut ur Egypten, och det övertäcker marken.
Så kom nu och förbanna det åt mig; kanhända skall jag då kunna giva mig i strid med det och förjaga det.'»
Då sade Gud till Bileam: »Du skall icke gå med dem; du skall icke förbanna detta folk, ty det är välsignat.»
Om morgonen, när Bileam hade stått upp, sade han alltså till Balaks furstar: »Gån hem till edert land, ty HERREN vill icke tillstädja mig att följa med eder.»
Då stodo Moabs furstar upp och gingo hem till Balak och sade: »Bileam vägrade att följa med oss.»
Men Balak sände ännu en gång åstad furstar, flera och förnämligare än de förra.
Och de kommo till Bileam och sade till honom: »Så säger Balak Sippors son: 'Låt dig icke avhållas från att komma till mig;
ty jag vill bevisa dig övermåttan stor ära, och allt vad du begär av mig skall jag göra.
Kom nu och förbanna åt mig detta folk.'»
Då svarade Bileam och sade till Balaks tjänare: »Om Balak än gåve mig så mycket silver och guld som hans hus rymmer, kunde jag dock icke överträda HERRENS min Guds befallning, så att jag gjorde något däremot, vare sig litet eller stort.
Men stannen nu också I kvar har över natten, för att jag må förnimma vad HERREN ytterligare kan vilja tala till mig.»
Och Gud kom till Bileam om natten och sade till honom: »Om dessa män hava kommit för att kalla dig, så stå upp och följ med dem.
Men allenast vad jag säger dig skall du göra.»
Om morgonen, när Bileam hade stått upp, sadlade han alltså sin åsninna och följde med Moabs furstar.
Men då han nu följde med, upptändes Guds vrede, och HERRENS ängel ställde sig på vägen för att hindra honom, där han red på sin åsninna, åtföljd av två sina tjänare.
När då åsninnan såg HERRENS ängel stå på vägen med ett draget svärd i sin hand, vek hon av ifrån vägen och gick in på åkern; men Bileam slog åsninnan för att driva henne tillbaka in på vägen.
Därefter ställde sig HERRENS ängel i en smal gata mellan vingårdarna, där murar funnos på båda sidor.
När nu åsninnan såg HERRENS ängel, trängde hon sig mot muren och klämde så Bileams ben mot muren; och han slog henne ännu en gång.
Då gick HERRENS ängel längre fram och ställde sig på ett trångt ställe, där ingen utväg fanns att vika undan, vare sig till höger eller till vänster.
När åsninnan nu såg HERRENS ängel, lade hon sig ned under Bileam.
Då upptändes Bileams vrede och han slog åsninnan med sin stav.
Men HERREN öppnade åsninnans mun, och hon sade till Bileam: »Vad har jag gjort dig, eftersom du nu tre gånger har slagit mig?»
Bileam svarade åsninnan: »Du har ju handlat skamligt mot mig; om jag hade haft ett svärd i min hand, skulle jag nu hava dräpt dig.»
Men åsninnan sade till Bileam: »Är icke jag din egen åsninna, som du har ridit på i all din tid intill denna dag?
Och har jag någonsin förut plägat göra så mot dig?
Han svarade: »Nej.»
Och HERREN öppnade Bileams ögon, så att han såg HERRENS ängel stå på vägen med ett draget svärd i sin hand.
Då bugade han sig och föll ned på sitt ansikte.
Och HERRENS ängel sade till honom: »Varför har du nu tre gånger slagit din åsninna?
Se, jag har gått ut för att hindra dig, ty denna väg leder till fördärv och är mig emot.
Och åsninnan såg mig, och hon har nu tre gånger vikit undan for mig.
Om hon icke hade vikit undan för mig, så skulle jag nu hava dräpt dig, men låtit henne leva.»
Då sade Bileam till HERRENS ängel: »Jag har syndat, ty jag visste icke att du stod mig emot på vägen.
Om nu min resa misshagar dig, så vill jag vända tillbaka.»
Men HERRENS ängel svarade Bileam: »Följ med dessa män; men intet annat än vad jag säger dig skall du tala.»
Så följde då Bileam med Balaks furstar.
När Balak hörde att Bileam kom, gick han honom till mötes till Ir i Moab, vid gränsen där Arnon flyter, vid yttersta gränsen.
Och Balak sade till Bileam: »Sände jag icke enträget bud till dig för att kalla dig hit?
Varför ville du då icke begiva dig till mig?
Skulle jag icke kunna bevisa dig tillräcklig ära?»
Bileam svarade Balak: »Du ser nu att jag har kommit till dig.
Men det står ingalunda i min egen makt att tala något.
Vad Gud lägger i min mun, det måste jag tala.»
Sedan följde Bileam med Balak, och de kommo till Kirjat-Husot.
Och Balak slaktade fäkreatur och småboskap och sände till Bileam och de furstar som voro med honom.
Och följande morgon tog Balak Bileam med sig och förde honom upp på Bamot-Baal; och han kunde från denna plats se en del av folket.
Och Bileam sade till Balak: »Bygg här åt mig sju altaren, och skaffa hit åt mig sju tjurar och sju vädurar.»
Balak gjorde såsom Bileam sade; och Balak och Bileam offrade en tjur och en vädur på vart altare
Därefter sade Bileam till Balak »Stanna kvar vid ditt brännoffer; jag vill gå bort och se om till äventyrs HERREN visar sig för mig; och vad helst han uppenbarar för mig, det skall jag förkunna för dig.»
Och han gick upp på en kal höjd.
Och Gud visade sig för Bileam; då sade denne till honom: »De sju altarna har jag uppfört, och på vart altare har jag offrat en tjur och en vädur.»
Och HERREN lade i Bileams mun vad han skulle tala; han sade: »Gå tillbaka till Balak och tala så och så.»
När han nu kom tillbaka till honom, fann han honom stående vid sitt brännoffer tillsammans med alla Moabs furstar.
Då hör han upp sin röst och kvad: »Från Aram hämtade mig Balak, från österns berg Moabs konung: 'Kom och förbanna åt mig Jakob, kom och tala ofärd över Israel.
Huru kan jag förbanna den gud ej förbannar, och tala ofärd över den som HERREN ej talar ofärd över?
Från klippornas topp ser jag ju honom, och från höjderna skådar jag honom: se, det är ett folk som bor för sig självt och icke anser sig likt andra folkslag.
Vem kan räkna Jakob, tallös såsom stoftet, eller tälja ens fjärdedelen av Israel?
Må jag få dö de rättfärdigas död, och blive mitt slut såsom deras!»
Då sade Balak till Bileam: »Vad har du gjort mot mig!
Till att förbanna mina fiender hämtade jag dig, och nu har du i stället välsignat dem.»
Men han svarade och sade: »Skulle jag då icke akta på vad HERREN lägger i min mun, och tala det?»
Och Balak sade till honom: »Följ nu med mig till ett annat ställe, varifrån du ser dem; du ser här allenast en del av dem, du ser dem icke allasammans.
Från det stället må du förbanna dem åt mig.»
Och han tog honom med sig till Väktarplanen på toppen av Pisga.
Där byggde han sju altaren och offrade en tjur och en vädur på vart altare.
Därefter sade han till Balak: »Stanna kvar har vid ditt brännoffer; jag själv vill därborta se till, om något visar sig.»
Och HERREN visade sig för Bileam och lade i hans mun vad han skulle tala; han sade: »Gå tillbaka till Balak och tala så och så.»
När han nu kom till honom, fann han honom stående vid sitt brännoffer, och Moabs furstar stodo där med honom.
Och Balak frågade honom: »Vad har HERREN talat?»
Då hov han upp sin röst och kvad: »Stå upp, Balak, och hör; lyssna till mig, du Sippors son.
Gud är icke en människa, så att han kan ljuga, icke en människoson, så att han kan ångra något.
Skulle han säga något och icke göra det, tala något och icke fullborda det?
Se, att välsigna har jag fått i uppdrag; han har välsignat, och jag kan icke rygga det.
Ofärd är icke att skåda i Jakob och olycka icke att se i Israel.
HERREN, hans Gud, är med honom, och jubel såsom mot en konung höres där.
Det är Gud som har fört dem ut ur Egypten; deras styrka är såsom vildoxars.
Ty trolldom båtar intet mot Jakob, ej heller spådom mot Israel.
Nej, nu måste sägas om Jakob och om Israel: 'Vad gör icke Gud!'
Se, det är ett folk som står upp likt en lejoninna, ett folk som reser sig likasom ett lejon.
Det lägger sig ej ned, förrän det har ätit rov och druckit blod av slagna man.»
Då sade Balak till Bileam: »Om du nu icke vill förbanna dem, så må du åtminstone icke välsigna dem.
Men Bileam svarade och sade till Balak: »Sade jag icke till dig: 'Allt vad HERREN säger, det måste jag göra'?»
Och Balak sade till Bileam: »Kom, jag vill taga dig med mig till ett annat ställe.
Kanhända skall det behaga Gud att du därifrån förbannar dem åt mig.
Och Balak tog Bileam med sig upp på toppen av Peor, där man kan se ut över ödemarken.
Och Bileam sade till Balak: »Bygg här åt mig sju altaren, och skaffa hit åt mig sju tjurar och sju vädurar.
Och Balak gjorde såsom Bileam sade; och han offrade en tjur och en vädur på vart altare.
Då nu Bileam såg att det var: HERRENS vilja att han skulle välsigna Israel, gick han icke, såsom de förra gångerna, bort och såg efter tecken, utan vände sitt ansikte mot öknen.
Och när Bileam lyfte upp sina ögon och såg Israel lägrad efter sina stammar, kom Guds Ande över honom.
Och han hov upp sin röst och kvad: »Så säger Bileam, Beors son, så säger mannen med det slutna ögat,
så säger han som hör Guds tal, han som skådar syner från den Allsmäktige, i det han sjunker ned och får sina ögon öppnade:
Huru sköna äro icke dina tält, du Jakob, dina boningar, du Israel!
De likna dalar som utbreda sig vida, de äro såsom lustgårdar invid en ström, såsom aloeträd, planterade av HERREN, såsom cedrar invid vatten.
Vatten flödar ur hans ämbar, hans sådd bliver rikligen vattnad.
Större än Agag skall hans konung vara, ja, upphöjd bliver hans konungamakt.
Det är Gud som har fört honom ut ur Egypten.
Hans styrka är såsom en vildoxes.
Han skall uppsluka de folk som stå honom emot, deras ben skall han sönderkrossa, och med sina pilar skall han genomborra dem.
Han har lagt sig ned, han vilar såsom ett lejon, såsom en lejoninna -- vem vågar oroa honom?
Välsignad vare den som välsignar dig, och förbannad vare den som förbannar dig!»
Då upptändes Balaks vrede mot Bileam, och han slog ihop händerna.
Och Balak sade till Bileam: »Till att förbanna mina fiender kallade jag dig hit, och se, du har i stället nu tre gånger välsignat dem.
Giv dig nu av hem igen.
Jag tänkte att jag skulle få bevisa dig stor ära; men se, HERREN har förmenat dig att bliva ärad.»
Bileam svarade Balak: »Sade jag icke redan till sändebuden som du skickade till mig:
'Om Balak än gåve mig så mycket silver och guld som hans hus rymmer, kunde jag dock icke överträda HERRENS befallning, så att jag efter eget tycke gjorde något, vad det vara må.'
Vad HERREN säger, det måste jag tala.
Se, jag går nu hem till mitt folk; men jag vill varsko dig om vad detta folk skall göra mot ditt folk i kommande dagar.»
Och han hov upp sin röst och kvad: »Så säger Bileam, Beors son, så säger mannen med det slutna ögat,
så säger han som hör Guds tal och har kunskap från den Högste, han som skådar syner från den Allsmäktige, i det han sjunker ned och får sina ögon öppnade:
Jag ser honom, men icke denna tid, jag skådar honom, men icke nära.
En stjärna träder fram ur Jakob, och en spira höjer sig ur Israel.
Den krossar Moabs tinningar och slår ned alla söner till Set.
Edom skall han få till besittning till besittning Seir -- sina fienders länder.
Ty Israel skall göra mäktiga ting;
ur Jakob skall en härskare komma; han skall förgöra i städerna dem som rädda sig dit.»
Och han fick se Amalek; då hov han upp sin röst och kvad: »En förstling bland folken är Amalek, men på sistone hemfaller han åt undergång.»
Och han fick se kainéerna; då hov han upp sin röst och kvad: »Fast är din boning, och lagt på klippan är ditt näste.
Likväl skall Kain bliva utrotad; ja, Assur skall omsider föra dig i fångenskap.»
Och han lov åter upp sin röst och kvad: »O ve!
Vem skall bliva vid liv, när Gud låter detta ske?
Skepp skola komma från kittéernas kust, de skola tukta Assur, tukta Eber; också han skall hemfalla åt undergång.»
Och Bileam stod upp och vände tillbaka hem; också Balak for sin väg.
Och medan Israel uppehöll sig i Sittim, begynte folket bedriva otukt med Moabs döttrar.
Dessa inbjödo folket till sina gudars offermåltider,
Och folket åt och tillbad deras gudar.
Och Israel slöt sig till Baal-Peor.
Då upptändes HERRENS vrede mot Israel.
Och HERREN sade till Mose: »Hämta folkets alla huvudman, och låt upphänga sådana i solen för HERREN, på det att HERRENS vredes glöd må vändas ifrån Israel.»
Då sade Mose till Israels domare: »Var och en av eder dräpe bland sina män dem som hava slutit sig till Baal-Peor.»
Nu kom en man av Israels barn och förde in bland sina bröder en midjanitisk kvinna, inför Moses och Israels barns hela menighets ögon, under det att dessa stodo gråtande vid ingången till uppenbarelsetältet.
När Pinehas, son till Eleasar, son till prästen Aron, såg detta, stod han upp i menigheten och tog ett spjut i sin hand
och följde efter den israelitiske mannen in i tältets sovrum och genomborrade dem båda, såväl den israelitiske mannen som ock kvinnan, i det att han stack henne genom underlivet.
Så upphörde hemsökelsen bland Israels barn.
Men de som hade omkommit genom hemsökelsen utgjorde tjugufyra tusen.
Och HERREN talade till Mose och sade:
»Pinehas, han som är son till prästen Arons son Eleasar, har avvänt min vrede från Israels barn, i det att han har nitälskat bland dem såsom jag nitälskar; därför har jag icke i min nitälskan förgjort Israels barn.
Säg fördenskull: Se, jag gör med honom ett fridsförbund;
och för honom, och för hans avkomlingar efter honom, skall detta vara ett förbund genom vilket han får ett evärdligt prästadöme, till lön för att han nitälskade för sin Gud och bragte försoning för Israels barn.»
Och den dödade israelitiske mannen, han som dödades jämte den midjanitiska kvinnan, hette Simri, Salus son, och var hövding för en familj bland simeoniterna.
Och den dödade midjanitiska kvinnan hette Kosbi, dotter till Sur; denne var stamhövding, hövding för en stamfamilj i Midjan.
Och HERREN talade till Mose och sade:
»Angripen midjaniterna och slån dem.
Ty de hava angripit eder genom de onda råd som de lade mot eder i saken med Peor och i saken med Kosbi, den midjanitiska hövdingdottern, deras syster, vilken dödades på den dag då hemsökelsen drabbade eder för Peors skull.»
Efter denna hemsökelse talade HERREN till Mose och till Eleasar, prästen Arons son, och sade:
»Räknen antalet av Israels barn, deras hela menighet, dem som äro tjugu år gamla eller därutöver, efter deras familjer, alla stridbara män i Israel.»
Och Mose och prästen Eleasar talade till dem på Moabs hedar, vid Jordan mitt emot Jeriko, och sade:
»De som äro tjugu år gamla eller därutöver skola räknas.»
Så hade ju HERREN bjudit Mose och Israels barn, dem som hade dragit ut ur Egyptens land.
Ruben var Israels förstfödde.
Rubens barn voro: Av Hanok hanokiternas släkt, av Pallu palluiternas släkt,
av Hesron hesroniternas släkt, av Karmi karmiternas släkt.
Dessa voro rubeniternas släkter.
Och de av dem som inmönstrades utgjorde fyrtiotre tusen sju hundra trettio.
Men Pallus söner voro Eliab.
Och Eliabs söner voro Nemuel, Datan och Abiram; det var den Datan och den Abiram, båda ombud för menigheten, som satte sig upp emot Mose och Aron, tillika med Koras hop, när dessa satte sig upp emot HERREN,
varvid jorden öppnade sin mun och uppslukade dem jämte Kora, vid det tillfälle då dennes hop omkom, i det att elden förtärde de två hundra femtio männen, så att de blevo till en varnagel.
Men Koras söner omkommo icke.
Simeons barn, efter deras släkter, voro: Av Nemuel nemueliternas släkt, av Jamin jaminiternas släkt, av Jakin jakiniternas släkt,
av Sera seraiternas släkt, av Saul sauliternas släkt.
Dessa voro simeoniternas släkter, tjugutvå tusen två hundra.
Gads barn, efter deras släkter, voro: Av Sefon sefoniternas släkt, av Haggi haggiternas släkt, av Suni suniternas släkt,
av Osni osniternas släkt, av Eri eriternas släkt,
av Arod aroditernas släkt, av Areli areliternas släkt.
Dessa voro Gads barns släkter, så många av dem som inmönstrades, fyrtio tusen fem hundra.
Judas söner voro Er och Onan; men Er och Onan dogo i Kanaans land.
Och Juda barn, efter deras släkter, voro: Av Sela selaniternas släkt, av Peres peresiternas släkt, av Sera seraiternas släkt.
Men Peres' barn voro: Av Hesron hesroniternas släkt, av Hamul hamuliternas släkt.
Dessa voro Juda släkter, så många av dem som inmönstrades, sjuttiosex tusen fem hundra.
Isaskars barn, efter deras släkter, voro: Av Tola tolaiternas släkt, av Puva puniternas släkt,
av Jasub jasubiternas släkt, av Simron simroniternas släkt.
Dessa voro Isaskars släkter, så många av dem som inmönstrades, sextiofyra tusen tre hundra.
Sebulons barn, efter deras släkter, voro: Av Sered serediternas släkt, av Elon eloniternas släkt, av Jaleel jaleeliternas släkt.
Dessa voro sebuloniternas släkter, så många av dem som inmönstrades, sextio tusen fem hundra.
Josefs barn, efter deras släkter voro Manasse och Efraim.
Manasse barn voro: Av Makir makiriternas släkt; men Makir födde Gilead; av Gilead kom gileaditernas släkt.
Dessa voro Gileads barn: Av Ieser ieseriternas släkt, av Helek helekiternas släkt,
av Asriel asrieliternas släkt, av Sikem sikemiternas släkt,
av Semida semidaiternas släkt och av Hefer heferiternas släkt.
Men Selofhad, Hefers son, hade inga söner, utan allenast döttrar; och Selofhads döttrar hette Mahela, Noa, Hogla, Milka och Tirsa.
Dessa voro Manasse släkter, och de av dem som inmönstrades utgjorde femtiotvå tusen sju hundra.
Dessa voro Efraims barn, efter deras släkter: Av Sutela sutelaiternas släkt, av Beker bekeriternas släkt, av Tahan tahaniternas släkt.
Men dessa voro Sutelas barn: Av Eran eraniternas släkt
Dessa voro Efraims barns släkter, så många av dem som inmönstrades trettiotvå tusen fem hundra.
Dessa voro Josefs barn, efter deras släkter.
Benjamins barn, efter deras släkter, voro: Av Bela belaiternas släkt, av Asbel asbeliternas släkt, av Ahiram ahiramiternas släkt,
av Sefufam sufamiternas släkt, av Hufam hufamiternas släkt.
Men Belas söner voro Ard och Naaman; arditernas släkt; av Naaman naamiternas släkt.
Dessa voro Benjamins barn, efter deras släkter, och de av dem som inmönstrades utgjorde fyrtiofem tusen sex hundra.
Dessa voro Dans barn, efter deras släkter: Av Suham suhamiternas släkt.
Dessa voro Dans släkter, efter deras släkter.
Suhamiternas släkter, så många av dem som inmönstrades, utgjorde tillsammans sextiofyra tusen fyra hundra.
Asers barn, efter deras släkter, voro: Av Jimna Jimnasläkten, av Jisvi jisviternas släkt, av Beria beriaiternas släkt.
Av Berias barn: Av Heber heberiternas släkt, av Malkiel malkieliternas släkt.
Och Asers dotter hette Sera.
Dessa voro Asers barns släkter, så många av dem som inmönstrades, femtiotre tusen fyra hundra.
Naftali barn, efter deras släkter, voro: Av Jaseel jaseeliternas släkt, av Guni guniternas släkt,
av Jeser jeseriternas släkt, av Sillem sillemiternas släkt.
Dessa voro Naftali släkter, efter deras släkter; och de av dem som inmönstrades utgjorde fyrtiofem tusen fyra hundra.
Dessa voro de av Israels barn som inmönstrades, sen hundra ett tusen sju hundra trettio.
Och HERREN talade till Mose och sade:
Åt dessa skall landet utskiftas till arvedel, efter personernas antal.
Åt en större stam skall du giva en större arvedel, och åt en mindre stam en mindre arvedel; åt var stam skall arvedel givas efter antalet av dess inmönstrade.
Men genom lottkastning skall landet utskiftas.
Efter namnen på sina fädernestammar skola de få sina arvedelar.
Efter lottens utslag skall var stam större eller mindre, få sin arvedel sig tillskiftad.
Och dessa voro de av Levi stam som inmönstrades, efter deras släkter: Av Gerson gersoniternas släkt av Kehat kehatiternas släkt, av Merari merariternas släkt.
Dessa voro leviternas släkter: libniternas släkt, hebroniternas släkt maheliternas släkt, musiternas släkt koraiternas släkt.
Men Kehat födde Amram.
Och Amrams hustru hette Jokebed, Levis dotter, som föddes åt Levi i Egypten; och hon födde åt Amram Aron och Mose och deras syster Mirjam.
Och åt Aron föddes Nadab och Abihu, Eleasar och Itamar.
Men Nadab och Abihu träffades av döden, när de buro fram främmande eld inför HERRENS ansikte.
Och de av dem som inmönstrades utgjorde tjugutre tusen, alla av mankön som voro en månad gamla eller därutöver.
De hade nämligen icke blivit inmönstrade bland Israels barn, eftersom icke någon arvedel var given åt dem bland Israels barn.
Dessa voro de som inmönstrades av Mose och prästen Eleasar, när dessa mönstrade Israels barn på Moabs hedar, vid Jordan mitt emot Jeriko.
Bland dessa var ingen av dem som förut hade blivit inmönstrade av Mose och prästen Aron, när dessa mönstrade Israels barn i Sinais öken,
ty om dem hade HERREN sagt: »De skola döden dö i öknen.»
Därför var ingen kvar av dem, förutom Kaleb, Jefunnes son, och Josua, Nuns son.
Och Selofhads döttrar trädde fram Selofhads, som var son till Hefer, son till Gilead, son till Makir son till Manasse, av Manasses, Josefs sons, släkter.
Och hans döttrar hette Mahela, Noa, Hogla, Milka och Tirsa.
Dessa kommo nu inför Mose och prästen Eleasar och stamhövdingarna och hela menigheten, vid ingången till uppenbarelsetältet, och sade:
»Vår fader har dött i öknen, men han var icke med i den hop som rotade sig samman mot HERREN, Koras hop, utan han dog genom egen synd, och han hade inga söner.
Icke skall nu vår faders namn utplånas ur hans släkt för det att han icke hade någon son?
Giv åt oss en besittning ibland vår faders bröder.»
och Mose bar fram deras sak inför HERREN.
Då talade HERREN till Mose och sade:
»Selofhads döttrar hava talat rätt.
Du skall giva också dem en arvsbesittning bland deras faders bröder genom att låta deras faders arvedel övergå till dem.
Och till Israels barn skall du tala och säga: När någon dör utan att efterlämna någon son, skolen I låta hans arvedel övergå till hans dotter.
Men om han icke har någon dotter, så skolen I giva hans arvedel åt hans bröder.
Har han icke heller några bröder, så skolen I giva hans arvedel åt hans faders bröder.
Men om hans fader icke har några broder, så skolen I giva hans arvedel åt närmaste blodsförvant inom hans släkt, och denne skall då taga den i besittning.»
Detta skall vara en rättsstadga för Israels barn, såsom HERREN har bjudit Mose.
Och HERREN sade till Mose: »Stig upp här på Abarimberget, så skall du få se det land som jag har givit åt Israels barn.
Men när du har sett det, skall också du samlas till dina fäder, likasom din broder Aron har blivit samlad till sina fäder;
detta därför att I, i öknen Sin, när menigheten tvistade med mig, voren gensträviga mot min befallning och icke villen hålla mig helig genom att skaffa fram vatten inför deras ögon.»
Detta gällde Meribas vatten vid Kades, i öknen Sin.
Och Mose talade till HERREN och sade:
»Må HERREN, den Gud som råder över allt kötts anda, sätta en man över menigheten,
som kan gå i spetsen för dem, när de draga ut eller vända åter, och som kan vara deras ledare och anförare, så att icke HERRENS menighet kommer att likna får som icke hava någon herde.»
HERREN svarade Mose: »Tag till dig Josua, Nuns son, ty han är en man i vilken ande är, och lägg din hand på honom.
Och för honom fram inför prästen Eleasar och hela menigheten, och insätt honom i hans ämbete inför deras ögon,
och lägg något av din värdighet på honom, för att Israels barns hela menighet må lyda honom.
Och hos prästen Eleasar skall han sedan hava att inställa sig, för att denne genom urims dom må hämta svar åt honom inför HERRENS ansikte.
Efter hans ord skola de draga ut och vända åter, han själv och alla Israels barn med honom, hela menigheten.»
och Mose gjorde såsom HERREN hade bjudit honom; han tog Josua och förde honom fram inför prästen Eleasar och hela menigheten.
Och denne lade sina händer på honom och insatte honom i hans ämbete, såsom HERREN hade befallt genom Mose.
Och HERREN talade till Mose och sade:
Bjud Israels barn och säg till dem: Mina offer, det som är min spis av mina eldsoffer, en välbehaglig lukt för mig, dem skolen I akta på, så att I offren dem åt mig på bestämd tid.
Och säg till dem: Detta är vad I skolen offra åt HERREN såsom eldsoffer: två årsgamla felfria lamm till brännoffer för var dag beständigt.
Det ena lammet skall du offra om morgonen, och det andra lammet skall du offra vid aftontiden,
och såsom spisoffer en tiondedels efa fint mjöl, begjutet med en fjärdedels hin olja av stötta oliver.
Detta är det dagliga brännoffret, som offrades på Sinai berg, till en välbehaglig lukt, ett eldsoffer åt HERREN.
Och såsom drickoffer därtill skall du offra en fjärdedels hin, till det första lammet; i helgedomen skall drickoffer av stark dryck utgjutas åt HERREN.
Det andra lammet skall du offra vid aftontiden; med likadant spisoffer och drickoffer som om morgonen skall du offra det: ett eldsoffer till en välbehaglig lukt för HERREN.
Men på sabbatsdagen skall du offra två årsgamla felfria lamm, så ock två tiondedels efa fint mjöl, begjutet med olja, såsom spisoffer, samt tillhörande drickoffer.
Detta är sabbatsbrännoffret, som skall offras var sabbat, jämte det dagliga brännoffret med tillhörande drickoffer.
Och på edra nymånadsdagar skolen I offra till brännoffer åt HERREN två ungtjurar och en vädur och sju årsgamla felfria lamm,
så ock tre tiondedels efa fint mjöl, begjutet med olja, såsom spisoffer till var tjur, två tiondedels efa fint mjöl, begjutet med olja, såsom spisoffer till väduren,
och en tiondedels efa fint mjöl begjutet med olja, såsom spisoffer till vart lamm: ett brännoffer till en välbehaglig lukt, ett eldsoffer åt HERREN.
Och de tillhörande drickoffren skola utgöras av en halv hin vin till var tjur och en tredjedels hin till väduren och en fjärdedels hin till vart lamm.
Detta är nymånadsbrännoffret, som skall offras i var och en av årets månader.
Tillika skolen I offra en bock till syndoffer åt HERREN; den skall offras jämte det dagliga brännoffret med tillhörande drickoffer.
Och i första månaden, på fjortonde dagen i månaden, är HERRENS påsk.
Och på femtonde dagen i samma månad är högtid; då skall man äta osyrat bröd, i sju dagar.
På den första dagen skall man hålla en helig sammankomst; ingen arbetssyssla skolen I då göra.
Och såsom eldsoffer, såsom brännoffer åt HERREN, skolen I offra två ungtjurar och en vädur och sju årsgamla lamm; felfria skola de vara.
Och såsom spisoffer därtill skolen I offra fint mjöl, begjutet med olja; tre tiondedels efa skolen I offra till var ungtjur och två tiondedels efa till väduren;
en tiondedels efa skall du offra till vart och ett av de sju lammen;
tillika skolen I offra en syndoffersbock till att bringa försoning för eder.
Förutom morgonens brännoffer, som utgör det dagliga brännoffret, skolen I offra detta.
Likadana offer skolen I offra var dag i sju dagar: en eldsoffersspis, till en välbehaglig lukt för HERREN.
Jämte det dagliga brännoffret skall detta offras, med tillhörande drickoffer.
Och på den sjunde dagen skolen I hålla en helig sammankomst; ingen arbetssyssla skolen I då göra.
Och på förstlingsdagen, då I bären fram ett offer av den nya grödan åt HERREN, vid eder veckohögtid, skolen I hålla en helig sammankomst; ingen arbetssyssla skolen I då göra.
Såsom brännoffer till en välbehaglig lukt för HERREN skolen I då offra två ungtjurar, en vädur, sju årsgamla lamm,
och såsom spisoffer därtill fint mjöl, begjutet med olja: tre tiondedels efa till var tjur, två tiondedels efa till väduren,
en tiondedels efa till vart och ett av de sju lammen;
tillika skolen I offra en bock till att bringa försoning för eder.
Förutom det dagliga brännoffret med tillhörande spisoffer skolen I offra detta -- felfria skola djuren vara -- och därjämte tillhörande drickoffer.
Och i sjunde månaden, på första dagen i månaden, skolen I hålla en helig sammankomst; ingen arbetssyssla skolen I då göra.
En basunklangens dag skall den vara för eder.
Såsom brännoffer till en välbehaglig lukt för HERREN skolen I då offra en ungtjur, en vädur, sju årsgamla felfria lamm,
och såsom spisoffer därtill fint mjöl, begjutet med olja: tre tiondedels efa till tjuren, två tiondedels efa till väduren
och en tiondedels efa till vart och ett av de sju lammen;
tillika skolen I offra en bock såsom syndoffer, till att bringa försoning för eder --
detta förutom nymånadsbrännoffret med tillhörande spisoffer, och förutom det dagliga brännoffret med tillhörande spisoffer, och förutom de drickoffer som på föreskrivet sätt skola offras till båda: allt till en välbehaglig lukt, ett eldsoffer åt HERREN.
På tionde dagen i samma sjunde månad skolen I ock hålla en helig sammankomst, och I skolen då späka eder; intet arbete skolen I då göra.
Och såsom brännoffer till en välbehaglig lukt för HERREN skolen I då offra en ungtjur, en vädur, sju årsgamla lamm -- felfria skola de vara --
och såsom spisoffer därtill fint mjöl, begjutet med olja: tre tiondedels efa till tjuren, två tiondedels efa till väduren,
en tiondedels efa till vart och ett av de sju lammen;
tillika skolen I offra en bock såsom syndoffer -- detta förutom försoningssyndoffret och det dagliga brännoffret med tillhörande spisoffer, och förutom de drickoffer som höra till båda.
På femtonde dagen i sjunde månaden skolen I ock hålla en helig sammankomst; ingen arbetssyssla skolen I då göra.
Då skolen I fira en HERRENS högtid, i sju dagar.
Och såsom brännoffer, såsom eldsoffer, skolen I då offra till en välbehaglig lukt för HERREN tretton ungtjurar, två vädurar, fjorton årsgamla lamm -- felfria skola de vara --
och såsom spisoffer därtill fint mjöl, begjutet med olja: tre tiondedels efa till var och en av de tretton tjurarna, två tiondedels efa till var och en av de två vädurarna,
en tiondedels efa till vart och ett av de fjorton lammen;
tillika skolen I offra en bock såsom syndoffer -- detta förutom det dagliga brännoffret med tillhörande spisoffer och drickoffer.
Och på den andra dagen: tolv ungtjurar, två vädurar, fjorton årsgamla felfria lamm,
med det spisoffer och de drickoffer som skola offras till dem, till tjurarna, vädurarna och lammen, efter deras antal, på föreskrivet sätt,
tillika också en bock såsom syndoffer -- detta förutom det dagliga brännoffret med tillhörande spisoffer och det drickoffer som hör till dem.
Och på den tredje dagen: elva tjurar, två vädurar, fjorton årsgamla felfria lamm,
med det spisoffer och de drickoffer som skola offras till dem, till tjurarna, vädurarna och lammen, efter deras antal, på föreskrivet sätt,
tillika också en syndoffersbock -- detta förutom det dagliga brännoffret med tillhörande spisoffer och drickoffer.
Och på den fjärde dagen; tio tjurar, två vädurar, fjorton årsgamla felfria lamm,
med det spisoffer och de drickoffer som skola offras till dem, till tjurarna, vädurarna och lammen, efter deras antal, på föreskrivet satt,
tillika också en bock såsom syndoffer -- detta förutom det dagliga brännoffret med tillhörande spisoffer och drickoffer.
Och på den femte dagen: nio tjurar, två vädurar, fjorton årsgamla felfria lamm,
med det spisoffer och de drickoffer som skola offras till dem, till tjurarna, vädurarna och lammen, efter deras antal, på föreskrivet sätt,
tillika också en syndoffersbock -- detta förutom det dagliga brännoffret med tillhörande spisoffer och drickoffer.
Och på den sjätte dagen: åtta tjurar, två vädurar, fjorton årsgamla felfria lamm,
med det spisoffer och de drickoffer som skola offras till dem, till tjurarna, vädurarna och lammen, efter deras antal, på föreskrivet sätt,
tillika också en syndoffersbock -- detta förutom det dagliga brännoffret med tillhörande spisoffer och drickoffer.
Och på den sjunde dagen: sju tjurar, två vädurar, fjorton årsgamla felfria lamm,
med det spisoffer och de drickoffer som skola offras till dem, till tjurarna, vädurarna och lammen, efter deras antal, på föreskrivet sätt,
tillika också en syndoffersbock -- detta förutom det dagliga brännoffret med tillhörande spisoffer och drickoffer.
På den åttonde dagen skolen I hålla en högtidsförsamling; ingen arbetssyssla skolen I då göra.
Och såsom brännoffer, såsom eldsoffer, skolen I då offra till en välbehaglig lukt för HERREN en tjur, en vädur, sju årsgamla felfria lamm,
med det spisoffer och de drickoffer som skola offras till dem, till tjuren, väduren och lammen, efter deras antal, på föreskrivet sätt,
tillika också en syndoffersbock -- detta förutom det dagliga brännoffret med tillhörande spisoffer och drickoffer.
Dessa offer skolen I offra åt HERREN vid edra högtider, förutom edra löftesoffer och frivilliga offer, dessa må nu vara brännoffer eller spisoffer eller drickoffer eller tackoffer.
Och Mose sade detta till Israels barn, alldeles såsom HERREN hade bjudit honom.
Och Mose talade till Israels barns stamhövdingar och sade: Detta är vad HERREN har bjudit:
om någon gör ett löfte åt HERREN, eller svär en ed genom vilken han förbinder sig till återhållsamhet i något stycke, så skall han icke sedan bryta sitt ord; han skall i alla stycken göra vad hans mun har talat.
Och om en kvinna, medan hon vistas i sin faders hus och ännu är ung, gör ett löfte åt HERREN och förbinder sig till återhållsamhet i något stycke,
och hennes fader hör hennes löfte och huru hon förbinder sig till återhållsamhet, och hennes fader icke säger något till henne därom, så skola alla hennes löften hava gällande kraft, och alla hennes förbindelser till återhållsamhet skola hava gällande kraft.
Men om hennes fader samma dag han hör det säger nej därtill, då skola hennes löften och hennes förbindelser till återhållsamhet alla vara utan gällande kraft; och HERREN skall förlåta henne, eftersom hennes fader sade nej till henne.
Och om hon bliver gift, och löften då vila på henne, eller något obetänksamt ord från hennes läppar, varmed hon har bundit sig,
och hennes man får höra därom, men icke säger något till henne därom samma dag han hör det, så skola hennes löften hava gällande kraft, och hennes förbindelser till återhållsamhet skola hava gällande kraft.
Men om hennes man samma dag han får höra det säger nej därtill, då upphäver han därmed hennes givna löfte och det obetänksamma ord från hennes läppar, varmed hon har bundit sig; och HERREN skall förlåta henne det.
Men en änkas eller en förskjuten hustrus löfte skall hava gällande kraft för henne, vartill hon än må hava förbundit sig.
Och om en kvinna i sin mans hus gör ett löfte, eller med ed förbinder sig till återhållsamhet i något stycke,
och hennes man hör det, men icke säger något till henne därom -- icke säger nej till henne -- så skola alla hennes löften hava gällande kraft, och alla hennes förbindelser till återhållsamhet skola hava gällande kraft.
Men om hennes man upphäver dem samma dag han hör dem, då skall allt som hennes läppar hava talat vara utan gällande kraft, det må nu vara löften eller någon förbindelse till återhållsamhet; hennes man har upphävt dem, därför skall HERREN förlåta henne.
Åt alla hennes löften och åt alla hennes edliga förbindelser till att späka sig kan hennes man giva gällande kraft, och hennes man kan ock upphäva dem.
Men om hennes man icke före påföljande dags ingång säger någonting till henne därom, så giver han gällande kraft åt alla hennes löften och åt alla de förbindelser till återhållsamhet, som vila på henne; han giver dem gällande kraft därigenom att han icke säger något till henne därom samma dag han hör dem.
Men om han upphäver dem först någon tid efter det han har hört dem, då kommer han att bära på hennes missgärning.
Dessa äro de stadgar som HERREN av Mose angående förhållandet mellan en man och hans hustru, och angående förhållandet mellan en fader och hans dotter, medan denna ännu är ung och vistas i sin faders hus.
Och HERREN talade till Mose och sade:
»Kräv ut hämnd för Israels barn midjaniterna; sedan skall du samlas till dina fäder.
Då talade Mose till folket och sade: »Låten en del av edra män väpna sig till strid; dessa skola tåga mot Midjan och utföra HERRENS hämnd på Midjan.
Tusen man ur var och en särskild av Israels alla stammar skolen I sända ut i striden.»
Så avlämnades då ur Israels ätter tusen man av var stam: tolv tusen man, väpnade till strid.
Och Mose sände dessa, tusen man av var stam, ut i striden; han sände med dem Pinehas, prästen Eleasars son, ut i striden, och denne tog med sig de heliga redskapen och larmtrumpeterna.
Och de gingo till strids emot Midjan, såsom HERREN hade bjudit Mose, och dräpte allt mankön.
Och jämte andra som då blevo slagna av dem dräptes ock de midjanitiska konungarna Evi, Rekem, Sur, Hur och Reba, fem midjanitiska konungar; Bileam, Beors son, dräpte de ock med svärd.
Och Israels barn förde Midjans kvinnor och barn bort såsom fångar; och alla deras dragare och all deras boskap och allt deras övriga gods togo de såsom byte.
Och alla deras städer, i de trakter där de bodde, och alla deras tältläger brände de upp i eld.
Och de togo med sig allt bytet, och allt vad de hade rövat, både människor och boskap.
Och de förde fångarna och det rövade och bytet fram till Mose och prästen Eleasar och Israels barns menighet i lägret på Moabs hedar, som ligga vid Jordan mitt emot Jeriko.
Och Mose och prästen Eleasar och alla menighetens hövdingar gingo dem till mötes utanför lägret.
Men Mose förtörnades på krigsbefälet, över- och underhövitsmännen, när de kommo tillbaka från sitt krigståg.
Mose sade till dem: »Haven I då låtit alla kvinnorna leva?
Det var ju de som, på Bileams inrådan, förledde Israels barn till att begå otrohet mot HERREN i saken med Peor, och som därigenom vållade att en hemsökelse kom över HERRENS menighet.
Så dräpen nu alla gossebarn, och dräpen alla kvinnor som hava haft med män, med mankön, att skaffa.
Men alla flickebarn som icke hava haft med mankön att skaffa, dem mån I låta leva för eder räkning.
Själva skolen I nu lägra eder utanför lägret, i sju dagar.
Var och en av eder som har dräpt någon människa, och var och en som har kommit vid någon slagen skall rena sig på tredje dagen och på sjunde dagen -- såväl I själva som edra fångar.
Alla kläder och allt som är förfärdigat av skinn och allt som är gjort av gethår och alla redskap av trä skolen I ock rena åt eder.»
Och prästen Eleasar sade till stridsmännen som hade deltagit i kriget: Detta är den lagstadga som HERREN har givit Mose:
Guld och silver, koppar, järn, tenn och bly,
allt sådant som tål eld, skolen I låta gå genom eld, så bliver det rent; dock bör det tillika renas med stänkelsevatten.
Men allt som icke tål eld skolen I låta gå genom vatten.
Och I skolen två edra kläder på sjunde dagen, så bliven I rena; därefter fån I gå in i lägret.
Och HERREN talade till Mose och sade:
Över det tagna rovet, både människor och boskap, skall du göra en beräkning, du tillsammans med prästen Eleasar och huvudmännen för menighetens familjer;
sedan skall du dela rovet i två delar, mellan de krigare som hava varit med i striden och hela den övriga menigheten.
Och du skall låta det krigsfolk som har varit med i striden giva var femhundrade av människor, fäkreatur, åsnor och får såsom skatt åt HERREN.
Så mycket skall tagas av den hälft som tillfaller dem, och du skall giva detta åt prästen Eleasar såsom en gärd åt HERREN.
Men ur den hälft som tillfaller de övriga israeliterna skall du uttaga var femtionde av människor, sammalunda av fäkreatur, åsnor och får, korteligen, av all boskap, och detta skall du giva åt leviterna, som det åligger att iakttaga vad som är att iakttaga vid HERRENS tabernakel.
Och Mose och prästen Eleasar gjorde såsom HERREN hade bjudit Mose.
Och rovet, nämligen återstoden av det byte som krigsfolket hade tagit utgjorde: av får sex hundra sjuttiofem tusen,
av fäkreatur sjuttiotvå tusen,
av åsnor sextioett tusen,
och av människor, sådana kvinnor som icke hade haft med mankön att skaffa, tillsammans trettiotvå tusen personer.
Och hälften därav, eller den del om tillföll dem som hade varit med striden, utgjorde: av får ett antal av tre hundra trettiosju tusen fem hundra,
varav skatten åt HERREN utgjorde sex hundra sjuttiofem får;
av fäkreatur trettiosex tusen, varav skatten åt HERREN sjuttiotvå;
av åsnor trettio tusen fem hundra, varav skatten åt HERREN sextioen;
av människor sexton tusen, varav skatten åt HERREN trettiotvå personer.
Och skatten, den för HERREN bestämda gärden, gav Mose åt prästen Eleasar, såsom HERREN hade bjudit Mose.
Och den hälft, som tillföll de övriga israeliterna, och som Mose hade avskilt från krigsfolkets,
denna hälft, den som tillföll menigheten, utgjorde: av får tre hundra trettiosju tusen fem hundra,
av fäkreatur trettiosex tusen,
av åsnor trettio tusen fem hundra
och av människor sexton tusen.
Och ur denna hälft, som tillföll de övriga israeliterna, uttog Mose var femtionde, både av människor och av boskap, och gav detta åt leviterna, som det ålåg att iakttaga vad som var att iakttaga vid HERRENS tabernakel, allt såsom HERREN hade bjudit Mose.
Och befälhavarna över härens avdelningar, över- och underhövitsmännen, trädde fram till Mose.
Och de sade till Mose: »Dina tjänare hava räknat antalet av de krigsmän som vi hava haft under vårt befäl, och icke en enda fattas bland oss.
Därför hava vi nu såsom en offergåva åt HERREN burit fram var och en del som han har kommit över av gyllene klenoder, armband av olika slag, ringar, örhängen och halssmycken, detta för att bringa försoning för oss inför HERRENS ansikte.»
Och Mose och prästen Eleasar togo emot guldet av dem, alla slags klenoder.
Och guldet som gavs såsom gärd åt HERREN av över- och underhövitsmännen utgjorde sammanlagt sexton tusen sju hundra femtio siklar.
Manskapet hade tagit byte var och en för sig.
Och Mose och prästen Eleasar togo emot guldet av över- och underhövitsmännen och buro in det i uppenbarelsetältet, för att det skulle bringa Israels barn i åminnelse inför HERRENS ansikte.
Och Rubens barn och Gads barn hade stora och mycket talrika boskapshjordar; och när de sågo Jaesers land och Gileads land, funno de att detta var en trakt för boskap.
Då kommo Gads barn och Rubens barn och sade till Mose och prästen Eleasar och menighetens hövdingar:
»Atarot, Dibon, Jaeser, Nimra, Hesbon, Eleale, Sebam, Nebo och Beon,
det land som HERREN har låtit Israels menighet intaga, är ett land för boskap, och dina tjänare hava boskap.»
Och de sade ytterligare: »Om vi hava funnit nåd inför dina ögon så må detta land givas åt dina tjänare till besittning.
Låt oss slippa att gå över Jordan.»
Men Mose sade till Gads barn och Rubens barn: »Skolen då I stanna här, under det att edra bröder draga ut i krig?
Varför viljen I avvända Israels barns hjärtan från att gå över floden, in i det land som HERREN har givit åt dem?
Så gjorde ock edra fäder, när jag sände dem från Kades-Barnea för att bese landet:
sedan de hade dragit upp till Druvdalen och besett landet, avvände de Israels barns hjärtan från att gå in i det land som HERREN hade givit åt dem.
Och på den dagen upptändes HERRENS vrede, och han svor och sade:
'Av de män som hava dragit upp ur Egypten skall ingen som är tjugu år gammal eller därutöver få se det land som jag med ed har lovat åt Abraham, Isak och Jakob -- eftersom de icke i allt hava efterföljt mig
ingen förutom Kaleb, Jefunnes son, kenaséen, och Josua, Nuns son; ty de hava i allt efterföljt HERREN.'
Så upptändes HERRENS vrede mot Israel, och han lät dem driva omkring i öknen i fyrtio år, till dess att hela det släkte hade dött bort som hade gjort vad ont var i HERRENS ögon.
Och se, nu haven I trätt i edra fäders fotspår, I, syndiga mäns avföda, och öken så ännu mer HERRENS vredes glöd mot Israel.
Då I nu vänden eder bort ifrån honom, skall han låta Israel ännu längre bliva kvar i öknen, och I dragen så fördärv över allt detta folk.»
Då trädde de fram till honom och sade: »Låt oss här bygga gårdar åt var boskap och städer åt våra kvinnor och barn.
Själva vilja vi sedan skyndsamt väpna oss och gå åstad i spetsen för Israels barn, till dess vi hava fört dem dit de skola.
Under tiden kunna våra kvinnor och barn bo i de befästa städerna och så vara skyddade mot landets inbyggare.
Vi skola icke vända tillbaka hem, förrän Israels barn hava fått var och en sin arvedel.
Ty vi vilja icke taga vår arvedel jämte dem, på andra sidan Jordan och längre bort, utan vår arvedel har tillfallit oss här på andra sidan Jordan, på östra sidan.»
Mose svarade dem: »Om I gören såsom I nu haven sagt, om I väpnen eder inför HERREN till kriget,
så att alla edra väpnade män gå över Jordan inför HERREN och stanna där, till dess han har fördrivit sina fiender för sig,
om I alltså vänden tillbaka först då landet har blivit HERREN underdånigt, så skolen I vara utan skuld mot HERREN och Israel, och detta land skall då bliva eder besittning inför HERREN.
Men om I icke så gören, se, då synden I mot HERREN, och I skolen då komma att förnimma eder synd, ty den skall drabba eder.
Byggen eder nu städer åt edra kvinnor och barn, och gårdar åt eder boskap, och gören vad eder mun har talat.»
Och Gads barn och Rubens barn talade till Mose och sade: »Dina tjänare skola göra såsom min herre bjuder.
Våra barn våra hustrur, vår boskap och alla våra dragare skola bliva kvar här i Gileads städer.
Men dina tjänare, vi så många som äro väpnade till strid, skola draga ditöver och kämpa inför HERREN, såsom min herre har sagt.»
Och Mose gav befallning om dem åt prästen Eleasar och åt Josua, Nuns son, och åt huvudmännen för familjerna inom Israels barns stammar.
Mose sade till dem: »Om Gads barn och Rubens barn gå över Jordan med eder, så många som äro väpnade till att kämpa inför HERREN, och landet så bliver eder underdånigt, då skolen I åt dem giva landet Gilead till besittning.
Men om de icke draga väpnade ditöver med eder, så skola de få sin besittning ibland eder i Kanaans land.»
Och Gads barn och Rubens barn svarade och sade: »Vad HERREN har sagt till dina tjänare, det vilja vi göra.
Vi vilja draga väpnade över till Kanaans land inför HERREN, och så få vår arvsbesittning har på andra sidan Jordan.»
Så gav då Mose åt dem, åt Gads barn, Rubens barn och ena hälften av Manasses, Josefs sons, stam, Sihons, amoréernas konungs, rike och Ogs rike, konungens i Basan: själva landet med dess städer och dessas områden, landets städer runt omkring.
Och Gads barn byggde upp Dibon, Atarot, Aroer,
Atrot-Sofan, Jaeser, Jogbeha,
Bet-Nimra och Bet-Haran, befästa städer och boskapsgårdar.
Och Rubens barn byggde upp Hesbon, Eleale, Kirjataim,
Nebo och Baal-Meon -- vilkas namn hava ändrats -- och Sibma.
Och de gåvo namn åt städerna som de byggde upp.
Och Makirs, Manasses sons, barn gingo åstad till Gilead och intogo det och fördrevo amoréerna som bodde där.
Och Mose gav Gilead åt Makir, Manasses son, och han bosatte sig där.
Och Jair, Manasses son, gick åstad och intog deras byar och kallade dem Jairs byar.
Och Noba gick åstad och intog Kenat, med underlydande orter, och kallade det Noba, efter sitt eget namn.
Dessa voro Israels barns lägerplatser, när de drogo ut ur Egyptens land, efter sina härskaror, anförda av Mose och Aron.
Och Mose upptecknade på HERRENS befallning deras uppbrottsorter, alltefter som de ändrade lägerplats.
Och dessa voro nu deras lägerplatser, alltefter som uppbrottsorterna följde på varandra:
De bröto upp från Rameses i första månaden, på femtonde dagen i första månaden.
Dagen efter påskhögtiden drogo Israels barn ut med upplyft hand inför alla egyptiers ögon,
under det att egyptierna begrovo dem som HERREN hade slagit bland dem, alla de förstfödda, då när HERREN höll dom över deras gudar.
Så bröto nu Israels barn upp från Rameses och lägrade sig i Suckot.
Och de bröto upp från Suckot och lägrade sig i Etam, där öknen begynte.
Och de bröto upp från Etam och vände om till Pi-Hahirot, som ligger mitt emot Baal-Sefon, och lägrade sig framför Migdol.
Och de bröto upp från Hahirot och gingo mitt igenom havet in i öknen och tågade så tre dagsresor i Etams öken och lägrade sig i Mara.
Och de bröto upp från Mara och kommo till Elim; och i Elim funnos tolv vattenkällor och sjuttio palmträd, och de lägrade sig där.
Och de bröto upp från Elim och lägrade sig vid Röda havet.
Och de bröto upp från Röda havet och lägrade sig i öknen Sin.
Och de bröto upp från öknen Sin och lägrade sig i Dofka.
Och de bröto upp från Dofka och lägrade sig i Alus.
Och de bröto upp från Alus och lägrade sig i Refidim, och där fanns intet vatten åt folket att dricka.
Och de bröto upp från Refidim och lägrade sig i Sinais öken.
Och de bröto upp från Sinais öken och lägrade sig i Kibrot-Hattaava.
Och de bröto upp från Kibrot-Hattaava och lägrade sig i Haserot.
Och de bröto upp från Haserot och lägrade sig i Ritma.
Och de bröto upp från Ritma och lägrade sig i Rimmon-Peres.
Och de bröto upp från Rimmon-Peres och lägrade sig i Libna.
Och de bröto upp från Libna och lägrade sig i Rissa.
Och de bröto upp från Rissa och lägrade sig i Kehelata.
Och de bröto upp från Kehelata och lägrade sig vid berget Sefer.
Och de bröto upp från berget Sefer och lägrade sig i Harada.
Och de bröto upp från Harada och lägrade sig i Makhelot.
Och de bröto upp från Makhelot och lägrade sig i Tahat.
Och de bröto upp från Tahat och lägrade sig i Tera.
Och de bröto upp från Tera och lägrade sig i Mitka.
Och de bröto upp från Mitka och lägrade sig i Hasmona.
Och de bröto upp från Hasmona och lägrade sig i Moserot.
Och de bröto upp från Moserot och lägrade sig i Bene-Jaakan.
Och de bröto upp från Bene-Jaakan och lägrade sig i Hor-Haggidgad.
Och de bröto upp från Hor-Haggidgad och lägrade sig i Jotbata.
Och de bröto upp från Jotbata och lägrade sig i Abrona.
och de bröto upp från Abrona och lägrade sig i Esjon-Geber.
Och de bröto upp från Esjon-Geber och lägrade sig i öknen Sin, det är Kades.
Och de bröto upp från Kades och lägrade sig vid berget Hor, på gränsen till Edoms land.
Och prästen Aron steg upp på berget Hor, efter HERRENS befallning, och dog där i det fyrtionde året efter Israels barns uttåg ur Egyptens land, i femte månaden, på första dagen i månaden.
Och Aron var ett hundra tjugutre år gammal, när han dog på berget Hor.
Och konungen i Arad, kananéen, som bodde i Sydlandet i Kanaans land, fick nu höra att Israels barn voro i antågande.
Och de bröto upp från berget Hor och lägrade sig i Salmona.
Och de bröto upp från Salmona och lägrade sig i Punon.
Och de bröto upp från Punon och lägrade sig i Obot.
Och de bröto upp från Obot och lägrade sig i Ije-Haabarim vid Moabs gräns.
Och de bröto upp från Ijim och lägrade sig i Dibon-Gad.
Och de bröto upp från Dibon-Gad och lägrade sig i Almon-Diblataima.
Och de bröto upp från Almon-Diblataima och lägrade sig vid Abarimbergen, framför Nebo.
Och de bröto upp från Abarimbergen och lägrade sig på Moabs hedar, vid Jordan mitt emot Jeriko.
Och deras läger vid Jordan sträckte sig från Bet-Hajesimot ända till Abel-Hassitim på Moabs hedar.
Och HERREN talade till Mose på Moabs hedar, vid Jordan mitt emot Jeriko, och sade:
Tala till Israels barn och säg till dem: När I haven gått över Jordan, in i Kanaans land,
skolen I fördriva landets alla inbyggare för eder, och I skolen förstöra alla deras stenar med inhuggna bilder, och alla deras gjutna beläten skolen I förstöra, och alla deras offerhöjder skolen I ödelägga.
Och I skolen intaga landet och bosätta eder där, ty åt eder har jag givit landet till besittning.
Och I skolen utskifta landet såsom arvedel åt eder genom lottkastning efter edra släkter; åt en större stam skolen I giva en större arvedel, och åt en mindre stam en mindre arvedel; var och en skall få sin del där lotten bestämmer att han skall hava den; efter edra fädernestammar skolen I utskifta landet såsom arvedel åt eder.
Men om I icke fördriven landets inbyggare för eder, så skola de som I låten vara kvar av dem bliva törnen i edra ögon och taggar i edra sidor, och skola tränga eder i landet där I bon.
Och då skall jag göra med eder så, som jag hade tänkt göra med dem.
Och HERREN talade till Mose och sade:
Bjud Israels barn och säg till dem: När I kommen till Kanaans land, då är detta det land som skall tillfalla eder såsom arvedel: Kanaans land, så långt dess gränser nå.
Edert land skall på södra sidan sträcka sig från öknen Sin utmed Edom; och eder södra gräns skall i öster begynna vid ändan av Salthavet.
Sedan skall eder gräns böja sig söder om Skorpionhöjden och gå fram till Sin och gå ut söder om Kades-Barnea.
Och den skall gå vidare ut till Hasar-Addar och fram till Asmon.
Och från Asmon skall gränsen böja sig mot Egyptens bäck och gå ut vid havet.
Och eder gräns i väster skall vara Stora havet; det skall utgöra gränsen.
Detta skall vara eder gräns i väster.
Och detta skall vara eder gräns i norr: Från Stora havet skolen I draga eder gränslinje fram vid berget Hor.
Från berget Hor skolen I draga eder gränslinje dit där vägen går till Hamat, och gränsen skall gå ut vid Sedad.
Sedan skall gränsen gå till Sifron och därifrån ut vid Hasar-Enan.
Detta skall vara eder gräns i norr.
och såsom eder gräns i öster skolen I draga upp en linje från Hasar-Enan fram till Sefam.
Och från Sefam skall gränsen gå ned till Haribla, öster om Ain, och gränsen skall gå vidare ned och intill bergsluttningen vid Kinneretsjön, österut.
Sedan skall gränsen gå ned till Jordan och ut vid Salthavet.
Detta skall vara edert land, med dess gränser runt omkring.
Och Mose bjöd Israels barn och sade: Detta är det land som I genom lottkastning skolen utskifta såsom arvedel åt eder, det land om vilket HERREN har bjudit att det skall givas åt de nio stammarna och den ena halva stammen.
Ty rubeniternas barns stam, efter dess familjer, och gaditernas barns stam, efter dess familjer, och den andra hälften av Manasse stam, dessa hava redan fått sin arvedel.
Dessa två stammar och denna halva stam hava fått sin arvedel på andra sidan Jordan mitt emot Jeriko, österut mot solens uppgång.
Och HERREN talade till Mose och sade:
Dessa äro namnen på de män som skola åt eder utskifta landet i arvslotter: först och främst prästen Eleasar och Josua, Nuns son;
vidare skolen I taga en hövding ur var stam till att utskifta landet,
och dessa äro de männens namn: av Juda stam Kaleb, Jefunnes son;
av Simeons barns stam Samuel Ammihuds son;
av Benjamins stam Elidad, Kislons son;
av Dans barns stam en hövding, Bucki, Joglis son;
av Josefs barn: av Manasse barns stam en hövding, Hanniel, Efods son,
och av Efraims barn stam en hövding, Kemuel, Siftans son;
av Sebulons barns stam en hövding, Elisafan, Parnaks son;
av Isaskars barns stam en hövding, Paltiel, Assans son;
av Asers barns stam en hövding, Ahihud, Selomis son;
av Naftali barns stam en hövding, Pedael, Ammihuds son.
Dessa äro de som HERREN bjöd att utskifta arvslotterna åt Israels barn i Kanaans land.
Och HERREN talade till Mose på Moabs hedar, vid Jordan mitt emot Jeriko, och sade:
Bjud Israels barn att de av de arvslotter de få till besittning skola åt leviterna giva städer att bo i; utmarker runt omkring dessa städer skolen I ock giva åt leviterna.
Städerna skola de själva hava att bo i, men de tillhörande utmarkerna skola vara för deras dragare och deras boskap och alla deras övriga djur.
Och städernas utmarker, som I skolen giva åt leviterna, skola sträcka sig tusen alnar från stadsmuren utåt på alla sidor.
Och utanför staden skolen I mäta upp på östra sidan två tusen alnar, på västra sidan två tusen alnar, på södra sidan två tusen alnar och på norra sidan två tusen alnar, med staden i mitten.
Detta skola de få såsom utmarker till sina städer.
Och de städer som I given åt leviterna skola först och främst vara de sex fristäderna, vilka I skolen giva till det ändamålet att en dråpare må kunna fly till dem; vidare skolen I jämte dessa städer giva dem fyrtiotvå andra,
så att de städer som I given åt leviterna tillsammans utgöra fyrtioåtta städer, med tillhörande utmarker.
Och av dessa städer, som I skolen giva av Israels barns besittningsområde, skolen I taga flera ur den stam som är större, och färre ur den som är mindre.
Var stam skall åt leviterna giva ett antal av sina städer, som svarar mot den arvedel han själv har fått.
Och HERREN talade till Mose och sade:
Tala till Israels barn och säg till dem: När I haven gått över Jordan, in i Kanaans land,
skolen I utse åt eder vissa städer, som I skolen hava till fristäder, till vilka en dråpare som ouppsåtligen har dödat någon må kunna fly.
Och dessa städer skolen I hava såsom tillflyktsorter undan blodshämnaren, så att dråparen slipper dö, förrän han har stått till rätta inför menigheten.
Och de städer som I skolen giva till fristäder skola vara sex.
Tre av städerna skolen I giva på andra sidan Jordan, och de tre övriga städerna skolen I giva i själva Kanaans land;
dessa skola vara fristäder.
Israels barn, såväl som främlingen och inhysesmannen som bor ibland dem skola hava dessa sex städer såsom tillflyktsorter, till vilka var och er som ouppsåtligen har dödat någon må kunna fly.
Men om någon slår en annan till döds med ett föremål av järn, så är han en sannskyldig dråpare; en sådan skall straffas med döden.
Likaledes, om någon i sin hand har en sten med vilken ett dråpslag kan givas, och han därmed slår en annan till döds, så är han en sannskyldig dråpare; en sådan skall straffas med döden.
Eller om någon i sin hand har ett föremål av trä varmed ett dråpslag kan givas, och han därmed slår en annan till döds, så är han en sannskyldig dråpare; en sådan skall straffas med döden.
Blodshämnaren må döda den dråparen; varhelst han träffar på honom må han döda honom.
Likaledes om någon av hat stöter till en annan, eller med berått mod kastar något på honom; så att han dör,
eller av fiendskap slår honom till döds med handen, då skall den som gav slaget straffas med döden, ty han är en sannskyldig dråpare; blodshämnaren må döda den dråparen, varhelst han träffar på honom
Men om någon av våda, utan fiendskap, stöter till en annan, eller utan berått mod kastar på honom något föremål, vad det vara må;
eller om han, utan att se honom, med någon sten varmed dråpslag kan givas träffar honom, så att han dör, och detta utan att han var hans fiende eller hade för avsikt att skada honom,
då skall menigheten döma mellan den som gav slaget och blodshämnaren, enligt här givna föreskrifter.
Och menigheten skall rädda dråparen ur blodshämnarens hand, och menigheten skall låta honom vända tillbaka till fristaden dit han hade flytt, och där skall han stanna kvar, till dess den med helig olja smorde översteprästen dör.
Men om dråparen går utom området för den fristad dit han har flytt,
och blodshämnaren då, när han träffar på honom utom hans fristads område, dräper dråparen, så vilar ingen blodskuld på honom.
Ty i sin fristad skall en dråpare stanna kvar, till dess översteprästen dör; men efter översteprästens död må han vända tillbaka till den ort där han har sin besittning.
Och detta skall vara en rättsstadga för eder från släkte till släkte, var I än ären bosatta.
Om någon slår ihjäl en annan, skall man, efter vittnens utsago, dräpa dråparen; men en enda persons vittnesmål är icke nog för att man skall kunna döma någon till döden.
I skolen icke taga lösen för en dråpares liv, om han är skyldig till döden, utan han skall straffas med döden.
Ej heller skolen I taga lösen för att den som har flytt till en fristad skall före prästens död få vända tillbaka och bo i landet.
I skolen icke ohelga det land där I ären; genom blod ohelgas landet, och försoning kan icke bringas för landet för det blod som har blivit utgjutet däri, annat än genom dens blod, som har utgjutit det.
I skolen icke orena landet där I bon, det i vars mitt jag har min boning, ty jag, HERREN, har min boning mitt ibland Israels barn.
Och huvudmännen för familjerna i Gileads barns släkt -- Gileads, som var son till Makir, Manasses son, av Josefs barns släkter -- trädde fram och talade inför Mose och de hövdingar som voro huvudmän för Israels barns familjer.
De sade: »HERREN har bjudit min herre att genom lottkastning göra landet såsom arvedel åt Israels barn och HERREN har vidare bjudit min herre att giva Selofhads, vår broders, arvedel åt hans döttrar.
Men om nu dessa bliva gifta med någon ur Israels barns andra stammar, så tages deras arvedel bort ifrån våra fäders arvedel, under det att den stam de komma att tillhöra får sin arvedel ökad; på detta sätt bliver en del av vår arvslott oss fråntagen.
När sedan jubelåret inträder för Israels barn, bliver deras arvedel lagd till den stams arvedel, som de komma att tillhöra, men från vår fädernestams arvedel tages deras arvedel bort.»
Då bjöd Mose Israels barn, efter HERRENS befallning, och sade: »Josefs barns stam har talat rätt.
Detta är vad HERREN bjuder angående Selofhads döttrar; han säger: De må gifta sig med vem de finna för gott, allenast de gifta sig inom en släkt som hör till deras egen fädernestam.
Ty en arvedel som tillhör någon, av Israels barn må icke gå över från en stam till en annan, utan Israels barn skola behålla kvar var och en sin fädernestams arvedel.
Och när en kvinna som inom någon av Israels barns stammar har kommit i besittning av en arvedel gifter sig, skall det vara med en man av någon släkt som hör till hennes egen fädernestam, så att Israels barn förbliva i besittning var och en av sina fäders arvedel.
Ty ingen arvedel må gå över från en stam till en annan, utan Israels barns stammar skola behålla kvar var och en sin arvedel.»
Selofhads döttrar gjorde såsom HERREN hade bjudit Mose.
Mahela, Tirsa, Hogla, Milka och Noa, Selofhads döttrar, gifte sig med sina farbröders söner.
De blevo alltså gifta inom Manasses, Josefs sons, barns släkter, och deras arvedel stannade så kvar inom deras fädernesläkts stam.
Dessa äro de bud och rätter som HERREN genom Mose gav Israels barn, på Moabs hedar, vid Jordan mitt emot Jeriko.
Dessa äro de ord som Mose talade till hela Israel på andra sidan Jordan, i öknen, på Hedmarken mitt emot Suf, mellan Paran och Tofel, Laban, Haserot och Di-Sahab
-- elva dagsresor från Horeb, åt Seirs bergsbygd till, fram till Kades-Barnea.
I det fyrtionde året, i elfte månaden. på första dagen i månaden, talade Mose till Israels barn, alldeles såsom Herren hade bjudit honom tala till dem.
Detta skedde sedan han hade slagit Sihon, amoréernas konung, som bodde i Hesbon, och Og, konungen i Basan, som bodde i Astarot, vid Edrei.
På andra sidan Jordan. i Moabs land, begynte Mose denna lagutläggning och sade:
HERREN, vår Gud, talade till oss på Horeb och sade: »Länge nog haven I uppehållit eder vid detta berg.
Vänden eder nu åt annat håll och bryten upp, och begiven eder till amoréernas bergsbygd och till alla deras grannfolk på Hedmarken, i Bergsbygden, i Låglandet, i Sydlandet och i Kustlandet vid havet -- in i kananéernas land och upp på Libanon, ända till den stora floden, floden Frat.
Se, jag har givit landet i edert våld.
Gån nu och intagen detta land, som HERREN med ed har lovat edra fäder, Abraham, Isak och Jakob, att giva åt dem och åt deras säd efter dem.»
Och jag talade till eder på den tiden och sade: »Jag förmår icke ensam bära eder.
HERREN, eder Gud, har förökat eder, och se, I ären nu talrika såsom stjärnorna på himmelen.
Må Herren, edra fäders Gud, än vidare föröka eder tusenfalt och välsigna eder, såsom han har lovat eder.
Men huru skall jag ensam kunna bära tyngden och bördan av eder och edert tvistande?
Utsen åt eder visa, förståndiga och välkända män inom edra särskilda stammar, så skall jag sätta dem till huvudmän över eder.»
I svaraden mig och saden: »Ditt förslag är gott.»
Då tog jag huvudmännen i edra stammar, visa och välkända män, och satte dem till huvudmän över eder, till föreståndare, somliga över tusen, andra över hundra, andra över femtio och somliga över tio, och till tillsyningsmän i edra särskilda stammar.
Och jag bjöd då också edra domare och sade: »Hören efter, vad edra bröder hava sig emellan; och om någon har en sak med sin broder eller med en främling som bor hos honom, så dömen rättvist mellan dem.
I skolen icke hava anseende till personen, när I dömen, utan höra den ringe likaväl dom den högre; I skolen icke frukta för någon människa, ty domen hör Gud till.
Men om något ärende bliven eder för svårt, skolen I hänskjuta det till mig, så att jag för höra det.»
Så bjöd jag eder på den tiden allt vad I skullen göra.
Och vi bröto upp från Horeb, och genom hela den stora och fruktansvärda öken som I haven sett vandrande vi åstad till amoréernas bergsbygd, såsom HERREN, vår Gud, hade bjudit oss; och vi kommo så till Kades-Barnea.
Och jag sade till eder: »I haven nu kommit till amoréernas bergsbygd, som HERREN vår Gud, vill giva oss.
Se, HERREN, din Gud, har givit landet i ditt våld.
Drag ditupp och intag det, såsom HERREN, dina fäders Gud, har tillsagt dig.
Frukta icke och var icke förfärad.»
Då trädden I fram till mig allasammans och saden: »Låt oss sända åstad några män framför oss, för att de må utforska landet åt oss och sedan avgiva sin berättelse inför oss, angående vägen på vilken vi skola draga ditupp, och angående de städer som vi skola komma till.»
Detta förslag behagade mig, och jag tog tolv män bland eder, en för var stam.
Dessa begåvo sig åstad och drogo upp till Bergsbygden och kommo till Druvdalen och bespejade landet.
Och de togo med sig av landets frukt ned till oss och avgåvo sin berättelse inför oss och sade: »Det land som Herren, vår Gud, vill giva oss är gott.»
Men I villen icke draga ditupp, utan voren gensträviga mot HERRENS, eder Guds, befallning.
Och I knorraden i edra tält och saden: »Herren hatar oss, därför har han fört oss ut ur Egyptens land för att giva oss i amoréernas hand och så förgöra oss.
Varthän skola vi då draga?
Våra bröder hava förfärat våra hjärtan, ty de säga: 'Där är ett folk, större och resligare än vi, där äro städer, stora och befästa upp mot himmelen; ja, vi sågo där också anakiter.'»
Då svarade jag eder: »I skolen icke förskräckas och icke frukta för dem.
HERREN, eder Gud, som går framför eder, skall själv strida för eder, alldeles såsom han handlade mot eder i Egypten inför edra ögon,
och alldeles såsom i öknen som du har sett, där HERREN, din Gud, bar dig, såsom en man bär sin son, hela den väg I haven vandrat, ända till dess att I nu haven kommit hit.»
Men detta oaktat trodden I icke på HERREN, eder Gud,
som gick framför eder på vägen, för att utse lägerplatser åt eder: om natten i eld, för att lysa eder på den väg I skullen gå, och om dagen i molnskyn.
Då nu HERREN hörde edra ord, blev han förtörnad och svor och sade:
»Sannerligen, ingen av dessa män, i detta onda släkte, skall få se det goda land som jag med ed har lovat giva åt edra fäder,
ingen utom Kaleb, Jefunnes son; han skall få se det, och åt honom och åt hans barn skall jag giva det land han har beträtt, därför att han i allt har efterföljt Herren.»
Också på mig vredgades HERREN, för eder skull, och sade: »Icke heller du skall komma ditin.
Josua, Nuns son, han som är din tjänare, han skall komma ditin.
Styrk honom att vara frimodig, ty han skall utskifta landet åt Israel såsom arv.
Och edra barn, om vilka I saden att de skulle bliva fiendens byte, och skola komma ditin, åt dem skall jag giva landet, och de skola taga det i besittning.
Men I själva mån vända eder åt annat håll; bryten nu upp och tagen vägen mot öknen, åt Röda havet till.»
Då svaraden I och saden till mig: »Vi hava syndat mot HERREN.
Vi vilja nu draga upp och strida, alldeles såsom HERREN, vår Gud, har bjudit oss.»
Och I omgjordaden eder, var och en tog sina vapen, och med lätt mod drogen I upp mot bergsbygden.
Men HERREN sade till mig: »Säg till dem: I skolen icke draga ditupp och giva eder i strid, ty jag är icke med bland eder; gören icke så, på det att I icke mån bliva slagna av edra fiender.»
Och jag talade till eder, men I hörden icke därpå, utan voren gensträviga mot HERRENS befallning och drogen i edert övermod upp mot bergsbygden.
Och amoréerna som bodde där i bergsbygden drogo mot eder och jagade eder, såsom bin göra, och slogo och förskingrade eder i Seir och drevo eder ända till Horma.
Då vänden I tillbaka och gräten inför HERRENS ansikte.
Men HERREN hörde icke eder röst och lyssnade icke till eder.
Och I stannaden länge i Kades, så länge det nu var.
Sedan vände vi oss åt annat håll, vi bröto upp och togo vägen mot öknen, åt Röda havet till, såsom Herren hade tillsagt mig, och vi höllo en lång tid på med att tåga omkring Seirs bergsbygd.
Och HERREN talade till mig och sade:
»Länge nog haven I hållit på med att tåga omkring denna bergsbygd; vänden eder nu mot norr.
Och bjud folket och säg: I kommen nu att draga fram genom det område som tillhör edra bröder, Esaus barn, vilka bo i Seir; men fastän de skola frukta för eder, mån I taga eder väl till vara.
I skolen icke inlåta eder i strid med dem, ty av deras land skall jag icke giva eder ens så mycket som en fotsbredd, eftersom jag redan har givit Seirs bergsbygd till besittning åt Esau.
Mat att äta skolen I köpa av dem för penningar; vatten att dricka skolen I ock köpa av dem för penningar.
HERREN, din Gud, har ju välsignat dig i alla dina händers verk; han har låtit sig vårda om din vandring i denna stora öken; nu i fyrtio år har HERREN, din Gud, varit med dig, och intet har fattats dig.
Så drog vi då åstad bort ifrån våra bröder, Esaus barn, som bodde i Seir, och lämnade Hedmarksvägen och Elat och Esjon-Geber.
Vi vände oss nu åt annat håll och drogo fram på vägen till Moabs öken.
Och Herren sade till mig: »Du skall icke angripa Moab eller inlåta dig i strid med dem, ty av deras land skall jag icke giva dig något till besittning, eftersom jag redan har givit Ar åt Lots barn till besittning.
(Eméerna bodde där fordom, ett stort och talrikt och resligt folk, sådant som anakiterna.
Och likasom anakiterna räknas också de för rafaéer; men moabiterna kalla dem eméer.
I Seir bodde däremot fordom horéerna, men Esaus barn fördrevo dem för sig och förgjorde dem och bosatte sig på det land som Herren hade givit dem till besittning.)
Stån nu upp och gån över bäcken Sered.»
Så gingo vi då över bäcken Sered.
Och den tid som åtgick för vår vandring från Kades-Barnea, till dess vi gingo över bäcken Sered. var trettioåtta år, och under denna tid förgicks hela den släktet, alla stridbara män i lägret, såsom Herren hade svurit att det skulle gå dem.
Ja, Herrens hand drabbade dem, och han sände förödelse i lägret bland dem och ryckte dem bort därur, så att de förgingos.
Då nu alla stridbara män i folket hade dött ut,
talade HERREN till mig och sade:
»Du drager nu över Moabs gräns, genom Ar,
och skall så komma i närheten av Ammons barn; men du må icke angripa dessa, ej heller inlåta dig i strid med dem, ty av Ammons barns land skall jag icke giva dig något till besittning, eftersom jag redan har givit det åt Lots barn till besittning.
(Såsom ett rafaéernas land räknas också detta; rafaéer bodde fordom där; men ammoniterna kalla dem samsummiter.
De voro ett stort och talrikt och resligt folk, sådant som anakiterna.
Men Herren förgjorde dessa för dem; de fördrevo dem och bosatte sig i deras land.
På samma sätt hade han gjort för Esaus barn, som bo i Seir, i det han för dem förgjorde horéerna; de fördrevo dem och bosatte sig i deras land, där de bo ännu i dag.
Likaså blevo avéerna, som bodde i byar ända fram till Gasa, förgjorda av kaftoréerna, som drogo ut från Kaftor och sedan bosatte sig i deras land.)
Stån nu upp, bryten upp och gån över bäcken Arnon.
Se, jag har givit Sihon, konungen i Hesbon, amoréen, och hans land i ditt våld.
Så begynn nu att intaga det, och bekriga honom.
Redan i dag vill jag begynna att låta förskräckelse och fruktan för dig komma över alla folk under himmelen, så att de skola darra och bäva för dig, när de höra berättas om dig.»
Och jag skickade sändebud från Kedemots öken till Sihon, konungen i Hesbon, med fridsam hälsning och lät säga:
»Låt mig tåga genom ditt land.
Raka vägen skall gå, utan att vika av vare sig till höger eller till vänster.
Mat att äta må du låta mig köpa för penningar; jag begär allenast att få tåga vägen fram härigenom
-- detsamma som tillstaddes mig av Esaus barn, Seirs inbyggare, och av moabiterna, Ars inbyggare -- så att jag kan gå över Jordan in i det land som HERREN, vår Gud, vill giva oss.»
Men Sihon, konungen i Hesbon, ville icke låta oss tåga genom sitt land, ty HERREN, din Gud, förhärdade hans sinne och förstockade hans hjärta, för att han skulle giva honom i din hand, såsom ock nu har skett.
Och Herren sade till mig: »Se, jag begynner nu att giva Sihon och hans land i ditt våld.
Begynn alltså du nu att intaga det, så att du får hans land till besittning.»
Och Sihon drog med allt sitt folk ut till strid mot oss, till Jahas.
Men HERREN, vår Gud, gav honom i vårt våld, och vi slogo honom jämte hans söner och allt hans folk.
Och vi intogo då alla hans städer och gåvo hela den manliga stadsbefolkningen till spillo, så ock kvinnor och barn; vi läto ingen slippa undan.
Allenast boskapen togo vi såsom byte, jämte rovet från de städer vi intogo.
Från Aroer, vid bäcken Arnons strand, och från staden i dalen ända till Gilead fanns ingen stad vars murar voro för höga för oss; allasammans gav HERREN, vår Gud, i vårt våld.
Men Ammons barns land lät du vara, hela landsträckan utefter bäcken Jabbok, och städerna i bergsbygden, och allt övrigt varom HERREN, vår Gud, hade så bjudit.
Sedan vände vi oss åt annat håll och drogo upp åt Basan till.
Och Og, konungen i Basan, drog med allt sitt folk ut i strid mot oss, till Edrei.
Men HERREN sade till mig: »Frukta icke för honom, ty i din hand har jag givit honom och allt hans folk och honom på samma sätt som du gjorde med Sihon, amoréernas konung, som bodde i Hesbon.»
Så gav HERREN, vår GUD, i vår hand också Og, konungen i Basan, och allt hans folk, och vi slogo honom och läto ingen av dem slippa undan.
Och vi intogo då alla hans städer, ingen stad fanns, som vi icke togo ifrån dem: sextio städer, hela landsträckan Argob, Ogs rike i Basan.
Alla dessa städer voro befästa med höga murar, med portar och bommar.
Därtill kom en stor mängd småstäder.
Och vi gåvo dem till spillo, likasom vi hade gjort med Sihon, konungen i Hesbon; hela den manliga stadsbefolkningen gåvo vi till spillo, så ock kvinnor och barn.
Men all boskapen och rovet från städerna togo vi såsom byte.
Från amoréernas två konungar, som härskade på andra sidan Jordan, togo vi alltså då deras land, från bäcken Arnon ända till berget Hermon
-- vilket av sidonierna kallas för Sirjon, men av amoréerna kallas för Senir --
alla städerna på slätten och hela Gilead och hela Basan, ända till Salka och Edrei, städerna i Ogs rike, i Basan.
Ty Og, konungen i Basan, var den ende som fanns kvar av de sista rafaéerna; hans gravkista, gjord av basalt, finnes, såsom känt är, i Rabba i Ammons barns land; den är nio alnar lång och fyra alnar bred, alnen beräknad efter längden av en mans underarm.
När vi då hade intagit detta land, gav jag den del därav, som sträcker sig från Aroer vid bäcken Arnon, samt hälften av Gileads bergsbygd med dess städer åt rubeniterna och gaditerna.
Återstoden av Gilead och hela Basan, Ogs rike, gav jag åt ena hälften av Manasse stam, hela landsträckan Argob, hela Basan; detta kallas rafaéernas land.
Jair, Manasses son, fick hela landsträckan Argob, ända till gesuréernas och maakatéernas område, och efter sitt eget namn kallade han landet -- nämligen Basan -- för Jairs byar, såsom det heter ännu i dag.
Och åt Makir gav jag Gilead.
Och åt rubeniterna och gaditerna gav jag landet från Gilead ända till Arnons dal, till dalens mitt -- den utgjorde gränsen -- och till bäcken Jabbok, som är Ammons barns gräns,
vidare Hedmarken med Jordan, som utgör gränsen, från Kinneret ända till Pisgas sluttningar, på östra sidan.
Och jag bjöd eder på den tiden och sade: »HERREN, eder Gud, har givit eder detta land till besittning.
Men nu skolen alla I som ären stridbara män draga väpnade åstad i spetsen för edra bröder, Israels barn.
Allenast edra hustrur och barn och eder boskap -- jag vet ju att I haven mycken boskap -- må stanna kvar i de städer som jag har givit eder,
till dess att HERREN har låtit edra bröder komma till ro, såväl som eder, när också de hava tagit i besittning det land som HERREN, eder Gud, vill giva dem på andra sidan Jordan; sedan mån I vända tillbaka till de besittningar jag har givit eder, var och en till sin besittning.»
Och jag bjöd Josua på den tiden och sade: »Du har med egna ögon sett allt vad HERREN, eder Gud, har gjort med dessa två konungar.
På samma sätt skall HERREN göra med alla riken där du drager fram.
Frukten icke för dem, ty HERREN, eder Gud, skall själv strida för eder.»
Och på den tiden bad jag till HERREN och sade:
»Herre, HERRE, du har begynt att låta sin tjänare se din storhet och din starka hand; ty vilken är den gud i himmelen eller på jorden, som kan göra sådana verk och sådana väldiga gärningar som du?
Så låt mig nu få gå ditöver och se det goda landet på andra sidan Jordan, det goda berglandet där och Libanon.»
Men HERREN hade blivit förgrymmad på mig för eder skull och ville icke höra mig, utan sade till mig: »Låt det vara nog; tala icke vidare till mig om denna sak.
Stig nu upp på toppen av Pisga, och lyft upp dina ögon mot väster och norr och söder och öster, och se med dina ögon; ty över denna Jordan skall du icke komma.
Och insätt Josua i hans ämbete, och styrk honom att vara frimodig och oförfärad; ty det är han som skall gå ditöver i spetsen för detta folk, och det är han som skall utskifta åt dem såsom arv det land du ser.»
Och så stannade vi i dalen mitt emot Bet-Peor.
Och nu, Israel, hör de stadgar och rätter som jag vill lära eder, för att I mån göra efter dem, på det att I mån leva och komma in i och taga i besittning det land som HERREN, edra fäders Gud, vill giva eder.
I skolen icke lägga något till det som jag bjuder eder, och I skolen icke taga något därifrån; I skolen hålla HERRENS, eder Guds, bud, som jag giver eder.
I haven med egna ögon sett vad HERREN har gjort i fråga om Baal-Peor, huru HERREN, din Gud, utrotade ur ditt folk var man som följde efter Baal-Peor.
Men I som höllen eder till HERREN, eder Gud, I leven alla ännu i dag.
Se, jag har lärt eder stadgar och rätter såsom HERREN, min Gud, har bjudit mig, på det att I mån göra efter dem i det land dit I nu kommen, för att taga det i besittning.
I skolen hålla dem och göra efter dem, ty det skall tillräknas eder såsom vishet och förstånd av andra folk.
När de få höra alla dessa stadgar, skola säga: »I sanning, ett vist och förståndigt folk är detta stora folk.»
Ty vilket annat stort folk finnes, vars gudar äro det så nära som HERREN, vår Gud, är oss, så ofta vi åkalla honom?
Och vilket annat stort folk finnes, som har stadgar och rätter så rättfärdiga som hela denna lag, vilken jag i dag förelägger eder?
Allenast tag dig till vara och akta dig väl, så att du icke förgäter vad dina ögon sågo, och icke låter vika ifrån ditt hjärta i all dina livsdagar, utan kungör det för dina barn och dina barnbarn:
vad som skedde den dag då du stod inför HERREN, din Gud, vid Horeb, då HERREN sade till mig: »Församla folket till mig, för att jag må låta dem höra mina ord; må de så lära sig att frukta mig, så länge de leva på jorden, och de lära sina barn detsamma.»
Och I trädden fram och blevo stående nedanför berget; och berget brann i eld ända upp till himmelen, och där var mörker, moln och töcken.
Och HERREN talade till eder ur elden orden hörden I, men I sågen ingen gestalt, I hörden allenast en röst.
Och han förkunnade eder sitt förbund, som han bjöd eder att hålla nämligen de tio orden; och han skrev dem på två stentavlor.
Och mig bjöd HERREN då att jag skulle lära eder stadgar och rätter, för att I skullen göra efter dem i det land dit I nu dragen, till att taga det i besittning.
Och eftersom I icke sågen någon gestalt den dag då HERREN talade till eder på Horeb ur elden, därför mån I nu noga hava akt på eder själva.
så att I icke tagen eder till, vad fördärvligt är, genom att göra eder någon beläte, något slags avgudabild, något bild av man eller av kvinna.
eller någon bild av något fyrfotadjur eller av någon bevingad fågel som flyger under himmelen,
eller av något kräldjur på marken eller av någon fisk i vattnet under jorden.
Och när du lyfter dina ögon upp till himmelen och ser solen, månen och stjärnorna, himmelens hela härskara, då må du icke heller låta förföra dig att tillbedja dem och tjäna dem; ty HERREN, din Gud, har givit dem åt alla folk under hela himmelen till deras del.
Men eder har HERREN tagit, och han har fört eder ut ur smältugnen, ur Egypten, för att I skullen bliva hans arvfolk, såsom nu har skett.
Och HERREN vredgades på mig för eder skull, och svor att jag icke skulle få gå över Jordan och komma in i de goda land som HERREN, din Gud, vill giva dig till arvedel.
Ty jag skall dö i detta land och icke gå över Jordan, men I skolen gå över den och taga detta goda land i besittning.
Tagen eder då till vara för att förgäta det förbund som HERREN, eder Gud, har slutit med eder, därigenom att I, alldeles emot HERRENS, eder Guds, bud, gören eder något beläte, något slags bild.
Ty, HERREN, din Gud, är en förtärande eld, en nitälskande Gud.
Om nu så sker, när du har fått barn och barnbarn och I haven blivit gamla i landet, att I tagen eder till, vad fördärvligt är, genom att göra eder något beläte, något slags bild, så att I gören vad som är ont i HERRENS, din Guds, ögon och därmed förtörnen honom,
då tager jag i dag himmel och jord till vittnen mot eder, att I med hast skolen förgås och utrotas ur det land dit I nu gån över Jordan, för att taga det i besittning; I skolen då icke längre leva där, utan skolen förvisso förgöras.
Och HERREN skall förströ eder bland folken, och allenast en ringa hop av eder skall bliva kvar bland de folk till vilka HERREN skall föra eder.
Och där skolen I tjäna gudar, gjorda av människohänder, gudar av trä och sten, som varken se eller höra eller äta eller lukta.
Men när I där söken HERREN, din Gud, då skall du finna honom, om du frågar efter honom av allt ditt hjärta och av all din själ.
När du är i nöd och allt detta vederfares dig, i kommande dagar, då skall du vända åter till HERREN, din Gud, och höra hans röst.
Ty HERREN, din Gud, är en barmhärtig Gud.
Han skall icke förgäta eller fördärva dig; han skall icke förgäta det förbund han har ingått med dina fäder och med ed bekräftat.
Ty fråga framfarna tider, dem som hava varit före dig, från den dag då Gud skapade människor på jorden, fråga ifrån himmelens ena ända till den andra om någonsin något så stort som detta har skett, eller om man har hört talas om något som är detta likt,
om något folk har hört Guds röst tala ur elden, såsom du har hört, och dock har blivit vid liv,
eller om någon gud har försökt att komma och hämta ett folk åt sig ut från ett annat folk, genom hemsökelser, tecken och under, genom krig, genom stark hand och uträckt arm, och genom stora, fruktansvärda gärningar, vilket allt HERREN, eder Guds, har gjort med eder i Egypten, inför dina ögon.
Du har själv fått se det, för att du skulle veta att HERREN är Gud, och ingen annan än han.
Från himmelen har han låtit dig höra sin röst för att undervisa dig, och på jorden har han låtit dig se sin stora eld, och du har hört hans ord ur elden.
Eftersom han nu älskade dina fäder och utvalde deras avkomlingar efter dem, och själv med sin stora kraft förde dig ut ur Egypten,
och fördrev för dig folk som voro större och mäktigare än du, och lät dig komma in i deras land och gav det åt dig till arvedel, såsom nu har skett,
därför skall du i dag veta och lägga på hjärtat att HERREN är Gud, uppe i himmelen och nere på jorden, han och ingen annan;
och du skall hålla hans stadgar och bud, som jag i dag giver dig, på det att det må gå dig väl och dina barn efter dig, och på det att du må länge leva i det land som HERREN, din Gud, vill giva dig för all tid.
Vid denna tid avskilde Mose tre städer på andra sidan Jordan, på östra sidan,
till vilka en dråpare skulle kunna fly, om han hade dräpt någon utan vett och vilja, och utan att förut hava burit hat till honom; om han flydde till någon av dessa städer, skulle han få bliva vid liv.
De voro: Beser i öknen på slättlandet för Rubens stam, Ramot i Gilead för Gads stam och Golan i Basan för Manasse stam.
Och detta är den lag som Mose förelade Israels barn,
dessa äro de vittnesbörd och stadgar och rätter som Mose föredrog för Israels barn, sedan de hade dragit ut ur Egypten,
på andra sidan Jordan i dalen, mitt emot Bet-Peor, i Sihons land, amoréernas konungs, som bodde i Hesbon, och som Mose och Israels barn slogo, när de hade dragit ut ur Egypten.
Ty de intogo hans land och Ogs land, konungens i Basan, amoréernas två konungars länder, på andra sidan Jordan, på östra sidan,
från Aroer vid bäcken Arnons strand ända till berget Sion, det är Hermon,
och hela Hedmarken på andra sidan Jordan på östra sidan, ända till Hedmarkshavet, nedanför Pisgas sluttningar.
Och Mose sammankallade hela Israel och sade till dem: Hör, Israel, de stadgar och rätter som jag i dag framställer för eder, och lären eder dem och hållen dem och gören efter dem.
HERREN, vår Gud, slöt ett förbund med oss på Horeb.
Icke med våra fäder slöt HERREN detta förbund, utan med oss själva som stå här i dag, oss alla som nu leva.
Ansikte mot ansikte talade HERREN till eder på berget ur elden.
Jag stod då mellan HERREN och eder, för att förkunna eder vad HERREN talade, ty I fruktaden för elden och stegen icke upp på berget.
Han sade:
Jag är HERREN, din Gud, som har fört dig ut ur Egyptens land, ur träldomshuset.
Du skall inga andra gudar hava jämte mig.
Du skall icke göra dig något beläte, som är en bild vare sig av det som är uppe i himmelen, eller av det som är i vattnet under jorden.
Du skall icke tillbedja sådana, ej heller tjäna dem; ty jag, HERREN, sin Gud, är en nitälskande Gud, som hemsöker fädernas missgärning på barn och efterkommande i tredje och fjärde led, när man hatar mig,
men som gör nåd med tusenden, när man älskar mig och håller mina bud.
Du skall icke missbruka HERRENS, din Guds namn, ty HERREN skall icke låta den bliva ostraffad, som missbrukar hans namn.
Håll sabbatsdagen, så att du helgar den, såsom HERREN, din Gud, har bjudit dig.
Sex dagar skall du arbeta och förrätta alla dina sysslor;
men den sjunde dagen är HERRENS, din Guds, sabbat; då skall du ingen syssla förrätta, ej heller din son eller sin dotter, eller din tjänare eller din tjänarinna, eller din oxe eller din åsna eller någon av dina dragare, ej heller främlingen som är hos dig inom dina portar; på det att din tjänare och din tjänarinna må hava ro såväl som du.
Du skall komma ihåg att du själv har varit träl i Egyptens land, och att HERREN, din Gud, har fört dig ut därifrån med stark hand och uträckt arm; därför har HERREN, din Gud bjudit dig att hålla sabbatsdagen.
Hedra din fader och din moder, såsom HERREN, din Gud har bjudit dig, på det att du må länge leva och det må gå dig väl i det land som HERREN, din Gud, vill giva dig.
Du skall icke dräpa.
Du skall icke heller begå äktenskapsbrott.
Du skall icke heller stjäla.
Du skall icke heller bära falsk vittnesbörd mot din nästa.
Du skall icke heller hava begärelse till din nästas hustru.
Du skall icke heller hava lust till din nästas hus, ej heller till hans åker eller hans tjänare eller hans tjänarinna, ej heller till hans oxe eller hans åsna, ej heller till något som tillhör din nästa.
Dessa ord talade HERREN till hela eder församling på berget, ur elden, molnskyn och töcknet, med hög röst, och han talade så intet mer.
Och han skrev dem på två stentavlor, som han gav åt mig.
När I hörden rösten ur mörkret, medan berget brann i eld, trädden I fram till mig, alla I som voren huvudmän för edra stammar, så ock edra äldste.
Och I saden: »Se, HERREN, vår Gud, har låtit oss se sin härlighet och sin storhet, och vi hava hört hans röst ur elden.
I dag hava vi sett att Gud kan tala med en människa och dock låta henne bliva vid liv.
Varför skola vi då likväl dö?
Denna stora eld kommer ju att förtära oss.
Om vi än vidare få höra HERRENS, vår Guds, röst, så måste vi dö.
Ty vem finnes väl bland allt kött som kan, såsom vi hava gjort, höra den levande Gudens röst tala ur elden och dock bliva vid liv?
Träd du fram och hör allt vad HERREN, vår Gud, säger, och tala du till oss allt vad HERREN, vår Gud, talar till dig, så vilja vi höra det och göra därefter.»
Och HERREN hörde edra ord, när I så taladen till mig; och HERREN sade till mig: »Jag har hört de ord som detta folk har talat till dig.
De hava rätt i allt vad de hava talat.
Ack att de hade sådana hjärtan, att de fruktade mig och hölle alla mina bud alltid!
Det skulle ju då gå dem och deras barn väl evinnerligen.
Gå nu och säg till dem: 'Vänden tillbaka till edra tält.'
Men du själv må stanna kvar här hos mig, så skall förkunna för dig alla de bud och stadgar och rätter som du skall lära dem, för att de må göra efter dem i det land som jag vill giva dem till besittning.»
Så hållen nu och gören vad HERREN, eder Gud, har bjudit eder.
I skolen icke vika av vare sig till höger eller till vänster.
På de vägar som HERREN, eder Gud, har bjudit eder gå skolen I alltid vandra, för att I mån bliva vid liv och det må gå eder väl, och för att I mån länge leva i det land som I skolen taga i besittning.
Och dessa äro de bud, stadgar och rätter som HERREN, eder Gud, har bjudit mig att lära eder, för att I skolen göra efter dem i det land dit I nu dragen, till att taga de i besittning --
detta på det att du må frukta HERREN, din Gud, så att du håller alla hans stadgar och bud, som jag giver dig, du med din som och din sonson, i all dina livsdagar, och på det att du må länge leva.
Så skall du nu höra, Israel, och hålla dem och göra efter dem, för att det må gå dig väl, och för att I mån föröka eder mycket, såsom HERREN, dina fäders Gud, har lovat dig -- ett land som flyter av mjölk och honung.
Hör, Israel!
HERREN, vår gud, HERREN är en.
Och du skall älska HERREN, din Gud, av allt ditt hjärta och av all din själ och av all din kraft.
Dessa ord som jag i dag giver dig skall du lägga på ditt hjärta.
Och du skall inskärpa dem hos dina barn och tala om för dem, när du sitter i ditt hus och när du går på vägen, när du lägger dig och när du står upp.
Och du skall binda dem såsom ett tecken på din hand, och de skola vara såsom ett märke på din panna.
Och du skall skriva dem på dörrposterna i ditt hus och på dina portar.
När nu HERREN, din Gud, låter dig komma in i det land som han med ed har lovat dina fäder, Abraham, Isak och Jakob, att giva dig -- stora och vackra städer, som du icke har byggt,
och hus, fulla med allt gott, vilka du icke har fyllt, och uthuggna brunnar, som du icke har huggit ut, vingårdar och olivplanteringar, som du icke har planterat -- och när du då äter och bliver mätt,
så tag dig till vara för att förgäta HERREN, som har fört dig ut ur Egyptens land, ur träldomshuset.
HERREN, din Gud, skall du frukta, och honom skall du tjäna, och vid hans namn skall du svärja.
I skolen icke följa efter andra gudar, någon av de folks gudar, som bo runt omkring eder,
ty en nitälskande Gud är HERREN, din Gud, mitt ibland dig, och du må taga dig till vara, så att icke HERRENS, din Guds, vrede upptändes mot dig, och han utrotar dig från jorden.
I skolen icke fresta HERREN, eder Gud, såsom I frestaden honom i Massa.
I skolen troget hålla HERRENS, eder Guds, bud och de vittnesbörd och stadgar som han hat givit dig.
Och du skall göra vad rätt och gott är i HERRENS ögon, för att det må gå dig väl, och för att du må komma in i det goda land som HERREN med ed har lovat åt dina fäder, och taga det i besittning,
därigenom att han driver undan för dig all dina fiender, såsom HERREN har lovat.
När din son i framtiden frågar dig: »Vad betyda de vittnesbörd och stadgar och rätter som HERREN, vår Gud, har givit eder?»
då skall du svara din son: »Vi voro Faraos trälar i Egypten, men med stark hand förde HERREN oss ut ur Egypten.
Och HERREN gjorde stora och gruvliga tecken och under i Egypten på Farao och hela hans hus inför våra ögon.
Men oss förde han ut därifrån, för att låta oss komma in och giva oss det land som han med ed har lovat åt våra fäder.
Och HERREN bjöd oss att göra efter all dessa stadgar och att frukta HERREN, vår Gud, för att det alltid skulle gå oss väl, i det att han behölle oss vid liv, såsom ock hittills har skett.
Och det skall lända oss till rättfärdighet, när vi hålla och göra efter alla dessa bud, inför HERREN, vår Guds, ansikte, såsom han har bjudit oss.»
När HERREN, din Gud låter dig komma in i det land di du nu går, för att taga i besittning, och när han för dig förjagar stora folk -- hetiterna, girgaséerna, amoréerna, kananéerna, perisséerna, hivéerna och jebuséerna, sju folk, större och mäktigare än du --
när HERREN, din Gud, giver dessa i ditt våld och du slår dem, då skall du giva dem till spillo; du skall icke sluta förbund med dem eller visa dem nåd.
Du skall icke befrynda dig med dem; dina döttrar skall du icke giva åt deras söner, och deras döttrar skall du icke taga till hustrur åt dina söner.
Ty de skola då förleda dina söner att vika av ifrån mig och tjäna andra gudar, och HERRENS vrede skall då upptändas mot eder och han skall med hast förgöra dig.
Utan så skolen I göra med dem I skolen bryta ned deras altaren och slå sönder deras stoder och hugga ned deras Aseror och bränna upp deras beläten i eld.
Ty du är ett folk som är helgat åt HERREN, din Gud; dig har HERREN, din Gud, utvalt till att vara hans egendomsfolk, framför alla andra folk på jorden.
Icke därför att I voren större än alla andra folk var det som HERREN fäste sig vid eder och utvalde eder, ty I ären ju mindre än alla andra folk;
utan därför att HERREN älskade eder och ville hålla den ed som han hade svurit fäder, därför förde HERREN eder ut med stark hand och förlossade dig ur träldomshuset, ur Faraos, den egyptiske konungens, hand.
Så skall du nu veta att HERREN, din Gud, är den rätte Guden, den trofaste Guden, som håller förbund och bevarar nåd intill tusende led, när man älskar honom och håller hans bud,
men som utan förskoning vedergäller och förgör dem som hata honom.
Han dröjer icke, när det gäller dem som hata honom; utan förskoning vedergäller han dem.
Så håll nu de bud och stadgar och rätter som jag i dag giver dig, och gör efter dem.
Om I nu hören dessa rätter och hållen dem och gören efter dem, så skall HERREN, din Gud, till lön därför låta sitt förbund och sin nåd bestå, vad han med ed lovade dina fäder.
Han skall då älska dig och välsigna sitt livs frukt och din marks frukt, din säd, ditt vin och din olja, dina fäkreaturs avföda och din småboskaps avel, i det land som han med ed har lovat dina fäder att giva dig.
Välsignad skall du bliva framför alla andra folk; bland dina män och kvinnor skall ingen vara ofruktsam, ej heller bland din boskap.
Och HERREN skall avvända från dig all krankhet; ingen av Egyptens alla svåra sjukdomar, som du väl känner, skall han lägga på dig; han skall i stället låta dem komma över alla dem som hata dig.
Och alla de folk som HERREN, din Gud, giver i din hand skall du utrota; du skall icke visa dem någon skonsamhet.
Du skall icke heller tjäna deras gudar, ty detta kunde bliva en snara för dig.
Om du ock säger vid dig själv: »Dessa folk äro större än jag; huru skall jag kunna fördriva dem?»,
så må du dock icke frukta för dem; du skall tänka på vad HERREN, din Gud gjorde med Farao och med all egyptierna,
på de stora hemsökelser som du med egna ögon såg, och på de tecken och under och på den starka hand och uträckta arm varmed HERREN, din Gud, förde dig ut.
På samma sätt skall HERREN, din Gud, nu göra med alla de folk som du fruktar för.
Därtill skall HERREN, din Gud, sända getingar över dem, till dess att de som äro kvar och hålla sig gömda för dig hava blivit utrotade.
Du må icke förskräckas för dem, ty HERREN, din Gud, är mitt ibland dig, en stod och fruktansvärd Gud.
Och HERREN, din Gud, skall förjaga dessa hedningar för dig, men blott småningom.
Du skall icke med hast få förgöra dem, på det att vilddjuren icke må föröka sig till din skada.
HERREN, din Gud, skall giva dem i ditt våld och sända stor förvirring bland dem, till dess att de förgöras.
Och han skall giva deras konungar i din hand, och du skall utrota till och med deras namn, så att de icke mer finnas under himmelen.
Ingen skall kunna stå dig emot, till dess du har förgjort dem.
Deras gudabeläten skola I bränna upp i eld.
Du skall icke hava begärelse till det silver och det guld som finnes på dem, och icke taga något av detta för din räkning, på det att du icke må snärjas därav; ty en styggelse är det för HERREN, din Gud.
Och du skall icke låta någon styggelse komma in i ditt hus, på det att du icke också själv må bliva given till spillo.
Du skall räkna det såsom en skändlighet och en styggelse, ty det är givet till spillo.
Alla de bud som jag i dag giver dig skolen I hållen, och efter dem skolen I göra, för att I mån komma in i och taga i besittning det land som HERREN med ed har lovat åt edra fäder.
Och du skall komma ihåg allt vad som har skett på den väg HERREN, din Gud, nu i fyrtio åt har låtit dig vandra i öknen, för att tukta dig och pröva dig, så att han kunde förnimma vad som var i ditt hjärta: om du ville hålla hans bud eller icke.
Ja, han tuktade dig och lät dig hungra, och han gav dig manna att äta, en mat som du förut icke visste av, och som icke heller dina fäder visste av; på det att han skulle lära dig förstå att människan lever icke allenast av bröd, utan att hon lever av allt det som utgår av HERRENS mun.
Dina kläder blevo icke utslitna på dig, och din fot svullnade icke under dessa fyrtio år.
Så skall du då förstå i ditt hjärta att HERREN, din Gud, fostrar dig, såsom en man fostrar sin son;
och du skall hålla HERRENS, din Guds, bud, så att du vandrar på hans vägar och fruktar honom.
Ty HERREN, din Gud, låter dig nu komma in i ett gott land, ett land där vattenbäckar, källor och djupa vatten flöda fram i dalar och på berg,
ett land med vete och korn, med vinträd, fikonträd och granatträd, ett land med ädla olivträd och med honung,
ett land där du icke skall äta ditt bröd i torftighet, där intet skall fattas dig, ett land vars stenar innehålla järn, och ur vars berg du skall bryta koppar.
Där skall du äta och bliva mätt, och du skall så lova HERREN, din Gud, för det goda land som han har givit dig.
Tag dig då till vara för att förgäta HERREN, din Gud, så att du icke håller hans bud och rätter och stadgar, som jag i dag giver dig.
Ja, när du äter och bliver mätt, och bygger vackra hus och bor i dem,
när dina fäkreatur och din småboskap förökas, och ditt silver och guld förökas, och allt annat du har förökas,
då må ditt hjärta icke bliva högmodigt, så att du förgäter HERREN, din Gud, som har fört dig ut ur Egyptens land, ur träldomshuset.
och som har lett dig genom den stora och fruktansvärda öknen, bland giftiga ormar och skorpioner, över förtorkad mark, där intet vatten åt dig komma ut ur den hårda klippan,
och som gav dig manna att äta i öknen, en mat som dina fäder icke visste av -- detta på det att han skulle tukta dig och pröva dig, för att sedan kunna göra dig gott.
Du må icke säga vid dig själv: »Min egen kraft och min hands styrka har förskaffat mig denna rikedom»,
utan du må komma ihåg att det är HERREN, din Gud, som giver dig kraft att förvärva rikedom, därför att han vill upprätta det förbund som han med ed har ingått med dina fäder -- såsom och hittills har skett.
Men om du förgäter HERREN, din Gud, och följer efter andra gudar och tjänar dem och tillbeder dem, så betygar jag i dag inför eder att I förvisso skolen förgås.
På samma sätt som hedningarna som HERREN förgör för eder skolen också I då förgås, därför att I icke hörden HERRENS, eder Guds röst.
Hör, Israel!
Du går nu över Jordan, för att komma ditin och underlägga dig folk, större och mäktigare än du, städer, stora och befästa upp mot himmelen,
anakiternas stora och resliga folkstam, som du själv känner, och om vilken du har hört att man säger: »Vem kan stå emot Anaks barn!»
Så skall du nu veta att HERREN, din Gud, är den som går framför dig, såsom en förtärande eld; han skall förgöra dem, och han skall förgöra dem, och han skall ödmjuka dem för dig, och du skall fördriva dem och utrota dem med hast, såsom HERREN har lovat dig.
Då nu HERREN, din Gud, driver dem undan för dig, må du icke säga vid dig själv: »För min rättfärdighets skull har HERREN låtit mig komma in i detta land och taga det i besittning.»
Ty dessa hedningars ogudaktighet är det som gör att HERREN fördriver dem för dig.
Icke din rättfärdighet och din rättsinnighet är det som gör att du får komma in i deras land och taga det i besittning, utan dessa hedningars ogudaktighet är det som gör att HERREN, din Gud, fördriver dem för dig.
Så vill ock HERREN uppfylla vad han med ed har lovat dina fäder, Abraham, Isak och Jakob.
Därför må du nu veta att det icke är din rättfärdighet som gör att HERREN, din Gud, vill giva dig detta goda land till besittning; ty du är ett hårdnackat folk.
Kom ihåg, förgät icke, huru du i öknen förtörnade HERREN, din Gud.
Allt ifrån den dag då du drog ut ur Egyptens land, ända till dess I nu haven kommit hit, haven I varit gensträviga mot HERREN.
Vid Horeb förtörnaden I HERREN, och HERREN vredgades på eder, så att han ville förgöra eder.
När jag hade stigit upp på berget för att taga emot stentavlorna, det förbunds tavlor, som HERREN hade slutit med eder, stannade jag på berget i fyrtio dagar och fyrtio nätter, utan att äta och utan att dricka.
Och HERREN gav mig de två stentavlorna, på vilka Gud hade skrivit med sitt finger; vad där stod var alldeles lika med de ord HERREN hade talat med eder på berget ur elden, den dag då I voren församlade där.
Och när de fyrtio dagarna och de fyrtio nätterna voro förlidna, gav HERREN mig de två stentavlorna, förbundets tavlor.
Och HERREN sade till mig: »Stå upp och gå med hast ned härifrån, ty ditt folk, som du har fört ut ur Egypten, har tagit sig till, vad fördärvligt är.
De hava redan vikit av ifrån den väg som jag bjöd dem gå; de hava gjort sig ett gjutet beläte.»
Och HERREN talade till mig och sade: »jag har sett att detta folk är ett hårdnackat folk.
Lämna mig i fred, ty jag vill förgöra dem och utplåna deras namn, så att det icke mer finnes under himmelen; dig vill jag sedan göra till ett folk som är mäktigare och större än detta.»
Då vände jag mig om och steg ned från berget, som brann i eld; och jag hade i mina båda händer förbundets två tavlor.
Och jag fick då se att I haven syndat mot HERREN, eder Gud: I haden gjort eder en gjuten kalv; så haden I redan vikit av ifrån den väg som HERREN hade bjudit eder gå.
Då fattade jag i de båda tavlorna och kastade dem ifrån mig med båda händerna och slog sönder dem inför edra ögon.
Och jag föll ned inför HERRENS ansikte och låg så, likasom förra gången i fyrtio dagar och fyrtio nätter, utan att äta och utan att dricka, för all den synds skulle som I haden begått genom att göra vad ont var i HERRENS ögon, till att förtörna honom.
Ty jag fruktade för den vrede och förbittring mot eder, av vilken HERREN hade blivit så uppfylld att han ville förgöra eder.
Och HERREN hörde mig även denna gång.
Också på Aron blev HERREN mycket vred, så att han ville förgöra honom, och jag bad då jämväl för Aron.
Sedan tog jag kalven, syndabelätet som I haden gjort, och brände den i eld och krossade sönder den väl, till dess att den blev fint stoft, och det stoftet kastade jag i bäcken som flöt ned från berget.
I Tabeera, i Massa och i Kibrot-Hattaava förtörnaden I ock HERREN.
Och när HERREN ville sända eder åstad från Kades-Barnea och sade: »Dragen upp och intagen det land som jag har givit eder», då voren I gensträviga mot HERREN, eder Guds, befallning och trodden honom icke och hörden icke hans röst.
Ja, gensträviga haven I varit mot HERREN allt ifrån den dag då jag lärde känna eder.
Så föll jag då ned inför HERRENS ansikte och låg så i de fyrtio dagarna och de fyrtio nätterna; ty HERREN hade sagt att han ville förgöra eder.
Och jag bad till HERREN och sade: »Herre, HERRE, fördärva icke ditt folk och din arvedel, som du har förlossat med din stora makt, och som du med stark hand har fört ut ur Egypten.
Tänk på dina tjänare Abraham, Isak och Jakob, se icke på detta folks hårdhet, ogudaktighet och synd;
på det att man icke må säga i det land varur du har fört oss ut: 'Därför att HERREN, icke förmådde föra dem in i det land som han hade lovat åt dem, och därför att han hatade dem, förde han dem ut och lät dem dö i öknen.'
De äro ju ditt folk och din arvedel, som du har fört ut med din stora kraft och din uträckta arm.»
På den tiden sade HERREN till mig: »Hugg ut åt dig två stentavlor, likadana som de förra voro, och stig upp till mig på berget; gör dig och en ark av trä.
Och sedan jag har skrivit på tavlorna samma ord som stodo på de förra tavlorna, vilka du slog sönder, skall du lägga dem i arken.»
Så gjorde jag då en ark av akacieträ och högg ut två stentavlor, likadana som de förra voro.
Och jag steg upp på berget och hade med mig de två tavlorna.
Och han skrev på tavlorna detsamma som var skrivet förra gången, de tio ord som HERREN hade talat till eder på berget ur elden, den dag då I voren församlade där.
Och HERREN gav dem åt mig.
Sedan vända jag mig om och steg ned från berget och lade tavlorna i arken som jag hade gjort, och där fingo de ligga, såsom HERREN hade bjudit mig.
Och Israels barn bröto upp från Beerot-Bene-Jaakan och tågade till Mosera.
Där dog Aron och blev där också begraven; och hans som Eleasar blev präst i hans ställe.
Därifrån bröto de upp och tågade till Gudgoda, och från Gudgoda, och från Gudgoda till Jotbata, en trakt som var rik på vattenbäckar.
På den tiden avskilde HERREN Levi stam till att bära HERRENS förbundsark, till att stå inför HERRENS ansikte och göra tjänst inför honom, och till att välsigna i hans namn, såsom den har att göra ännu i dag.
Därför fick Levi ingen lott eller arvedel jämte sina bröder.
HERREN är hans arvedel, såsom HERREN, din Gud, har sagt honom.
Och jag stannade på berget lika länge som förra gången, fyrtio dagar och fyrtio nätter; och HERREN hörde mig också denna gång: HERREN ville icke fördärva mig.
Och HERREN sade till mig: »Stå upp och gå åstad framför folket, och låt dem bryta upp, för att de må komma in i och taga i besittning det land som jag med ed har lovat deras fäder att giva dem.»
Och nu Israel, var är det som HERREN, din Gud, fordrar av dig annat än att du fruktar HERREN, din Gud, att du alltid vandrar på hans vägar och älskar honom, och att du tjänar HERREN, din Gud, av allt ditt hjärta och av all din själ,
så att du håller HERRENS bud och stadgar, som jag i dag giver dig, på det att det må gå dig väl?
Se, HERREN, din Gud, tillhör himlarna och himlarnas himmel, jorden och allt vad därpå är;
men allenast vid dina fäder fäste sig HERREN och älskade dem; och han utvalde deras avkomlingar efter dem, han utvalde eder bland alla folk, såsom I nu själva sen.
Omskären därför edert hjärtas förhud, och varen icke länge hårdnackade.
Ty HERREN, eder Gud, är gudarnas Gud och herrarnas Herre, den store, den väldige och fruktansvärde Guden, som icke har anseende till personen och icke tager mutor;
som skaffar den faderlöse och änkan rätt, och som älskar främlingen och giver honom mat och kläder.
Därför skolen också I älska främlingen; I haven ju själva varit främlingar i Egyptens land.
HERREN, din Gud, skall du frukta, honom skall du tjäna, och till honom skall du hålla dig, och vid hans namn skall du svärja.
Han är ditt lov, och han din Gud, som har gjort med dig de stora och underbara gärningar som du med egna ögon har sett.
Sjuttio personer voro dina fäder, som drogo ned till Egypten, men nu har HERREN, din Gud, gjort dig talrik såsom himmelens stjärnor.
Så skall du nu älska HERREN, din Gud, och hålla vad han bjuder dig hålla, hans stadgar och rätter och bud, alltid.
Och besinnen i dag -- jag talar nu icke om edra barn, som icke hava förnummit och sett det -- huru HERREN, eder Gud, har fostrat eder, besinnen hans storhet, hans starka hand och hans uträckta arm,
de tecken och gärningar som han gjorde i Egypten, med Farao, konungen i Egypten, och med hela hans land,
och vad han gjorde med egyptiernas här, med deras hästar och vagnar, huru han lät Röda havets vatten strömma över dem, när de förföljde eder, och huru HERREN då förgjorde dem, så att de nu icke mer äro till;
och vad han gjorde med eder i öknen, ända till dess I kommen hit,
och vad han gjorde med Datan och Abiram, Eliabs, Rubens sons, söner, huru jorden öppnade sin mun och uppslukade dem med deras hus och deras tält och allt levande som följde dem, och detta mitt i hela Israel.
Ty I haven ju med egna ögon sett alla de stora gärningar som HERREN har gjort.
Så hållen då alla de bud som jag i dag giver dig, på det att I med frimodighet mån kunna gå in i och intaga det land dit I nu dragen, för att taga det i besittning,
och på det att I mån länge leva i det land som HERREN med ed har lovat edra fäder att giva åt dem och deras efterkommande, ett land som flyter av mjölk och honung.
Ty det land dit du nu kommer, för att taga det i besittning, är icke såsom Egyptens land, varifrån I haven dragit ut, där du måste trampa upp vatten till den säd du sådde, såsom man gör i en köksträdgård;
nej, det land dit I nu dragen, för att taga det i besittning, är ett land med berg och dalar, som får vatten att dricka genom himmelens regn,
ett land som HERREN, din Gud, låter sig vårda om, och på vilket HERRENS, din Guds, ögon beständigt vila, från årets begynnelse till årets slut.
Om i nu hören de bud som jag i dag giver eder, så att I älsken HERREN, eder Gud, och tjänen honom av allt edert hjärta och av all eder själ,
så skall jag giva åt edert land regn i rätt tid, höstregn och vårregn, och du skall få inbärga din säd och ditt vin och din olja.
Och jag skall giva din boskap gräs på din mark; och du skall äta och bliva mätt.
Men tagen eder till vara, låten icke edra hjärtan bliva förförda, så att I viken av och tjänen andra gudar och tillbedjen dem;
ty då skall HERRENS vrede upptändas mot eder, och han skall tillsluta himmelen, så att regn icke faller och marken icke giver sin gröda; och I skolen med hast bliva utrotade ur det goda land som HERREN vill giva eder.
Så skolen I nu lägga dessa mina ord på edert hjärta och edert sinne, och I skolen binda dem såsom ett tecken på eder hand, och de skola vara såsom ett märke på eder panna;
och I skolen lära edra barn dem, i det att du talar om dem, när du sitter i ditt hus och när du står upp.
och du skall skriva dem på dörrposterna i ditt hus och på dina portar;
på det att I och edra barn mån länge få bo i det land som HERREN med ed har lovat edra fäder att giva dem, lika länge som himmelen välver sig över jorden.
Ty om I hållen alla dessa bud som jag giver eder och gören efter dem, så att I älsken HERREN, eder Gud, och alltid vandren på hans vägar och hållen eder till honom,
då skall HERREN fördriva alla dessa folk för eder, och I skolen underlägga eder folk som äro större och mäktigare än I.
Var ort eder fot beträder skall bliva eder.
Från öknen till Libanon, ifrån floden -- floden Frat -- ända till Västra havet skall edert område sträcka sig.
Ingen skall kunna stå eder emot.
Fruktan och förskräckelse för eder skall HERREN, eder Gud, låta komma över hela det land I beträden, såsom han har lovat eder.
Se, jag förelägger eder i dag välsignelse och förbannelse:
välsignelse, om I hören HERRENS eder Guds, bud, som jag i dag giver eder,
och förbannelse, om I icke hören HERRENS, eder Guds, bud, utan viken av ifrån den väg jag i dag bjuder eder gå och följen efter andra gudar, som I icke kännen.
Och när HERREN, din Gud, har låtit dig komma in i det land dit du nu går, för att taga det i besittning, skall du låta berget Gerissim bliva platsen för välsignelsen och berget Ebal platsen för förbannelsen.
(Dessa berg ligga, såsom känt är, på andra sidan Jordan, bortom Västra vägen, i hedmarkskananéernas land, mitt emot Gilgal, bredvid Mores terebintlund.)
Ty I gån nu över Jordan, för att komma in i och taga i besittning det land som HERREN, eder Gud, vill giva eder; I skolen taga det i besittning och bo där.
Hållen då alla de stadgar och rätter som jag i dag förelägger eder, och gören efter dem.
Dessa äro de stadgar och rätter som I skolen hålla och iakttaga i det land som HERREN, dina fäders Gud, har givit dig till besittning; så länge I leven på jorden skolen I hålla dem.
I skolen i grund föröda alla platser där de folk som I fördriven hava hållit sin gudstjänst, vare sig detta har skett på höga berg och höjder eller någonstädes under gröna träd.
I skolen bryta ned deras altaren och slå sönder deras stoder och bränna upp deras Aseror i eld och hugga ned deras gudabeläten, och I skolen utrota deras namn från sådana platser.
När I tillbedjen HERREN, eder Gud, skolen I icke göra såsom de,
utan den plats som HERREN, eder Gud, utväljer inom någon av edra stammar till att där fästa sitt namn, denna boning skolen I söka och dit skall du gå.
Och dit skolen I föra edra brännoffer och slaktoffer, eder tionde, vad edra händer bära fram såsom offergärd, edra löftesoffer och frivilliga offer och det förstfödda av edra fäkreatur och eder småboskap.
Och där skolen I äta inför HERRENS, eder Guds, ansikte, och glädja eder med edert husfolk över allt vad I haven förvärvat, allt varmed HERREN, din Gud, vara rättast;
I skolen då icke göra såsom vi nu göra här, var och en vad honom tyckes vara rättast.
I haven ju ännu icke kommit till ro och till den arvedel som HERREN, din Gud, vill giva dig.
Men när I haven gått över Jordan och bon i det land som HERREN, eder Gud, vill giva eder till arvedel, och när han har låtit eder få ro för alla edra fiender runt omkring, då att I bon i trygghet,
då skolen I till den plats som HERREN, eder Gud, utväljer till boning åt sitt namn föra allt vad jag nu bjuder eder: edra brännoffer och slaktoffer, eder tionde, vad edra händer bära fram såsom offergärd, så ock alla de utvalda löftesoffer som I loven HERREN.
Och så skolen I glädja eder inför HERREN, eder Guds, ansikte, med edra söner och döttrar, edra tjänare och tjänarinnor, och med leviten som bor inom edra portar, ty han har ju ingen lott eller arvedel med eder.
Tag dig till vara för att offra dina brännoffer på någon annan plats som kan falla din in;
nej, på den plats HERREN utväljer inom en av dina stammar, där skall du offra dina brännoffer, och där skall du göra allt vad jag eljest bjuder dig.
Dock får du, så mycket dig lyster, slakta och äta kött inom vilken som helst av dina städer, i mån av den välsignelse som HERREN, din Gud, giver dig.
Både den som är oren och den som är ren må äta därav, såsom vore det gasell- eller hjortkött.
Men blodet skolen I icke förtära I skolen gjuta ut det på jorden såsom vatten.
Du får alltså icke hemma inom dina portar äta tionde av din säd, ditt vin och din olja, ej heller det förstfödda av dina fäkreatur och din småboskap, ej heller något av de löftesoffer som du lovar, eller av dina frivilliga offer, eller av det din hand bär fram såsom offergärd;
utan inför HERREN, din Guds, ansikte, på den plats som HERREN, din Gud, utväljer skall du äta sådant, med din son och din dotter, din tjänare och din tjänarinna, och med leviten som bor inom dina portar; och så skall du glädja dig inför HERRENS, din Guds, ansikte över allt vad du har förvärvat.
Tag dig till vara för att glömma bort leviten, så länge du lever i ditt land.
Om du alltså, när HERREN, din Gud, har utvidgat ditt område, såsom han har lovat dig, tänker så: »Jag vill äta kött» -- ifall det nu lyster för dig att äta kött -- så må du då äta kött, så mycket dig lyster.
Om den plats som HERREN, din Gud, utväljer till att där fästa sitt namn ligger för avlägset för dig, så må du, i enlighet med vad jag har bjudit dig, slakta av de fäkreatur och av den småboskap som HERREN har givit dig, och äta därav hemma inom dina portar, så mycket av din lyster.
Men du skall äta på samma sätt som man äter gasell- eller hjortkött; både den som är oren och den som är ren må äta därav.
Allenast skall du vara ståndaktig i att icke förtära blodet; ty blodet är själen, och själen skall du icke förtära med köttet.
Du skall icke förtära det; du skall gjuta ut det på jorden såsom vatten.
Du skall icke förtära det, på det att det må gå dig väl och dina barn efter dig, när du göra vad rätt är i HERRENS ögon.
Men de heliga gåvor som du vill bära fram, och dina löftesoffer, dem skall du föra med dig till den plats som HERREN utväljer.
Och av dina brännoffer skall du offra både köttet och blodet på HERRENS, din Guds, altare.
Av dina slaktoffer däremot skall väl blodet gjutas ut på HERRENS, din Guds, altare, men köttet må du äta.
Alla dessa bud som jag giver dig skall du hålla och höra, för att det må gå dig väl och dina barn efter dig, till evig tid, när du gör var gott och rätt är i HERRENS, din Guds, ögon.
När HERREN, din Gud, har utrotat de folk till vilka du nu kommer, för att fördriva dem för dig, när du alltså har fördrivit dessa och bosatt dig i deras land,
tag dig då till vara för att bliva snärjd, så att du efterföljer dem, sedan de hava blivit förgjorda för dig; fråga icke efter deras gudar, så att du säger: »På vad sätt höllo dessa folk sin gudstjänst?
Så vill också jag göra.»
Nej, på det sättet skall icke du göra, när du tillbeder HERREN, din Gud, ty allt som är en styggelse för HERREN, och som han hatar, det hava de gjort till sina gudars ära; ja, de gå så långt att de bränna upp sina söner och döttrar i eld åt sina gudar.
Allt vad jag bjuder eder, det skolen I hålla och göra.
Du skall icke lägga något därtill och icke taga något därifrån.
Om en profet eller en som har drömmar uppstår bland dig, och han utlovar åt dig något tecken eller under,
och sedan det tecken eller under, verkligen inträffar, varom han talade med dig, i det att han sade: »Låt oss efterfölja och tjäna andra gudar, som I icke kännen»,
så skall du ändå icke höra på den profetens ord eller på den drömmaren, ty HERREN, eder Gud, sätter eder därmed allenast på prov, för att förnimma om I älsken HERREN, eder Gud, av allt edert hjärta och av all eder själ.
HERREN, eder Gud, skolen I efterfölja, honom skolen I frukta, hans bud skolen I hålla, hans röst skolen I höra, honom skolen I tjäna, och till honom skolen I hålla eder.
Men den profeten eller drömmaren skall dödas, ty han predikade avfall från HERREN, eder Gud, som har fört eder ut ur Egyptens land och förlossat dig ur träldomshuset; och han ville förföra dig till att övergiva den väg som HERREN, din Gud, har bjudit dig att vandra.
Du skall skaffa bort ifrån dig vad ont är.
Om din broder, din moders son, eller din son eller din dotter, eller hustrun i din famn, eller din vän som är för dig såsom ditt eget liv, om någon av dessa i hemlighet vill förleda dig, i det han säger: »Låt oss gå åstad och tjäna andra gudar, som varken du eller dina fäder hava känt»
-- gudar hos de folk som bo runt omkring eder, nära dig eller fjärran ifrån dig, från jordens ena ända till den andra --
så skall du icke göra honom till viljes eller höra på honom.
Du skall icke visa honom någon skonsamhet eller hava misskund och undseende med honom,
utan du skall dräpa honom: först skall din egen hand lyftas mot honom för att döda honom, och sedan hela folkets hand.
Och du skall stena honom till döds, därför att han sökte förföra dig till att övergiva HERREN, din Gud, som har fört dig ut ur Egyptens land, ur träldomshuset.
Och hela Israel skall höra detta och frukta, och man skall sedan icke mer göra något sådant ont bland dig.
Om du får höra att man i någon av de städer, som HERREN vill giva dig till att bo i, berättar
att män hava uppstått bland dig, onda män som förföra invånarna i sin stad, i det att de säga: »Låt oss gå åstad och tjäna andra gudar, som I icke kännen»,
så skall du noga undersöka och rannsaka och efterforska; om det då befinnes vara sant och visst att en sådan styggelse har blivit förövad bland dig,
så skall du slå den stadens invånare med svärdsegg; du skall giva den och allt vad däri är till spillo; också boskapen där skall du slå med svärdsegg.
Och allt byte du får där skall du samla ihop mitt på torget, och därefter skall du bränna upp staden i eld, med allt byte du får där, såsom ett heloffer åt HERREN, din Gud; den skall bliva en grushög för evärdlig tid, aldrig mer skall den byggas upp.
Låt intet av det tillspillogivna låda vi din hand, på det att HERREN må vända sig ifrån sin vredes glöd och låta barmhärtighet vederfaras dig och förbarma sig över dig och föröka dig, såsom han med ed har lovat dina fäder att göra,
om du nämligen hör HERRENS, din Guds, röst, så att du håller alla hans bud, som jag i dag giver dig, och gör vad rätt är i HERRENS, din Guds, ögon.
I ären Herrens, eder Guds, barn.
I skolen icke rista några märken på eder eller göra eder skalliga ovanför pannan för någon död;
ty du är ett folk som är helgat åt Herren, din Gud, och dig har Herren utvalt till att vara hans egendomsfolk framför alla andra folk på jorden.
Du skall icke äta något som är en styggelse.
Dessa äro de fyrfotadjur som I fån äta: fäkreatur, får och getter, hjort,
gasell, dovhjort, stenbock, dison, teoantilop och semer,
alla de fyrfotadjur som hava klövar och hava dem helkluvna i två hälfter, och som idissla; sådana fyrfotadjur fån I äta.
Men dessa skolen I icke äta av de idisslande djuren och av dem som hava genomkluvna klövar: kamelen, haren och klippdassen, ty de idissla väl, men de hava icke klövar, de skola gälla för eder som orena;
svinet, ty det har väl klövar, men det idisslar icke, det skall gälla för eder såsom orent.
Av dessa djurs kött skolen I icke äta, ej heller skolen I komma vid deras döda kroppar.
Detta är vad I fån äta av allt det som lever i vattnet: allt det som har fenor och fjäll fån I äta.
Men intet som icke har fenor och fjäll skolen I äta; det skall gälla för eder så som orent.
Alla rena fåglar fån I äta.
Men dessa fåglar skolen I icke äta: örnen, lammgamen, havsörnen,
raafågeln, falken, gladan med dess arter,
alla slags korpar efter deras arter,
strutsen tahemasfågeln, fiskmåsen, höken med dess arter,
ugglan, uven tinsemetfågeln,
pelikanen, asgamen, dykfågeln,
hägern, regnpiparen med dess arter, härfågeln och flädermusen.
Alla flygande smådjur skola ock gälla för eder såsom orena, de skola icke ätas.
Men alla rena flygande djur fån I äta.
I skolen icke äta något självdött; åt främlingen som bo inom dina portar må du giva sådant, och han må äta det; eller ock må du sälja det åt en utlänning.
Ty du är ett folk som är helgat HERREN, din Gud.
Du skall icke koka en killing i dess moders mjölk.
Tionde skall du giva av all sädesgröda som för vart år växer på din åker,
och du skall äta den inför Herrens, din Guds, ansikte, på den plats som han utväljer till boning åt sitt namn: tionden av din säd, ditt vin och din olja, så ock din förstfödda av dina fäkreatur och din småboskap; ty du skall lära att frukta Herren, din Gud, alltid.
Men om vägen är dig för lång, så att du icke förmår föra det dit, eftersom den plats som Herren, din Gud, utväljer till att där fästa sitt namn ligger för avlägset för dig -- då nu Herren, din Gud, välsigna dig --
så må du sälja det och knyta in penningarna och taga dem med dig och gå till den plats som Herren, din Gud, utväljer.
Och du må köpa för penningarna vadhelst dig lyster fäkreatur eller småboskap, eller vin eller andra starka drycker eller vad du eljest kan åstunda; och så skall du hålla måltid där inför HERRENS, din Guds, ansikte och glädja dig med ditt husfolk.
Och leviten som bor inom dina portar skall du då icke glömma bort, ty han har ingen lott eller arvedel jämte dig.
Vid slutet av vart tredje år skall du avskilja all tionde av vad du har fått i avkastning under det året och lägga upp det inom dina städer.
Och sedan skall leviten få komma, han som ingen lott eller arvedel har jämte dig, så ock främlingen och den faderlöse och änkan som bo inom dina portar; och då skola äta och bliva mätta.
Så skall du göra, för att Herren din Gud, må välsigna dig i alla dina händers verk, i allt vad du gör.
Vart sjunde år skall du låta vara ett friår.
Och så skall förhålla sig med det friåret: Var långivare som har lånat något åt sin nästa skall då efterskänka sin fordran.
Han får då icke kräva sin nästa och broder, ty ett HERRENS friår har då blivit utlyst.
En utlänning må du kräva, men om du har något att fordra av din broder, skall du efterskänka det.
Dock borde rätteligen ingen fattig finnas hos dig, ty Herren skall rikligen välsigna dig i det land som HERREN, din Gud, vill giva dig till besittning, såsom din arvedel,
allenast du hör HERRENS, din Guds, röst, så att du håller alla dessa bud som jag i dag giver dig och gör efter dem.
Ty Herren, din Gud, skall välsigna dig, såsom han har lovat dig; och du skall giva lån åt många folk, men själv skall du icke behöva låna av någon, och du skall råda över många folk, men de skola icke råda över dig.
Om någon fattig finnes hos dig, en av dina bröder inom någon av dina städer, i det land som Herren, din Gud, vill giva dig, så skall du icke förstocka ditt hjärta och tillsluta din hand för denne din fattige broder,
utan du skall gärna öppna din hand för honom och gärna låna honom vad han behöver i sin brist.
Tag dig till vara, så att icke den onda tanken uppstår i ditt hjärta: »Det sjunde året, friåret, är nära», och att du så ser med ont öga på din fattige broder och icke giver honom något; han kan då ropa över dig till Herren, och så kommer synd att vila på dig.
Gärna skall du giva åt honom, och ditt hjärta skall icke vara motvilligt, när du giver åt honom, ty för en sådan gåvas skull skall Herren, din Gud, välsigna dig i alla dina verk, i allt vad du företager dig.
Fattiga skola ju aldrig saknas i landet, därför bjuder jag dig och säger: Du skall gärna öppna din hand för din broder, för de arma och fattiga som du har i ditt land.
Om någon av ditt folk, en hebreisk man eller en hebreisk kvinna, har sålt sig till dig och tjänat dig i sex år, så skall du på det sjunde året släppa honom fri ur din tjänst;
och när du släpper honom fri ur din tjänst, skall du icke låta honom gå med tomma händer.
Du skall fastmer förse honom med gåvor från din hjord, från din loge och från din vinpress; av det varmed Herren, din Gud, har välsignat dig skall du giva honom.
Du skall komma ihåg att du själv har varit en träl i Egyptens land, och att Herren, din Gud, har förlossat dig; därför bjuder jag dig detta i dag.
Men om så skulle hända, att han säger till dig att han icke vill lämna dig, därför att han älskar dig och ditt hus, eftersom han har haft det gott hos dig,
så skall du taga en syl och sticka den genom hans öra in i dörren; därefter skall han vara din träl evärdligen.
Med din tjänarinna skall du göra på samma sätt.
Du skall icke tycka det vara hårt att du måste släppa din tjänare fri ur din tjänst; i sex år har han ju berett dig dubbelt så stor förmån som någon avlönad legodräng.
Så skall Herren, din Gud, välsigna dig i allt vad du gör.
Allt förstfött av hankön, som födes bland dina fäkreatur och din småboskap, skall du helga åt Herren, din Gud; du skall icke vid ditt arbete begagna det som är förstfött bland dina fäkreatur, icke heller skall du klippa ullen på det som är förstfött bland din småboskap.
Inför Herrens, din Guds, ansikte skall du med ditt husfolk för vart år äta det på den plats som Herren utväljer.
Men om djuret har något lyte, om det är halt eller blint eller har något annat ont lyte, så skall du icke offra det åt Herren, din Gud.
Inom dina städer må du då äta det; både den som är oren och den som är ren må äta därav, såsom vore det gasell- eller hjortkött.
Men blodet skall du icke förtära; du skall gjuta ut det på jorden såsom vatten.
Tag i akt månaden Abib och håll Herrens, din Guds, påskhögtid; ty i månaden Abib förde Herren, din Gud, dig ut ur Egypten om natten.
Du skall då slakta påskoffer åt Herren. din Gud, av småboskap och fäkreatur, på den plats som Herren utväljer till boning åt sitt namn.
Du skall icke äta något syrat därtill; i sju dagar skall du äta osyrat bröd därtill, betryckets bröd.
Ty med hast måste du draga ut ur Egyptens land.
I alla dina livsdagar må du därför komma ihåg den dag då du drog ut ur Egyptens land.
I sju dagar må man icke se någon surdeg hos dig, i hela ditt land; och av det som du slaktar om aftonen på den första dagen skall intet kött lämnas kvar över natten till morgonen.
Du får icke slakta påskoffret inom vilken som helst av de städer som Herren, din Gud, vill giva dig,
utan du skall gå till den plats som Herren, din Gud, utväljer till boning åt sitt namn, och där skall du slakta påskoffret om aftonen, när solen går ned den tid på dagen, då den drog ut ur Egypten.
Och du skall koka det och äta det på den plats som Herren, din Gud, utväljer; sedan må du om morgonen vända tillbaka och gå hem till dina hyddor.
I sex dagar skall du äta osyrat bröd, och på sjunde dagen är Herrens, din Guds, högtidsförsamling; då skall du icke göra något arbete.
Sju veckor skall du räkna åt dig; från den dag då man begynner skära säden skall du räkna sju veckor.
Därefter skall du hålla Herrens, din Guds, veckohögtid och bära fram din hands frivilliga gåva, som du må giva efter råd och lägenhet, alltefter måttet av den välsignelse som Herren, din Gud, har givit dig.
Och inför Herrens, din Guds, ansikte skall du glädja dig på den plats som Herren, din Gud, utväljer till boning åt sitt namn, du själv med din son och din dotter, din tjänare och tjänarinna, och med leviten som bor inom dina portar, och främlingen, den faderlöse och änkan som du har hos dig.
Och du skall komma ihåg att du själv har varit en träl i Egypten, och så hålla dessa stadgar och göra efter dem.
Lövhyddohögtiden skall du hålla, i sju dagar, när du inbärgar avkastningen av din loge och av din vinpress.
Och du skall glädja dig vid denna din högtid, med din son och din dotter, din tjänare och din tjänarinna, med leviten, med främlingen, den faderlöse och änkan som bo inom dina portar.
I sju dagar skall du hålla Herrens, din Guds, högtid, på den plats som Herren utväljer; ty Herren, din Gud, skall välsigna dig i all den avkastning du får och i dina händers alla verk, och du skall vara uppfylld av glädje.
Tre gånger om året skall allt ditt mankön träda fram inför Herrens, din Guds, ansikte, på den plats som han utväljer: vid det osyrade brödets högtid, vid veckohögtiden och vid lövhyddohögtiden.
Men med tomma händer skall ingen träda fram inför Herrens ansikte,
utan var och en skall: giva vad hans hand förmår, alltefter måttet av den välsignelse som Herren, din Gud, har givit dig.
Domare och tillsyningsmän skall du tillsätta åt dig inom alla de städer som Herren, din Gud, vill giva dig, för dina särskilda stammar; de skola döma folket med rättvis dom.
Du skall icke vränga rätten och icke hava anseende till personen; och du skall icke taga mutor, ty mutor förblinda de visas ögon och förvrida de rättfärdigas sak.
Rättfärdighet, rättfärdighet skall du eftertrakta, för att du må leva och taga i besittning det land som Herren, din Gud, vill giva dig.
Du skall icke plantera åt dig Aseror av något slags träd, vid sidan av Herrens, din Guds, altare, det som du skall göra åt dig;
icke heller skall du resa åt dig någon stod, ty sådant hatar Herren, din Gud.
Du skall icke offra åt Herren, din Gud, något djur av fäkreaturen eller av småboskapen, som har något lyte eller något annat fel, ty sådant är en styggelse för Herren, din Gud.
Om bland dig, inom någon av de städer som Herren, din Gud, vill giva dig, någon man eller kvinna befinnes göra vad ont är i Herrens, din Guds, ögon, i det att han överträder hans förbund,
och går åstad och tjänar andra gudar och tillbeder dem, eller ock solen eller månen eller himmelens hela härskara, mot mitt bud,
och detta bliver berättat för dig, så att du får höra därom, då skall du noga undersöka saken; om det då befinnes vara sant och visst att en sådan styggelse har blivit förövad i Israel,
så skall du föra den man eller den kvinna som har gjort denna onda gärning ut till din stadsport det må nu vara en man eller en kvinna-och stena den skyldige till döds.
Efter två eller tre vittnens utsago skall han dödas; ingen skall dömas till döden efter allenast ett vittnes utsago.
Först skall vittnenas hand lyftas mot honom för att döda honom, och sedan hela folkets hand: du skall skaffa bort ifrån dig vad ont är.
Om det i något fall bliver dig för svårt att själv döma i en blodssak eller i en rättsfråga eller i ett misshandlingsmål eller överhuvud i någon sak varom man tvistar i dina portar, så skall du-stå upp och begiva dig till den plats som HERREN, din Gud, utväljer,
och gå till de levitiska prästerna, och till den som på den tiden är domare; dem skall du fråga, och de skola förkunna för dig vad som är rätt.
Och i enlighet med vad de förkunna för dig där, på den plats som Herren utväljer. skall du göra; du skall i alla stycken hålla och göra vad de lära dig.
Efter den lag som de lära dig, och efter den dom som de avkunna för dig skall du göra.
Från det som de förkunna för dig skall du icke vika av, vare sig till höger eller till vänster.
Men om någon gör sig skyldig till den förmätenheten att icke vilja lyssna till prästen, som står och gör tjänst där inför Herren, din Gud, eller till domaren, så skall den mannen dö: du skall skaffa bort ifrån Israel vad ont är.
Och allt folket skall höra det och frukta, och de skola icke mer göra sig skyldiga till sådan förmätenhet.
När du kommer in i det land som Herren, din Gud, vill giva dig, och du tager det i besittning och bor där om du då säger: »Jag vill sätta en konung över mig, såsom alla folk omkring mig hava»,
så skall du till konung över dig sätta den som Herren, din Gud, utväljer.
En av dina bröder skall du sätta till konung över dig; du får icke sätta till konung över dig en utländsk man, som icke är din broder.
Men han må icke skaffa sig hästar i mängd, och icke sända sitt folk tillbaka till Egypten för att skaffa de många hästarna, ty Herren har ju sagt till eder: »I skolen icke mer återvända denna väg.»
Icke heller skall han skaffa sig hustrur i mängd, på det att hans hjärta icke må bliva avfälligt; och icke heller skall han skaffa sig alltför mycket silver och guld.
Och när han har blivit uppsatt på sin konungatron, skall han hämta denna lag från de levitiska prästerna och taga en avskrift därav åt sig i en bok.
Och den skall han hava hos sig och läsa i den i alla sina livsdagar, för att han må lära att frukta Herren, sin Gud, så att han håller alla denna lags ord och dessa stadgar och gör efter dem.
Så skall han göra, för att hans hjärta icke må förhäva sig över hans bröder, och för att han icke må vika av ifrån buden, vare sig till höger eller till vänster; på det att han och hans söner må länge regera; sitt rike, bland Israels folk.
De levitiska prästerna, hela Levi stam, skola ingen lott eller arvedel hava med det övriga Israel; av HERRENS eldsoffer och hans arvedel skola de hava sitt underhåll.
De skola icke hava någon arvedel bland sina bröder; Herren är deras arvedel, såsom han har sagt dem.
Och detta skall vara vad prästerna hava rätt att få av folket, av dem som offra ett slaktoffer, vare sig av fäkreaturen eller av småboskapen: man skall giva prästen bogen, käkstyckena och vommen.
Förstlingen av din säd, ditt vin och din olja, och förstlingen av dina fårs ull skall du giva honom.
Ty honom har Herren, din Gud, utvalt bland alla dina stammar, för att han och hans söner alltid skola stå och göra tjänst i Herrens namn.
Och om leviten vill komma från någon av dina städer, inom vilken han vistas någonstädes i Israel, så må det stå honom fritt att komma, såsom honom lyster, till den plats som Herren utväljer,
och han må då göra tjänst i HERRENS, sin Guds, namn, likasom alla hans bröder, leviterna, som stå där inför HERRENS ansikte.
De skola alla hava lika mycket till sitt underhåll, oberäknat vad någon kan äga genom försäljning av sitt fädernearv.
När du kommer in i det land som HERREN, din Gud, vill giva dig, skall du icke lära dig att göra efter hedningarnas styggelser.
Hos dig må icke finnas någon som låter sin son eller dotter gå genom eld, eller som befattar sig med trolldom eller teckentydning eller svartkonst eller häxeri,
ingen som förehar besvärjelsekonster, ingen som frågar andar, eller som är en spåman, eller som söker råd hos de döda.
Ty en styggelse för Herren är var och en som gör sådant, och för sådana styggelsers skull fördriver HERREN, din Gud, dem för dig.
Du skall vara ostrafflig inför HERREN, din Gud.
Hedningarna som du nu fördriver lyssna väl till sådana som öva teckentydning och trolldom, men dig har HERREN, din Gud, icke tillstatt sådant.
En profet bland ditt folk, av dina bröder, en som är mig lik, skall HERREN, din Gud, låta uppstå åt dig; honom skolen I lyssna till.
Det skall bliva alldeles såsom du begärde av HERREN, din Gud, vid Horeb, den dag då I voren där församlade och du sade: »Låt mig icke vidare höra HERRENS, min Guds, röst, och låt mig slippa att längre se denna stora eld, på det att jag icke må dö.»
Och HERREN sade till mig: »De hava rätt i vad de hava talat.
En profet skall jag låta uppstå åt dem bland deras bröder, en som är dig lik, och jag skall lägga mina ord i hans mun, och han skall tala till dem allt vad jag bjuder honom.
Och om någon icke lyssnar till mina ord, de ord han talar i mitt namn, så skall jag själv utkräva det av honom.
Men den profet som är så förmäten, att han i mitt namn talar vad jag icke har bjudit honom tala, eller som talar i andra gudars namn, den profeten skall dö.
Och om du säger vid dig själv: 'Huru skola vi känna igen det som icke är talat av HERREN?',
så må du veta: när profeten talar i HERRENS namn, och det som han har talat icke sker och icke inträffar, då är detta något som HERREN icke har talat; i förmätenhet har då profeten talat det; du skall icke frukta för honom.»
När HERREN, din Gud, har utrotat de folk vilkas land HERREN, din Gud, vill giva dig, och när du har fördrivit dem och bosatt dig i deras städer och i deras hus,
då skall du avskilja åt dig tre städer i ditt land, det som HERREN, din Gud, vill giva dig till besittning.
Du skall försätta vägarna till dem i gott skick åt dig; och du skall dela i tre delar det landområde som HERREN, din Gud, giver dig till arvedel.
Så skall du göra, för att var och en som har dräpt någon må kunna fly dit.
Och under följande villkor må en dråpare fly till någon av dem och så bliva vid liv; om någon dödar sin nästa utan vett och vilja, och utan att förut hava burit hat till honom
-- såsom när någon går med sin nästa ut i skogen för att hugga ved, och hans hand hugger till med yxan för att fälla trädet, och järnet då far av skaftet och träffar den andre, så att denne dör -- då må en sådan fly till någon av dessa städer och så bliva vid liv.
Detta vare stadgat, för att blodshämnaren, om han i sitt hjärtas vrede förföljer dråparen, icke må hinna upp honom, ifall vägen är för lång, och slå ihjäl honom, fastän han icke hade förtjänat döden, eftersom han icke förut hade burit hat till den andre.
Därför är det som jag bjuder dig och säger: »Tre städer skall du avskilja åt dig.»
Och när HERREN, din Gud, utvidgar ditt område, såsom han med ed har lovat dina fäder, och giver dig allt det land som han har sagt att han skulle giva åt dina fäder --
om du då håller och gör efter alla dessa bud som jag i dag giver dig, så att du älskar HERREN, din Gud, och alltid vandrar på hans vägar, då skall du lägga ännu tre städer till dessa tre,
för att oskyldigt blod icke må utgjutas i ditt land, det som HERREN, din Gud, vill giva dig till arvedel, och blodskuld så komma att vila på dig.
Men om någon bär hat till sin nästa och lägger sig i försåt för honom och överfaller honom och slår honom till döds, och sedan flyr till någon av dessa städer,
då skola de äldste i hans stad sända bort och hämta honom därifrån och lämna honom i blodshämnarens hand, och han skall dö.
Du skall icke visa honom någon skonsamhet, utan du skall skaffa bort ifrån Israel skulden för den oskyldiges blod, för att det må gå dig väl.
Du skall icke flytta din nästas råmärke, något råmärke som förfäderna hava satt upp i den arvedel du får i det land som HERREN, din Gud, vill giva dig till besittning.
Det är icke nog att allenast ett vittne träder upp mot någon angående någon missgärning eller synd, vad det nu må vara för en synd som någon kan hava begått.
Efter två eller efter tre vittnens utsago skall var sak avgöras.
Om ett orättfärdigt vittne träder upp mot någon för att vittna mot honom angående någon förbrytelse,
så skola båda parterna träda fram inför HERRENS ansikte, inför de män som på den tiden äro präster och domare.
Och domarna skola noga undersöka saken; om då vittnet befinnes vara ett falskt vittne, som har burit falskt vittnesbörd mot sin broder,
så skolen I låta detsamma vederfaras honom som han hade tilltänkt sin broder: du skall skaffa bort ifrån dig vad ont är.
Och det övriga folket skall höra det och frukta, och man skall icke vidare göra något sådant ont bland eder.
Du skall icke visa honom någon skonsamhet: liv för liv, öga for öga, tand för tand, hand för hand, fot för fot.
Om du drager ut i krig mot dina fiender, och du då får se hästar och vagnar och ett folk som är större än du. så skall du dock icke frukta för dem, ty HERREN, din Gud, är med dig, han som har fört dig upp ur Egyptens land.
När I då stån färdiga att gå i striden, skall prästen träda fram och tala till folket;
han skall säga till dem: »Hör, Israel!
I stån nu färdiga att gå i strid mot edra fiender.
Edra hjärtan vare icke försagda; frukten icke och ängslens icke, och varen icke förskräckta för dem,
ty HERREN, eder Gud, går själv med eder; till att strida för eder mot edra fiender och giva eder seger.»
Och tillsyningsmännen skola tala till folket och säga: »Om någon finnes här, som har byggt sig ett nytt hus, men ännu icke invigt det, så må han vända tillbaka hem, för att icke. om han faller i striden, en annan må komma att inviga det.
Och om någon finnes här, som har planterat en vingård, men ännu icke fått skörda någon frukt därav, så må han vända tillbaka hem, för att icke, om han faller i striden, en annan må komma att hämta första skörden av den.
Och om någon finnes här, som har trolovat sig med en kvinna, men ännu icke tagit henne till sig, så må han vända tillbaka hem, för att icke om han faller i striden, en annan man må taga henne till sig.»
Vidare skola tillsyningsmännen tala till folket och säga: »Om någon finnes här, som fruktar och har ett försagt hjärta, så må han vända tillbaka hem, för att icke också hans bröders hjärtan må bliva uppfyllda av räddhåga, såsom hans eget hjärta är.»
Och när tillsyningsmännen så hava talat till folket, skola hövitsmän tillsättas övar härens avdelningar, till att gå i spetsen för folket.
När du kommer till någon stad för att belägra den, skall du först tillbjuda den fred.
Om den då giver dig ett fridsamt svar och öppnar sina portar för dig, så skall allt folket som finnes där bliva arbetspliktigt åt dig och vara dina tjänare.
Men om den icke vill hava fred med dig, utan vill föra krig mot dig, så må du belägra den.
Och om HERREN, din Gud, då giver den i din hand, skall du slå allt mankön där med svärdsegg.
Men kvinnorna och barnen och boskapen och allt annat som finnes i staden, allt rov du får där, skall du hava såsom ditt byte; och du må då njuta av det rov som HERREN. din Gud, låter dig taga från dina fiender.
Så skall du göra med alla de städer som äro mer avlägsna från dig, och som icke höra till dessa folks städer.
Men i de städer som tillhöra dessa folk, och som HERREN, din Gud, vill giva dig till arvedel, skall du icke låta något som anda har bliva vid liv,
utan du skall giva dem alla till spillo: hetiterna och amoréerna, kananéerna och perisséerna, hivéerna och jebuséerna, såsom HERREN din Gud, har bjudit dig.
Så skall du göra, för att de icke må lära eder att bedriva alla de styggelser som de själva hava bedrivit till sina gudars ära, och så komma eder att synda mot HERREN, eder Gud.
Om du måste länge belägra en stad för att erövra och intaga den, så skall du icke förstöra träden däromkring genom att höja din yxa mot dem; du må äta av deras frukt, men du skall icke hugga ned dem; träden på marken äro ju icke människor som skola belägras av dig.
Men de träd om vilka du vet att de icke bära ätbar frukt, dem må du förstöra och hugga ned för att av dem bygga bålverk mot den fientliga staden, till dess att den faller
Om i det land som HERREN, din Gud, vill giva dig till besittning en ihjälslagen människa påträffas liggande på marken, och man icke vet vem som har dödat honom,
så skola dina äldste och dina domare gå ut och mäta upp avståndet från platsen där den ihjälslagne påträffas till de städer som ligga där runt omkring.
Och de äldste i den stad som ligger närmast denna plats skola taga en kviga som icke har blivit begagnad till arbete, och som icke såsom dragare har gått under ok.
Och de äldste i staden skola föra kvigan ned till en dalgång som icke har varit plöjd eller besådd; och där i dalen skola de krossa nacken på kvigan.
Och prästerna, Levi söner, skola träda fram, ty dem har HERREN, din Gud, utvalt till att göra tjänst inför honom och till att välsigna i HERRENS namn, och såsom de bestämma skola alla tvister och alla misshandlingsmål behandlas.
Och alla de äldste i den staden, de som bo närmast platsen där den ihjälslagne påträffades, skola två sina händer över kvigan på vilken man hade krossat nacken i dalen;
och de skola betyga och säga: »Våra händer hava icke utgjutit detta blod, och våra ögon hava icke sett dådet.
Förlåt ditt folk Israel, som du har förlossat, HERRE, och låt icke oskyldigt blod komma över någon i ditt folk Israel.»
Så bliver denna blodskuld dem förlåten.
Du skall skaffa bort ifrån dig skulden för det oskyldiga blodet, ty du skall göra vad rätt är i HERRENS ögon.
Om HERREN, din Gud, när du drager ut i krig mot dina fiender, giver dem i din hand, så att du tager fångar,
och du då bland fångarna får se någon skön kvinna som du fäster dig vid, och som du vill taga till hustru åt dig,
så skall du föra henne in i ditt hus, och hon skall raka sitt huvud och ansa sina naglar.
Och hon skall lägga av de kläder hon bar såsom fånge och skall bo i ditt hus och få begråta sin fader och sin moder en månads tid; därefter må du gå in till henne och äkta henne, så att hon bliver din hustru.
Och om du sedan icke mer finner behag i henne, så må du låta henne gå vart hon vill; du får icke sälja henne för penningar.
Du får icke heller behandla henne såsom trälinna, då du nu har kränkt henne.
Om en man har två hustrur, en som han älskar och en som han försmår, och båda hava fött honom söner, såväl den han älskar som den han försmår, och hans förstfödde son till den försmådda,
så får mannen icke, när han åt sina söner utskiftar sin egendom såsom arv, giva förstfödslorätten åt sonen till den älskar, till förfång för sonen till den han försmår, då nu denne är den förstfödde,
utan han skall såsom sin förstfödde erkänna sonen till den försmådda och giva honom dubbel lott av allt vad han äger.
Ty denne är förstlingen av hans kraft; honom tillhör förstfödslorätten.
Om någon har en vanartig och uppstudsig son, som icke lyssnar till sin faders och sin moders ord, och som, fastän de tukta honom, ändå icke hör på dem,
så skola hans fader och hans moder taga honom och föra honom ut till de äldste i staden, till stadens port.
Och de skola säga till de äldste i staden: »Denne vår son är vanartig och uppstudsig och vill icke lyssna till våra ord, utan är en frossare och drinkare.»
Då skall allt folket i staden stena honom till döds: du skall skaffa bort ifrån dig vad ont är.
Och hela Israel skall höra det och frukta.
Om på någon vilar en sådan synd som förtjänar döden, och han så bliver dödad och du hänger upp honom på trä,
så skall den döda kroppen icke lämnas kvar på träet över natten, utan du skall begrava den på samma dag, ty en Guds förbannelse är den som har blivit upphängd; och du skall icke orena det land som HERREN, din Gud, vill giva dig till arvedel.
Om du ser din broders oxe eller får gå vilse, skall du icke undandraga dig att taga vara på djuret; du skall föra det tillbaka till din broder.
Och om din broder icke bor i din närhet, eller om du icke vet vem det är, så skall du taga djuret in i ditt hus, och det skall vara hos dig, till dess din broder frågar efter det; då skall du lämna det tillbaka åt honom.
På samma sätt skall du göra med hans åsna, på samma sätt med hans kläder, och på samma sätt skall du göra med allt annat som din broder kan hava förlorat, och som du hittar; du får icke draga dig undan.
Om du ser din broders åsna eller oxe falla på vägen, skall du icke undandraga dig att bistå djuret; du skall hjälpa honom att resa upp det.
En kvinna skall icke bära vad till en man hör, ej heller skall en man sätta på sig kvinnokläder; ty var och en som så gör är en styggelse för HERREN, din Gud.
Om du på din väg träffar på ett fågelbo, i något träd eller på marken, med ungar eller ägg i, och modern ligger på ungarna eller på äggen, så skall du icke taga både modern och ungarna.
Du skall låta modern flyga och taga allenast ungarna; så skall du göra, för att det må gå dig väl och du må länge leva.
När du bygger ett nytt hus, skall du förse taket med bröstvärn, för att du icke må draga blodskuld över ditt hus, om någon faller ned därifrån.
Du skall icke, för att få två slags skörd i din vingård, så säd däri, på det att icke alltsammans, både vad du har sått och vad själva vingården avkastar, må hemfalla till helgedomen.
Du skall icke plöja med oxe och åsna tillsammans.
Du skall icke kläda dig i tyg av olika garn, av ull och lin tillsammans.
Du skall göra dig tofsar i de fyra hörnen på överklädnaden som du höljer dig i.
Om en man har tagit sig en hustru och gått in till henne, men sedan får motvilja mot henne,
och då påbördar henne skamliga ting och sprider ut ont rykte om henne och säger: »Denna kvinna tog jag till hustru; men när jag låg hos henne, fann jag icke tecknen till att hon var jungfru»,
så skola flickans fader och moder taga tecknen till att flickan var jungfru och bära dem ut till de äldste i staden, där de sitta i porten.
Och flickans fader skall säga till de äldste: »Jag gav min dotter till hustru åt denne man, men han har fått motvilja mot henne.
Och nu påbördar han henne skamliga ting och säger: 'Jag har icke funnit tecknen till att din dotter var jungfru'; men här äro tecknen till att min dotter var jungfru.»
Och de skola breda ut klädet inför de äldste i staden.
Då skola de äldste i staden taga mannen och tukta honom.
Och de skola ålägga honom att böta hundra siklar silver, vilka han skall giva åt flickans fader, därför att han har spritt ut ont rykte om en jungfru i Israel.
Och hon skall vara hans hustru, och han får icke skilja sig från henne, så länge han lever.
Men om det var sanning, om tecknen till att flickan var jungfru icke funnos,
då skall man föra ut flickan utanför dörren till hennes faders hus, och männen i staden skola stena henne till döds därför att hon har gjort vad som var en galenskap i Israel, då hon bedrev otukt i sin faders hus: du skall skaffa bort ifrån dig vad ont är.
Om en man ertappas med att ligga hos en kvinna som är en annan mans äkta hustru, så skola båda dö, både mannen som låg hos kvinnan, och jämväl kvinnan: du skall skaffa bort ifrån Israel vad ont är.
Om en jungfru är trolovad med en man, och en annan man träffar henne i staden och lägrar henne,
så skolen I föra dem båda ut till stadens port och stena dem till döds, flickan, därför att hon icke ropade på hjälp i staden, och mannen, därför att han kränkte en annans trolovade: du skall skaffa bort ifrån dig vad ont är.
Men om det var ute på marken som mannen träffade den trolovade flickan, och han där tog henne med våld och lägrade henne, så skall mannen som lägrade henne ensam dö.
Men flickan skall du icke göra något, flickan har icke begått någon synd som förtjänar döden; utan det är med denna sak, såsom när en man överfaller en annan och dräper honom.
Ty då det var ute på marken som han träffade den trolovade flickan, kan hon hava ropat, utan att någon fanns där, som kunde frälsa henne.
Om däremot en man träffar en jungfru som icke är trolovad, och han tager fatt henne och lägrar henne, och de ertappas,
så skall mannen som lägrade flickan giva åt flickans fader femtio siklar silver och taga henne själv till sin hustru, därför att han har kränkt henne; han får icke skilja sig från henne, så länge han lever.
Ingen skall taga sin faders hustru och lyfta på sin faders täcke.
Ingen som är snöpt, vare sig genom krossning eller genom stympning, skall komma in i HERRENS församling.
Ingen som är född i äktenskapsbrott eller blodskam skall komma in i HERRENS församling; icke ens den som i tionde led är avkomling av en sådan skall komma in i HERRENS församling.
Ingen ammonit eller moabit skall komma in i HERRENS församling; icke ens den som i tionde led är avkomling av en sådan skall någonsin komma in i HERRENS församling --
detta därför att de icke kommo eder till mötes med mat och dryck på vägen, när I drogen ut ur Egypten, och därför att han mot dig lejde, Bileam, Beors son, från Petor i Aram-Naharaim, för att denne skulle förbanna dig.
Men HERREN, din Gud, ville icke höra på Bileam, utan HERREN, din Gud, förvandlade förbannelsen till välsignelse för dig, ty HERREN, din Gud, älskade dig.
Du skall aldrig, i all din tid, fråga efter deras välfärd och lycka.
Edoméen skall däremot icke för dig vara en styggelse, ty han är din broder.
Egyptiern skall icke heller för dig vara en styggelse, ty i hans land har du bott såsom främling.
Barn som födas av dessa i tredje led må komma in i HERRENS församling.
När du drager ut mot dina fiender och slår läger, skall du taga, dig till vara för allt vad orent är.
Om bland dig finnes någon som icke är ren, därigenom att något har hänt honom under natten, så skall han gå ut till något ställe utanför lägret; han får icke komma in i lägret.
Och mot aftonen skall han bada sig i vatten, och när solen går ned, får han gå in i lägret. --
Du skall hava en särskild plats utanför lägret, dit du kan gå avsides.
Och du skall jämte annat som du bär hava en pinne, och när du vill sätta dig därute, skall du med den gräva en grop och sedan åter täcka över din uttömning.
Ty HERREN, din Gud, vandrar fram i ditt läger för att hjälpa dig och giva dina fiender i ditt våld; därför skall ditt läger vara heligt, så att han icke hos dig ser något som väcker hans leda och fördenskull vänder sig bort ifrån dig.
En träl som har flytt till dig från sin herre skall du icke utlämna till hans herre.
Han skall få stanna hos dig, mitt ibland dig, på det ställe som han utväljer inom någon av dina städer, var han finner för gott; och du skall icke förtrycka honom.
Ingen tempeltärna skall finnas bland Israels döttrar, och ingen tempelbolare bland Israels söner.
Du skall icke bära skökolön och hundpenningar in i HERRENS, din Guds, hus, till gäldande av något löfte; ty det ena som det andra är en styggelse för HERREN, din Gud.
Du skall icke taga ränta av din broder, varken på penningar eller på livsmedel eller på något annat varpå ränta kan tagas.
Av utlänningen må du taga ränta, men icke av din broder, på det att HERREN, din Gud, i allt vad du företager dig, må välsigna dig i det land dit du nu kommer, för att taga det i besittning.
Om du har gjort ett löfte åt HERREN, din Gud, skall du icke dröja att infria det, ty HERREN, din Gud, skall förvisso utkräva det av dig, och synd kommer att vila på dig.
Men om du underlåter att göra något löfte, så kommer icke därigenom synd att vila på dig.
Vad dina läppar hava talat skall du hålla och göra, i enlighet med det frivilliga löfte du har givit HERREN, din Gud, och uttalat med din mun.
När du kommer in i din nästas vingård, får du där äta druvor, så mycket dig lyster, till dess du bliver mätt, men du får icke lägga något i ditt kärl.
När du kommer in på din nästas sädesfält, får du plocka ax med din hand, men med skära får du icke komma vid din nästas säd.
Om en man har tagit sig en hustru och äktat henne, men hon sedan icke längre finner nåd för hans ögon, därför att han hos henne har funnit något som väcker hans leda, och om han fördenskull har skrivit skiljebrev åt henne och givit henne det i handen och skickat bort henne från sitt hus,
och kvinnan sedan, när hon har lämnat hans hus, går åstad och bliver en annans hustru,
och nu också denne andre man får motvilja mot henne och skriver skiljebrev åt henne och giver henne det i handen och skickar henne bort ifrån sitt hus, eller om denne andre man som har tagit henne till sin hustru dör,
då får icke hennes förste man, som skickade bort henne, åter taga henne till sin hustru, sedan hon har låtit orena sig, ty detta vore en styggelse inför HERREN; du skall icke draga synd över det land som HERREN, din Gud, vill giva dig till arvedel.
Om en man nyligen har tagit sig hustru, behöver han icke gå i krigstjänst, ej heller må någon annan tjänstgöring åläggas honom.
Han skall vara fri ett år för att stanna hemma och glädja den hustru han har tagit.
Man skall icke taga handkvarnen eller ens kvarnens översten i pant, ty den så gör tager livet i pant.
Om en man befinnes hava stulit någon av sina bröder, Israels barn, och han behandlar denne såsom träl eller säljer honom, så skall tjuven dö: du skall skaffa bort ifrån dig vad ont är.
Tag dig till vara, så att du, när någon bliver angripen av spetälska, noga håller och gör allt som de levitiska prästerna lära eder.
Vad jag har bjudit dem skolen I hålla och göra.
Kom ihåg vad HERREN, din Gud, gjorde med Mirjam på vägen, när I drogen ut ur Egypten.
Om du giver något lån åt din nästa, så skall du icke gå in i hans hus och taga pant av honom.
Du skall stanna utanför, och mannen som du har lånat åt skall bära ut panten till dig.
Och om det är en fattig man, så skall du icke hava hans pant till täcke, när du ligger och sover.
Du skall giva honom panten tillbaka, när solen går ned, så att han kan hava sin mantel på sig när han ligger och sover, och så välsigna dig; och detta skall lända dig till rättfärdighet inför HERREN, din Gud.
Du skall icke göra en arm och fattig daglönare orätt, evad han är en dina bröder, eller han är en av främlingarna som äro hos dig i ditt land, inom dina portar.
Samma dag han har gjort sitt arbete skall du giva honom hans lön och icke låta solen gå ned däröver, eftersom han är arm och längtar efter sin lön; han kan eljest ropa över dig till HERREN, och så kommer synd att vila på dig.
Föräldrarna skola icke dödas för sina barns skull och barnen skola icke dödas för sina föräldrars skull; var och en skall lida döden genom sin egen synd.
Du skall icke vränga rätten för främlingen eller den faderlöse, och en änkas kläder skall du icke taga i pant;
du skall komma ihåg att du själv har varit en träl i Egypten, och att HERREN, din Gud, har förlossat dig därifrån; därför bjuder jag dig att iakttaga detta.
Om du, när du inbärgar skörden på din åker, glömmer en kärve kvar på åkern, skall du icke gå tillbaka för att hämta den, ty den skall tillhöra främlingen, den faderlöse och änkan.
Detta skall du iakttaga, för att HERREN, din Gud, må välsigna dig i alla dina händers verk.
När du har slagit ned dina oliver, skall du icke sedan genomsöka grenarna; vad där finnes kvar skall tillhöra främlingen den faderlöse och änkan.
När du har avbärgat din vingård, skall du sedan icke göra någon efterskörd; vad där finnes kvar skall tillhöra främlingen, den faderlöse och änkan.
Du skall komma ihåg att du själv har varit en träl i Egyptens land; därför bjuder jag dig att iakttaga detta.
Om en tvist uppstår mellan män, och de komma inför rätta, för att man där skall döma mellan dem, så skall man fria den oskyldige och fälla den skyldige.
Om då den skyldige dömes till hudflängning, skall domaren befalla honom att lägga sig ned, och skall i sin åsyn låta giva honom det antal slag, som svarar emot hans brottslighet.
Fyrtio slag får han giva honom, men icke mer, så att din broder icke bliver vanärad i dina ögon, därigenom att man giver honom oskäligt många slag, flera än som sades.
Du skall icke binda munnen till på oxen som tröskar.
När bröder bo tillsammans, och en av dem dör barnlös, då skall den dödes hustru icke gifta sig med någon främmande man utom släkten; hennes svåger skall gå in till henne och taga henne till hustru, och så äkta henne i sin broders ställe.
Och den förste son hon föder skall upptaga den döde broderns namn, för att dennes namn icke må utplånas ur Israel.
Men om mannen icke vill taga sin svägerska till äkta, så skall svägerskan gå upp i porten, till de äldste, och säga: Min svåger vägrar att upprätthålla sin broders namn i Israel; han vill icke äkta mig i sin broders ställe.»
Då skola de äldste i staden där han bor kalla honom till sig och tala med honom.
Om han då står fast och säger: »Jag vill icke taga henne till äkta»,
så skall hans svägerska träda fram till honom inför de äldstes ögon och draga skon av hans fot och spotta honom i ansiktet och betyga och säga: »Så gör man med den man som icke vill uppbygga sin broders hus.»
Och hans hus skall sedan i Israel heta »den barfotades hus».
Om två män träta med varandra, och den enes hustru kommer för att hjälpa sin man mot den andre, när denne slår honom, och hon därvid räcker ut sin hand och fattar i hans blygd,
så skall du hugga av henne handen, utan att visa henne någon skonsamhet.
Du skall icke hava två slags vikt i din pung, ett större slag och ett mindre,
ej heller skall du i ditt hus hava två slags efa-mått, ett större och ett mindre.
Full och riktig vikt skall du hava, fullmåligt och riktigt efa-mått skall du ock hava, för att du må länge leva i det land som HERREN, din Gud, vill giva dig.
Ty en styggelse för HERREN, din Gud, är var och en som så gör, var och en som gör orätt.
Kom ihåg vad Amalek gjorde mot dig på vägen, när I drogen ut ur Egypten,
huru han, utan att frukta Gud, gick emot dig på vägen och slog din eftertrupp, alla de svaga som hade blivit efter, medan du var trött och utmattad.
Därför, när HERREN, din Gud, har låtit dig få ro för alla dina fiender runt omkring, i det land som HERREN, din Gud, vill giva dig till besittning såsom din arvedel, skall du så utplåna minnet av Amalek, att det icke mer skall finnas under himmelen.
Förgät icke detta.
När du du kommer in i det land som HERREN, din Gud, vill giva dig till arvedel, och du tager det i besittning och bor där,
då skall du taga förstling av all markens frukt, av vad du får i avkastning av landet som HERREN, din Gud, vill giva dig, och lägga detta i en korg och gå därmed till den plats som HERREN, din Gud, utväljer till boning åt sitt namn.
Och du skall gå till den som på den tiden är präst och säga till honom: »Jag förklarar i dag för HERREN, din Gud, att jag har kommit in i det land som HERREN med ed har lovat våra fäder att giva oss.»
Och prästen skall taga korgen ur din hand och sätta den ned inför HERRENS, din Guds, altare.
Och du skall betyga och säga inför HERRENS, din Guds, ansikte: »Min fader var en hemlös aramé, som drog ned till Egypten och bodde där såsom främling med en ringa hop, och där blev av honom ett stort, mäktigt och talrikt folk.
Men sedan behandlade egyptierna oss illa och förtryckte oss och lade hårt arbete på oss.
Då ropade vi till HERREN, våra fäders Gud, och HERREN hörde vår röst och såg vårt lidande och vår vedermöda och vårt betryck.
Och HERREN förde oss ut ur Egypten med stark hand och uträckt arm, med stora och fruktansvärda gärningar, med tecken och under.
Och han lät oss komma hit och gav oss detta land, ett land som flyter av mjölk och honung.
Och här bär jag nu fram förstlingen av frukten på den mark som du, HERRE, har givit mig.»
Och du skall sätta korgen ned inför HERRENS, din Guds, ansikte och tillbedja inför HERRENS, din Guds, ansikte.
Och över allt det goda som HERREN, din Gud har givit åt dig och ditt hus skall du glädja dig, och jämte dig leviten och främlingen som bor hos dig.
När du under det tredje året, tiondeåret, har lagt av all tionde av vad du då har fått i avkastning och givit den åt leviten, främlingen, den faderlöse och änkan, och de hava ätit därav inom dina portar och blivit mätta,
då skall du så säga inför HERRENS, din Guds, ansikte: »Jag har nu fört bort ur mitt hus det heliga, och jag har givit det åt leviten och främlingen, åt den faderlöse och änkan, alldeles såsom du har bjudit mig; jag har icke överträtt eller förgätit något av dina bud.
Jag åt intet därav, när jag hade sorg, och jag förde icke bort något därav, när jag var oren, ej heller använde jag något därav för någon död.
Jag har lyssnat till HERRENS, min Guds, röst; jag har i alla stycken gjort såsom du har bjudit mig.
Skåda nu ned från din heliga boning, himmelen, och välsigna ditt folk Israel och det land som du har givit oss, såsom du med ed lovade våra fäder, ett land som flyter av mjölk och honung.»
I dag bjuder dig HERREN, din Gud, att göra efter dessa stadgar och rätter; du skall hålla dem och göra efter dem av allt ditt hjärta och av all din själ.
Du har i dag hört HERREN förklara att han vill vara din Gud, och att du skall vandra på hans vägar och hålla hans stadgar och bud och rätter och lyssna till hans röst.
Och HERREN har i dag hört dig förklara att du vill vara hans egendomsfolk, såsom han har sagt till dig, och att du vill hålla alla hans bud;
på det att han över alla folk som han har gjort må upphöja dig till lov, berömmelse och ära, och på det att du må vara ett folk som är helgat åt HERREN, din Gud, såsom han har sagt.
Och Mose och de äldste i Israel bjödo folket och sade: »Hållen alla de bud som jag i dag giver eder.
Och när I kommen över Jordan, in i det land som HERREN, din Gud, vill giva dig, då skall du resa åt dig stora stenar och bestryka dem med kalk.
På dessa skall du, när du har gått över floden, skriva alla denna lags ord, för att du må komma in i det land som HERREN, din Gud, vill giva dig, ett land som flyter av mjölk och honung, såsom HERREN, dina fäders Gud, har lovat dig.
Och när I haven gått över Jordan, skolen I på berget Ebal resa dessa stenar om vilka jag i dag giver eder befallning; och du skall bestryka dem med kalk.
Och du skall där åt HERREN, din Gud, bygga ett altare, ett altare av stenar, vid vilka du icke skall komma med något järn.
Av ohuggna stenar skall du bygga HERRENS, din Guds, altare; och du skall på det offra brännoffer åt HERREN, din Gud.
Du skall där ock offra tackoffer och skall äta och glädja dig inför HERRENS, din Guds. ansikte.
Och du skall på stenarna skriva alla denna lags ord, klart och tydligt.»
Och Mose och de levitiska prästerna talade till hela Israel och sade: »Var stilla och hör, Israel!
I dag har du blivit HERRENS, din Guds, folk.
Så skall du då höra HERRENS, din Gud röst och göra efter hans bud och stadgar, som jag i dag giver dig.»
Och Mose bjöd folket på den dagen och sade:
Dessa stammar skola stå och välsigna folket på berget Gerissim, när I haven gått över Jordan: Simeon, Levi, Juda.
Isaskar, Josef och Benjamin.
Och dessa skola stå och uttala förbannelsen på berget Ebal: Ruben, Gad, Aser, Sebulon, Dan och Naftali.
Och leviterna skola taga till orda och skola med hög röst inför var man i Israel säga så:
Förbannad vare den man som gör ett beläte, skuret eller gjutet, en styggelse för HERREN, ett verk av en konstarbetares händer, och som sedan i hemlighet sätter upp det.
Och allt folket skall svara och säga: »Amen.»
Förbannad vare den som visar förakt för sin fader eller sin moder.
Och allt folket skall säga: »Amen.»
Förbannad vare den som flyttar sin nästas råmärke.
Och allt folket skall säga: »Amen.»
Förbannad vare den som leder en blind vilse på vägen.
Och allt folket skall säga: »Amen.»
Förbannad vare den som vränger rätten för främlingen, den faderlöse och änkan.
Och allt folket skall säga: »Amen.»
Förbannad vare den som ligger hos sin faders hustru, ty han lyfter på sin faders täcke.
Och allt folket skall säga: »Amen.»
Förbannad vare den som beblandar sig med något djur Och allt folket skall säga: »Amen.»
Förbannad vare den som ligger hos sin syster, sin faders dotter eller sin moders dotter.
Och allt folket skall säga: »Amen.»
Förbannad vare den som ligger hos sin svärmoder.
Och allt folket skall säga: »Amen.»
Förbannad vare den som lönnligen mördar sin nästa.
Och allt folket skall säga: »Amen.»
Förbannad vare den som tager mutor för att slå ihjäl en oskyldig och utgjuta hans blod.
Och allt folket skall säga: »Amen.»
Förbannad vare den som icke håller denna lags ord och icke gör efter dem.
Och allt folket skall säga: »Amen.»
Om du hör HERRENS, din Guds, röst, så att du håller alla hans bud, som jag i dag giver dig, och gör efter dem, så skall HERREN, din Gud, upphöja dig över alla folk på jorden.
Och alla dessa välsignelser skola då komma över dig och träffa dig när du hör HERRENS, din Guds, röst:
Välsignad skall du vara i staden, och välsignad skall du vara på marken.
Välsignad skall ditt livs frukt vara, och din marks frukt och din boskaps frukt, dina fäkreaturs avföda och din småboskaps avel.
Välsignad skall din korg vara, och välsignat ditt baktråg.
Välsignad skall du vara vid din ingång. och välsignad skall du vara vid din utgång.
När dina fiender resa sig upp mot dig, skall HERREN låta dem bliva slagna av dig; på en väg skola de draga ut mot dig, men på sju vägar skola de fly för dig.
HERREN skall bjuda välsignelsen vara med dig i dina visthus och i allt vad du företager dig; han skall välsigna dig i det land som HERREN, din Gud, vill giva dig.
HERREN skall upphöja dig till ett folk som är helgat åt honom, såsom han med ed har lovat dig, om du håller HERRENS, din Guds, bud och vandrar på hans vägar.
Och alla folk på jorden skola se att du är uppkallad efter HERRENS namn; och de skola frukta dig.
Och HERREN skall giva dig överflöd och lycka i ditt livs frukt och i din boskaps frukt och i din marks frukt, i det land som HERREN med ed har lovat dina fäder att giva dig.
HERREN skall öppna för dig sitt rika förrådshus, himmelen, till att giva åt ditt land regn i rätt tid, och till att välsigna alla dina händers verk; och du skall giva lån åt många folk, men själv skall du icke behöva låna av någon.
Och HERREN skall göra dig till huvud och icke till svans, du skall alltid ligga över och aldrig ligga under, om du hör HERRENS, din Guds, bud, som jag i dag giver dig, för att du skall hålla och göra efter dem,
och om du icke viker av, vare sig till höger eller till vänster, från något av alla de bud som jag i dag giver eder, så att du följer efter andra gudar och tjänar dem.
Men om du icke hör HERRENS, din Guds, röst och icke håller alla hans bud och stadgar, som jag i dag giver dig, och gör efter dem, så skola alla dessa förbannelser komma över dig och träffa dig:
Förbannad skall du vara i staden, och förbannad skall du vara på marken.
Förbannad skall din korg vara, och förbannat ditt baktråg.
Förbannad skall ditt livs frukt vara, och din marks frukt, dina fäkreaturs avföda och din småboskaps avel.
Förbannad skall du vara vid din ingång, och förbannad skall du vara vid din utgång.
HERREN skall sända över dig förbannelse, förvirring och näpst, vad det än må vara som du företager dig, till dess du förgöres och med hast förgås, för ditt onda väsendes skull, då du nu har övergivit mig.
HERREN skall låta dig bliva ansatt av pest, till dess han har utrotat dig ur det land dit du nu kommer, för att taga det i besittning.
HERREN skall slå dig med tärande sjukdom, feber och hetta, med brand och med svärd, med sot och rost; och av sådant skall du förföljas, till dess du förgås.
Och himmelen över ditt huvud skall vara såsom koppar, och jorden under dig skall vara såsom järn.
Damm och stoft skall vara det regn HERREN giver åt ditt land; från himmelen skall det komma ned över dig, till dess du förgöres.
HERREN skall låta dig bliva slagen av dina fiender; på en väg skall du draga ut mot dem, men på sju vägar skall du fly för dem; och du skall bliva en varnagel för alla riken på jorden.
Och dina dödas kroppar skola bliva mat åt alla himmelens fåglar och åt markens djur, och ingen skall skrämma bort dem.
HERREN skall slå dig med Egyptens bulnader och med bölder, med skabb och skorv, så att du icke skall kunna botas.
HERREN skall slå dig med vanvett och blindhet och sinnesförvirring.
Du skall famla mitt på ljusa dagen, såsom en blind famlar i mörkret, och du skall icke lyckas finna vägen; förtryck allenast och plundring skall du utstå i all din tid, och ingen skall frälsa dig.
Du skall trolova dig med en kvinna, men en annan man skall sova hos henne; du skall bygga ett hus, men icke få bo däri; du skall plantera en vingård, men icke få skörda dess frukt.
Din oxe skall slaktas inför dina ögon, men du skall icke få äta av den; din åsna skall i din åsyn rövas ifrån dig och icke givas tillbaka åt dig; dina får skola komma i dina fienders våld, och ingen skall hjälpa dig.
Dina söner och döttrar skola komma i främmande folks våld, och dina ögon skola se det och försmäkta av längtan efter dem beständigt, men du skall icke förmå göra något därvid.
Frukten av din mark och av allt ditt arbete skall förtäras av ett folk som du icke känner; förtryck allenast och övervåld skall du lida i all din tid.
Och du skall bliva vanvettig av de ting du skall se för dina ögon.
HERREN skall slå dig med svåra bulnader på knän och ben, ja, ifrån fotbladet ända till hjässan, så att du icke skall kunna botas.
HERREN skall föra dig och den konung som du sätter över dig bort till ett folk som varken du eller dina fäder hava känt, och där skall du få tjäna andra gudar, gudar av trä och sten.
Och du skall bliva ett föremål för häpnad, ett ordspråk och en visa bland alla de folk till vilka HERREN skall föra dig.
Mycken säd skall du föra ut på åkern, men litet skall du inbärga, ty gräshoppor skola förtära den.
Vingårdar skall du plantera och skall arbeta i dem, men intet vin skall du få att dricka och intet att lägga i förvar, ty maskar skola äta upp allt.
Olivplanteringar skall du hava överallt inom ditt land, men med oljan skall du icke få smörja din kropp, ty oliverna skola falla av.
Söner och döttrar skall du föda, men du skall icke få behålla dem, ty de skola draga bort i fångenskap.
Alla dina träd och din marks frukt skall ohyra taga i besittning.
Främlingen som bor hos dig skall höja sig över dig, allt mer och mer, men du skall stiga ned, allt djupare och djupare.
Han skall giva lån åt dig, och du skall icke giva lån åt honom.
Han skall bliva huvudet, och du skall bliva svansen.
Alla dessa förbannelser skola komma över dig och förfölja dig och träffa dig, till dess du förgöres, därför att du icke hörde HERRENS, din Guds, röst och icke höll de bud och stadgar som han har givit dig.
De skola komma över dig såsom tecken och under, och över dina efterkommande till evig tid.
Eftersom du icke tjänade HERREN, din Gud, med glädje och hjärtans lust, medan du hade överflöd på allt,
skall du få tjäna fiender som HERREN skall sända mot dig, under hunger och törst och nakenhet och brist på allt; och han skall lägga ett järnok på din hals, till dess han har förgjort dig.
HERREN skall skicka över dig ett folk fjärran ifrån, ifrån jordens ända. likt örnen i sin flykt,
ett folk vars språk du icke förstår, ett folk med grym uppsyn, utan försyn för de gamla och utan misskund med de unga.
Det skall äta upp frukten av din boskap och frukten av din mark, till dess du förgöres, ty det skall icke lämna kvar åt dig vare sig säd eller vin eller olja, icke dina fäkreaturs avföda eller dina fårs avel, till dess det har gjort slut på dig.
Och det skall tränga dig i alla dina portar, till dess dina höga och fasta murar, som du förtröstade på, falla i hela ditt land.
Ja, det skall tränga dig i alla dina portar över hela ditt land, det land som HERREN, din Gud, har givit dig.
Och då skall du nödgas äta din egen livsfrukt, köttet av dina söner och döttrar, dem som HERREN, din Gud, har givit dig.
I sådan nöd och sådant trångmål skall din fiende försätta dig.
En man hos dig, som levde i veklighet och stor yppighet, skall då så missunnsamt se på sin broder och på hustrun i sin famn och på de barn han ännu har kvar,
att han icke skall vilja åt någon av dem dela med sig av sina barns kött, ty han äter det själv, eftersom han icke har något annat kvar.
I sådan nöd och sådant trångmål skall din fiende försätta dig i alla dina portar.
En kvinna hos dig, som levde i veklighet och yppighet, i sådan yppighet och veklighet, att hon icke ens försökte sätta sin fot på jorden, hon skall då så missunnsamt se på mannen i sin famn och på sin son och sin dotter,
att hon missunnar dem efterbörden som kommer fram ur hennes liv, och barnen som hon föder; ty då hon nu lider brist på allt annat, skall hon själv i hemlighet äta detta.
I sådan nöd och sådant trångmål skall din fiende försätta dig i dina portar.
Om du icke håller alla denna lags ord, som äro skrivna i denna bok, och gör efter dem, så att du fruktar detta härliga och fruktansvärda namn »HERREN, din Gud»,
så skall HERREN sända underliga plågor över dig och dina efterkommande, stora och långvariga plågor, svåra och långvariga krankheter.
Han skall låta komma över dig alla Egyptens sjukdomar, som du fruktar för, och de skola ansätta dig.
Och allahanda andra krankheter och plågor, om vilka icke är skrivet i denna lagbok, skall HERREN ock låta gå över dig, till dess du förgöres.
Och allenast en ringa hop skall bliva kvar av eder, i stället för att I förut haven varit talrika såsom stjärnorna på himmelen; så skall det gå dig, därför att du icke hörde HERRENS. din Guds, röst.
Och det skall ske, att likasom HERREN förut fröjdade sig över eder när han fick göra eder gott och föröka eder, så skall HERREN nu fröjda sig över eder, när han utrotar och förgör eder.
Och I skolen ryckas bort ur det land dit du nu kommer, för att taga det i besittning.
Och HERREN skall förströ dig bland alla folk, ifrån jordens ena ända till den andra, och där skall du tjäna andra gudar, som varken du eller dina fäder hava känt, gudar av trä och sten.
Och bland de folken skall du icke få någon ro eller någon vila för din fot; HERREN skall där giva dig ett bävande hjärta och förtvinande ögon och en försmäktande själ.
Och ditt liv skall synas dig likasom hänga på ett hår; du skall känna fruktan både natt och dag och icke vara säker för ditt liv.
Om morgonen skall du säga: »Ack att det vore afton!», och om aftonen skall du säga: »Ack att det vore morgon!»
Sådan fruktan skall du känna i ditt hjärta, och sådana ting skall du se för dina ögon.
Och HERREN skall föra dig tillbaka till Egypten på skepp, på den väg om vilken jag sade dig: »Du skall icke se den mer.»
Och där skolen I nödgas bjuda ut eder till salu åt edra fiender, till trälar och trälinnor; men ingen skall finnas, som vill köpa.
Dessa äro förbundets ord, det förbunds som HERREN bjöd Mose att sluta med Israels barn i Moabs land, ett annat förbund än det som han hade slutit med dem på Horeb.
Och Mose sammankallade hela Israel och sade till dem: I haven sett allt vad HERREN har gjort inför edra ögon i Egyptens land, med Farao och alla hans tjänare och hela hans land,
de stora hemsökelser som du med egna ögon såg, de stora tecknen och undren.
Men HERREN har ännu intill denna dag icke givit eder hjärtan att förstå med, ögon att se med och öron att höra med.
Och jag lät eder vandra i öknen i fyrtio år; edra kläder blevo icke utslitna på eder, och din sko blev icke utsliten på din fot.
Bröd fingen I icke att äta, icke vin eller starka drycker att dricka, på det att I skullen veta att jag är HERREN, eder Gud.
Och när I kommen till dessa trakter, drogo Sihon, konungen i Hesbon, och Og, konungen i Basan, ut till strid mot oss, men vi slogo dem.
Och vi intogo deras land och gåvo det till arvedel åt rubeniterna, gaditerna och ena hälften av Manasse stam.
Så hållen nu detta förbunds ord och gören efter dem, för att I mån hava framgång i allt vad I gören.
I stån i dag allasammans inför HERREN, eder Gud: edra huvudmän, edra stammar, edra äldste och edra tillsyningsmän, var man i Israel,
så ock edra barn och hustrur, och främlingen som är hos dig i ditt läger, din vedhuggare såväl som din vattenbärare,
för att du må inträda i HERRENS, din Guds, förbund, det edsförbund som HERREN, din Gud, i dag vill sluta med dig.
Ty han vill i dag upphöja dig, så att du skall vara hans folk och han din Gud, såsom han har sagt dig, och såsom han med ed har lovat dina fäder, Abraham, Isak och Jakob.
Och det är icke med eder allenast som jag i dag sluter detta förbund, detta edsförbund,
utan jag gör det både med dem som i dag stå här med oss inför HERREN, vår Gud, och med dem som icke äro här med oss i dag.
I veten ju själva huru vi bodde i Egyptens land, och huru vi drogo mitt igenom de folks land, som I nu haven lämnat
Och I sågen deras styggelser och eländiga avgudar, de gudar av trä och sten, silver och guld, som funnos hos dem.
Så må då bland eder icke finnas någon man eller kvinna, någon släkt eller stam vars hjärta i dag vänder sig bort ifrån HERREN, vår Gud, för att gå åstad och tjäna dessa folks gudar; bland eder må icke finnas någon rot varifrån gift och malört växer upp,
så att någon som hör detta edsförbunds ord välsignar sig i sitt hjärta och tänker att det skall gå honom väl, där han vandrar i sitt hjärtas hårdhet.
Ty då skall hela landet, både vått och torrt, förgås.
HERREN skall icke vilja förlåta honom; nej, Herrens vrede och nitälskan skall då vara såsom en rykande eld mot de männen, och all den förbannelse som är uppskriven i denna bok skall komma att vila på honom, och Herren skall så utplåna hans namn, att det icke mer skall finnas under himmelen.
Och HERREN skall avskilja honom från alla Israels stammar till att drabbas av olycka, efter alla de förbannelser som äro fästa vid det förbund som är uppskrivet i denna lagbok.
Och ett kommande släkte, edra barn som uppstå efter eder, och främlingen, som kommer ifrån fjärran land, de skola säga, när de se de plågor och sjukdomar som HERREN har skickat över detta land,
när de se huru all jord där är förbränd och förvandlad till svavel och salt, så att den icke kan besås eller framalstra växter, och så att inga örter där kunna komma upp -- såsom det blev, när Sodom och Gomorra, Adma och Seboim omstörtades, då HERREN i sin vrede och harm omstörtade dem --
ja, alla folk skola då säga: »Varför har Herren gjort så mot detta land?
Varför brinner hans vrede så starkt?»
Och man skall svara: »Därför att de övergåvo HERRENS, sina fäders Guds, förbund, det som han slöt med dem, när han förde dem ut ur Egyptens land,
och därför att de gingo åstad och tjänade andra gudar och tillbådo dem, gudar som de icke kände, och som han icke hade givit dem till deras del,
därför upptändes HERRENS vrede mot detta land, så att han lät komma över det all den förbannelse som är uppskriven i denna bok.
Ja, därför ryckte HERREN dem upp ur deras land, med vrede och harm och stor förtörnelse, och kastade dem bort till ett annat land, såsom nu har skett.»
Vad som ännu är fördolt hör HERREN, vår Gud, till; men vad som är uppenbarat, det gäller för oss och våra barn till evig tid, för att vi skola göra efter alla denna lags ord.
Om du nu, när allt detta kommer över dig -- välsignelsen och förbannelsen som jag har förelagt dig -- om du lägger detta på hjärtat bland alla de folk till vilka HERREN, din Gud, då har drivit dig bort,
och du så vänder åter till HERREN, din Gud, och hör hans röst, du med dina barn, av allt ditt hjärta och av all din själ, i alla stycken såsom jag i dag bjuder dig,
då skall HERREN, din Gud, åter upprätta dig och förbarma sig över dig; HERREN, din Gud, skall då åter församla dig från alla folk bland vilka han har förstrött dig.
Om ock dina fördrivna vore vid himmelens ända, skulle HERREN, din Gud, församla dig därifrån och hämta dig därifrån.
Och HERREN, din Gud, skall låta dig komma in i det land som dina fäder hava haft till besittning; och du skall taga det i besittning, och han skall göra dig gott och skall föröka dig mer än han har gjort med dina fäder.
Och HERREN, din Gud. skall omskära ditt hjärta och dina efterkommandes hjärtan, så att du skall älska HERREN, din Gud, av allt ditt hjärta och av all din själ, för att du må leva.
Och HERREN, din Gud, skall lägga alla dessa förbannelser på dina fiender och på dem som hata och förfölja dig.
Och du skall åter höra HERRENS röst och göra efter alla hans bud, som jag i dag giver dig.
Och HERREN, din Gud, skall giva dig överflöd och lycka i alla dina händers verk, i ditt livs frukt och i din boskaps frukt och i din marks frukt.
Ty såsom HERREN fröjdade sig över dina fäder, skall han då åter fröjda sig över dig och göra dig gott,
när du hör HERRENS, din Guds, röst, så att du håller hans bud och stadgar, det som är skrivet i denna lagbok, och när du vänder åter till HERREN, din Gud, av allt ditt hjärta och av all din själ.
Ty det bud som jag i dag giver dig är dig icke för svårt och är icke långt borta.
Det är icke i himmelen, så att du skulle behöva säga: »Vem vill för oss fara upp till himmelen och hämta det åt oss och låta oss höra det, så att vi kunna göra därefter?»
Det är icke heller på andra sidan havet, så att du skulle behöva säga: »Vem vill för oss fara över till andra sidan havet och hämta det åt oss och låta oss höra det, så att vi kunna göra därefter?»
Nej, ordet är dig mycket nära, i din mun och i ditt hjärta, så att du kan göra därefter.
Se, jag förelägger dig i dag livet och vad gott är, döden och vad ont är,
då jag nu i dag bjuder dig att älska HERREN, din Gud, att vandra på hans vägar och hålla hans bud och stadgar och rätter, för att du må leva och föröka dig, och för att HERREN, din Gud, må välsigna dig i det land dit du nu kommer, för att taga det i besittning.
Men om ditt hjärta vänder sig bort och du icke vill höra, om du låter förföra dig, så att du tillbeder andra gudar och tjänar dem,
så förkunnar jag eder i dag att I förvisso skolen förgås.
I skolen då icke länge leva i det land dit du nu drager över Jordan, för att komma och taga det i besittning.
Jag tager i dag himmel och jord till vittnen mot eder, att jag har förelagt dig liv och död, välsignelse och förbannelse, Så må du då välja livet, för att du och dina efterkommande mån leva,
i det att du älskar HERREN, din Gud, och hör hans röst och håller dig till honom; ty detta betyder för dig liv och lång levnad, så att du får bo i det land som HERREN med ed har lovat dina fäder, Abraham, Isak och Jakob, att giva dem.
Och Mose gick åstad och talade följande till hela Israel;
han sade till dem: »Jag är nu ett hundra tjugu år gammal; jag kan icke mer vara ledare och anförare, och HERREN har sagt till mig: 'Du skall icke komma över denna Jordan.'
Men HERREN, din Gud, går framför dig; han skall förgöra dessa folk för dig, och du skall fördriva dem, och Josua skall anföra dig, såsom HERREN har sagt.
Och HERREN skall göra med dem såsom han gjorde med Sihon och Og, amoréernas konungar. vilka han lät förgås, och såsom han gjorde med deras land.
HERREN skall giva dem i edert våld, och I skolen göra med dem alldeles såsom jag har bjudit eder.
Varen frimodiga och oförfärade, frukten icke och varen icke förskräckta för dem; ty HERREN, din Gud, går själv med dig; han skall icke lämna dig eller övergiva dig.»
Och Mose kallade Josua till sig och sade till honom inför hela Israel: »Var frimodig och oförfärad; ty du skall med detta folk gå in i det land som HERREN med ed har lovat deras fäder att giva dem; och du skall utskifta det åt dem såsom arv.
Och HERREN är den som går framför dig, han skall vara med dig, han skall icke lämna dig eller övergiva dig; du må icke frukta och icke vara förfärad.»
Och Mose skrev upp denna lag och gav den åt prästerna, Levi söner, som buro HERRENS förbundsark, och åt alla de äldste i Israel.
Och Mose bjöd dem och sade: »Vid slutet av vart sjunde år, när friåret är inne, vid lövhyddohögtiden,
då hela Israel kommer för att träda fram inför HERRENS, din Guds, ansikte, på den plats som han utväljer, då skall du läsa upp denna lag inför hela Israel, så att de höra den.
Församla då folket, män, kvinnor och barn, och främlingarna som äro hos dig inom dina portar, på det att de må höra och lära, och på det att de må frukta HERREN, eder Gud, och hålla och göra efter alla denna lags ord;
och på det att deras barn, som då ännu icke känna den, må höra den och lära den, så att de frukta HERREN, eder Gud.
Detta skolen I göra, så länge I leven i det land dit I nu dragen över Jordan, för att taga det i besittning.
Och HERREN sade till Mose: »Se, tiden närmar sig att du skall dö.
Kalla till dig Josua, och inställen eder därefter i uppenbarelsetältet, så vill jag insätta honom i hans ämbete.»
Och Mose gick åstad med Josua, och de inställde sig i uppenbarelsetältet.
Då visade sig HERREN i tältet i en molnstod, och molnstoden blev stående vid ingången till tältet.
Och HERREN sade till Mose: »Se, när du vilar hos dina fäder, skall detta folk stå upp och i trolös avfällighet löpa efter främmande gudar, som dyrkas i det land dit de nu komma, och de skola övergiva mig och bryta det förbund som jag har slutit med dem.
Och min vrede skall då upptändas mot dem, och jag skall övergiva dem och fördölja mitt ansikte för dem, och de skola förgöras, och mycken olycka och nöd skall träffa dem; och då skola de säga: 'Förvisso är det därför att vår Gud icke är ibland oss som dessa olyckor hava träffat oss.'
Men jag skall på den tiden alldeles fördölja mitt ansikte, för allt det ondas skull som de hava gjort, i det att de hava vänt sig till andra gudar.
Så tecknen nu upp åt eder följande sång.
Och du skall lära Israels barn den och lägga den i deras mun.
Och så skall denna sång vara mig ett vittne mot Israels barn.
Ty jag skall låta dem komma in i det land som jag med ed har lovat åt deras fäder, ett land som flyter av mjölk och honung, och de skola äta och bliva mätta och feta; men de skola då vända sig till andra gudar och tjäna dem och förakta mig och bryta mitt förbund.
Och när då mycken olycka och nöd träffar dem, skall denna sång avlägga sitt vittnesbörd inför dem; ty den skall icke förgätas och försvinna ur deras avkomlingars mun.
Jag vet ju med vilka tankar de umgås redan nu, innan jag har låtit dem komma in i det land som jag med ed lovade dem.»
Så tecknade då Mose upp sången på den dagen och lät Israels barn lära den.
Och han insatte Josua, Nuns son, i hans ämbete och sade: »Var frimodig och oförfärad; ty du skall föra Israels barn in i det land som jag med ed har lovat åt dem, och jag skall vara med dig.»
Då nu Mose hade fullständigt tecknat upp denna lags ord i en bok,
bjöd han leviterna som buro HERRENS förbundsark och sade:
»Tagen denna lagbok och läggen den vid sidan av HERRENS, eder Guds, förbundsark, så att den ligger där till ett vittne mot dig.
Ty jag känner din gensträvighet och hårdnackenhet.
Se, ännu medan jag har levat kvar bland eder, haven I varit gensträviga mot HERREN; huru mycket mer skolen I ej då bliva det efter min död!
Församlen nu till mig alla de äldste i edra stammar, så ock edra tillsyningsmän, för att jag må inför dem tala dessa ord och taga himmel och jord till vittnen mot dem.
Ty jag vet att I efter min död skolen taga eder till, vad fördärvligt är, och vika av ifrån den väg som jag har bjudit eder gå; därför skall olycka träffa eder i kommande dagar, när I gören vad ont är i HERRENS ögon, så att I förtörnen honom genom edra händers verk.»
Och Mose föredrog inför Israels hela församling följande sång från början till slutet.
Lyssnen, I himlar, ty jag vill tala; och jorden höre min muns ord.
Såsom regnet drype min lära, såsom daggen flöde mitt tal, såsom rikligt regn på grönska och såsom en regnskur på gräsets brodd.
Ty HERRENS namn vill jag förkunna; ja, given ära åt vår Gud.
Vår klippa -- ostraffliga äro hans gärningar, ty alla hans vägar äro rätta.
En trofast Gud och utan svek, rättfärdig och rättvis är han.
De åter handlade illa mot honom; de voro icke hans barn, utan en skam för Israel, det vrånga och avoga släktet!
Är det så du lönar HERREN, du dåraktiga och ovisa folk?
Är han då icke din fader, som skapade dig?
Han danade ju dig och beredde dig.
Tänk på de dagar som fordom voro; akta på förgångna släktens år.
Fråga din fader, han skall förkunna dig det, dina äldste, de skola säga dig det.
När den Högste gav arvslotter åt folken, när han fördelade människors barn, då utstakade han gränserna för folken efter antalet av Israels barn.
Ty HERRENS folk är hans del, Jakob är hans arvedels lott.
Han fann honom i öknens land, i ödsligheten, där ökendjuren tjöto.
Då tog han honom i sitt beskärm och sin vård, han bevarade honom såsom sin ögonsten.
Likasom en örn lockar sin avkomma ut till flykt och svävar upp ovanför sina ungar, så bredde han ut sina vingar och tog honom och bar honom på sina fjädrar.
HERREN allena ledsagade honom, och ingen främmande gud jämte honom.
Han förde honom fram över landets höjder och lät honom äta av markens gröda; han lät honom suga honung ur hälleberget och olja ur den hårda klippan.
Gräddmjölk av kor, söt mjölk av får, fett av lamm fick du ock, vädurar från Basan och bockar, därtill fetaste märg av vete; och av druvors blod drack du vin.
Då blev Jesurun fet och istadig; du blev fet och tjock och stinn.
Han övergav Gud, sin skapare, och föraktade sin frälsnings klippa.
Ja, de retade honom genom sina främmande gudar, med styggelser förtörnade de honom.
De offrade åt onda andar, skengudar, åt gudar som de förut icke kände, nya, som nyss hade kommit till, och som edra fäder ej fruktade för.
Din klippa, som hade fött dig, övergav du, du glömde Gud, som hade givit dig livet.
När HERREN såg detta, förkastade han dem, ty han förtörnades på sina söner och döttrar.
Han sade: »Jag vill fördölja mitt ansikte för dem, jag vill se vilket slut de få; ty ett förvänt släkte äro de, barn i vilka ingen trohet är.
De hava retat mig med gudar som icke äro gudar, förtörnat mig med de fåfängligheter de dyrka; därför skall jag reta dem med ett folk som icke är ett folk, med ett dåraktigt hednafolk skall jag förtörna dem.
Ty eld lågar fram ur min näsa, och den brinner ända till dödsrikets djup; den förtär jorden med dess gröda och förbränner bergens grundvalar.
Jag skall hopa olyckor över dem, alla mina pilar skall jag avskjuta på dem.
De skola utsugas av hunger och förtäras av feberglöd, av farsoter som bittert pina; jag skall sända över dem vilddjurs tänder och stoftkrälande ormars gift.
Ute skall svärdet förgöra deras barn, och inomhus skall förskräckelsen göra det: ynglingar såväl som jungfrur, spenabarn tillsammans med gråhårsmän.
Jag skulle säga: 'Jag vill blåsa bort dem, göra slut på deras åminnelse bland människor',
om jag icke fruktade att deras fiender då skulle vålla mig grämelse, att deras ovänner skulle misstyda det, att de skulle säga: 'Vår hand var så stark, det var icke HERREN som gjorde allt detta.'»
Ty ett rådlöst folk äro de, och förstånd finnes icke i dem.
Vore de visa, så skulle de begripa detta, de skulle första vilket slut de måste få.
Huru kunde en jaga tusen framför sig och två driva tiotusen på flykten, om icke deras klippa hade sålt dem, och om icke HERREN hade prisgivit dem?
Ty de andras klippa är icke såsom vår klippa; våra fiender kunna själva döma därom.
Ty av Sodoms vinträd är deras ett skott, det stammar från Gomorras fält; deras druvor äro giftiga druvor, deras klasar hava bitter smak.
Deras vin är drakars etter, huggormars gruvligaste gift.
Ja, sådant ligger förvarat hos mig, förseglat i mina förrådshus.
Min är hämnden och vedergällningen, sparad till den tid då deras fot skall vackla.
Ty nära är deras ofärds dag, och vad dem väntar kommer med hast.
Ty HERREN skall skaffa rätt åt sitt folk, och över sina tjänare skall han förbarma sig, när han ser att deras kraft är borta, och att det är ute med alla och envar.
Då skall han fråga: Var äro nu deras gudar, klippan till vilken de togo sin tillflykt?
Var äro de som åto deras slaktoffers fett och drucko deras drickoffers vin?
Må de stå upp och hjälpa eder, må de vara edert beskärm.
Sen nu att jag allena är det, och att ingen Gud finnes jämte mig.
Jag dödar, och jag gör levande, jag har slagit, men jag helar ock.
Ingen finnes, som kan rädda ur min hand.
Se, jag lyfter min hand upp mot himmelen, jag säger: Så sant jag lever evinnerligen:
när jag har vässt mitt ljungande svärd och min hand tager till att skipa rätt, då skall jag utkräva hämnd av mina ovänner och vedergällning av dem som hata mig.
Jag skall låta mina pilar bliva druckna av blod, och mitt svärd skall mätta sig av kött, av de slagnas och fångnas blod, av fiendehövdingars huvuden.
Jublen, I hedningar, över hans folk, ty han hämnas sina tjänares blod, han utkräver hämnd av sina ovänner och bringar försoning för sitt land, för sitt folk.
Och Mose kom med Hosea, Nuns son, och föredrog hela denna sång inför folket.
Och när Mose hade föredragit alltsammans till slut för hela Israel,
sade han till dem: »Akten på alla de ord som jag i dag gör till vittnen mot eder, så att I given edra barn befallning om dem, att de skola hålla alla denna lags ord och göra efter dem.
Ty det är icke ett tomt ord, som ej angår eder, utan det gäller edert liv; och genom detta ord skolen I länge leva i det land dit I nu dragen över Jordan, för att taga det i besittning.»
Och HERREN talade till Mose på denna samma dag och sade:
»Stig upp här på Abarimberget, på berget Nebo i Moabs land, gent emot Jeriko, så skall du få se Kanaans land, som jag vill giva åt Israels barn till besittning.
Och du skall dö där på berget, dit du stiger upp, och du skall samlas till dina fäder, likasom din broder Aron dog på berget Hor och blev samlad till sina fäder;
detta därför att I handladen trolöst mot mig bland Israels barn vid Meribas vatten vid Kades, i öknen Sin, i det att I icke höllen mig helig bland Israels barn.
Mitt framför dig skall du se landet; men du skall icke komma dit, in i det land som jag vill giva åt Israels barn.»
Och detta är den välsignelse gudsmannen Mose gav Israels barn före sin död;
han sade: »HERREN kom från Sinai, och från Seir gick hans sken upp för dem; man kom fram i glans från berget Paran, ut ur hopen av mångtusen heliga; på hans högra sida brann i eld en lag för dem.
Ja, han vårdar sig om folken; folkets heliga äro alla under din hand.
De ligga vid din fot, de hämta upp av dina ord.
Mose gav åt oss en lag, en arvedel for Jakobs menighet.
Och Jesurun fick en konung, när folkets hövdingar församlades, Israels stammar allasammans.»
»Må Ruben leva och icke dö; dock blive hans män en ringa hop.
Och detta sade han om Juda: »Hör, o HERRE, Judas röst, och låt honom komma till sitt folk.
Med sina händer utförde han dess sak; bliv du honom en hjälp mot hans ovänner.»
Och om Levi sade han: »Dina tummim och dina urim, de tillhöra din frommes skara, dem du frestade i Massa, dem du tvistade med vid Meribas vatten,
dem som sade om fader och moder: 'Jag ser dem icke', och som icke ville kännas vid sina bröder, ej heller veta av sina barn.
Ty de aktade på ditt tal, och ditt förbund höllo de.
De lära Jakob dina rätter och Israel din lag, de bära fram rökverk för din näsa och heloffer på ditt altare.
Välsigna, HERRE, hans kraft, och låt hans händers verk behaga dig.
Krossa länderna på hans motståndare, på hans fiender, så att de icke kunna resa sig.»
Om Benjamin sade han: »HERRENS vän är han, han skall bo i trygghet hos honom, hos honom som överskygger honom alltid, och som har sin boning mellan hans höjder.»
Och om Josef sade han: »Välsignat av HERREN vare hans land med himmelens ädlaste gåvor, med dagg, med gåvor från djupet som utbreder sig därnere,
med solens ädlaste alster och månvarvens ädlaste frukter,
med de uråldriga bergens yppersta skatter och de eviga höjdernas ädlaste frukt,
med jordens ädlaste frukt och allt vad hon bär, och med nåd från honom som bodde i busken.
Detta komme över Josefs huvud, över hans hjässa, furstens bland bröder.
Härlig är den förstfödde bland hans tjurar, såsom en vildoxes äro hans horn; med dem stångar han ned alla folk, ja ock dem som bo vid jordens ändar.
Sådana äro Efraims tiotusenden. sådana Manasses tusenden.»
Och om Sebulon sade han: »Gläd dig, Sebulon, när du drager ut, och du, Isaskar, i dina tält.
Folk inbjuda de till sitt berg; där offra de rätta offer.
Ty havens rikedom få de suga, och de skatter som sanden döljer.»
Och om Gad sade han: »Lovad vare han som gav så rymligt land åt Gad!
Lik en lejoninna har han lägrat sig, han krossar både arm och hjässa.
Han utsåg åt sig förstlingslandet, ty där var hans härskarlott förvarad.
Dock drog han med bland folkets hövdingar; HERRENS rätt utförde han och hans domar, tillsammans med det övriga Israel.»
Och om Dan sade han: »Dan är ett ungt lejon, som rusar ned från Basan.»
Och om Naftali sade han: »Naftali har fått riklig nåd och välsignelse till fyllest av HERREN.
Västern och södern tage du i besittning.»
Och om Aser sade han: »Välsignad bland söner vare Aser!
Han blive älskad av sina bröder, och han doppe sin fot i olja.
Av järn och koppar vare dina riglar; och så länge du lever, må din kraft bestå.»
»Ingen är lik Gud, o Jesurun; till din hjälp far han fram på himmelen och i sin höghet på skyarna.
En tillflykt är han, urtidens Gud, och härnere råda hans eviga armar.
Han förjagade fienderna för dig, han sade: Förgör dem.
Så fick Israel bo i trygghet, Jakobs källa vara i ro, i ett land med säd och vin, under en himmel som dryper av dagg.
Säll är du, Israel; ja, vem är dig lik?
Du är ett folk som får seger genom HERREN, genom honom som är din skyddande sköld, honom som är ditt ärorika svärd.
Ja, dina fiender skola visa dig underdånighet, och du skall gå fram över deras höjder.»
Och Mose gick från Moabs hedar upp på berget Nebo, på toppen av Pisga, gent emot Jeriko.
Och HERREN lät honom se hela landet: Gilead ända till Dan,
och hela Naftali och Efraims och Manasses land, och hela Juda land, ända till Västra havet,
och Sydlandet och Jordanslätten, det är lågslätten vid Jeriko -- Palmstaden -- ända till Soar.
Och HERREN sade till honom: »Detta är det land som jag med ed har lovat åt Abraham.
Isak och Jakob, i det jag sade: 'Åt din säd skall jag giva det.'
Jag har nu låtit dig se det med dina ögon, men ditin skall du icke komma.»
Och HERRENS tjänare Mose dog där i Moabs land, såsom HERREN hade sagt.
Och han begrov honom i dalen i Moabs land, mitt emot Bet-Peor; men ännu intill denna dag har ingen fått veta var hans grav är.
Och Mose var ett hundra tjugu år gammal, när han dog, men hans ögon voro icke skumma, och hans livskraft hade icke försvunnit.
Och Israels barn begräto Mose på Moabs hedar i trettio dagar; därmed voro gråtodagarna ute, vid sorgefesten efter Mose.
Och Josua, Nuns son, var full med vishetens ande, ty Mose hade lagt sina händer på honom; och Israels barn lydde honom och gjorde såsom HERREN hade bjudit Mose.
Men i Israel uppstod icke mer någon profet sådan som Mose, med vilken HERREN hade umgåtts ansikte mot ansikte --
ingen, om man tänker på alla de tecken och under som HERREN hade sänt honom att göra i Egyptens land, med Farao och alla hans tjänare och med hela hans land,
och om man tänker på all den väldiga kraft som Mose visade, och på alla de stora och fruktansvärda gärningar som han gjorde inför hela Israel.
Efter HERRENS tjänare Moses död sade HERREN till Josua, Nuns son, Moses tjänare:
»Min tjänare Mose är död; så stå nu upp och gå över denna Jordan, du med allt detta folk, in i det land som jag vill giva dem, giva åt Israels barn.
Var ort som eder fot beträder har jag givit eder, såsom jag lovade Mose.
Från öknen till Libanon däruppe och ända till den stora floden, floden Frat, över hetiternas land och ända till Stora havet västerut skall edert område sträcka sig.
Ingen skall kunna stå dig emot i alla dina livsdagar; såsom jag har varit med Mose, så skall jag ock vara med dig; jag skall icke lämna dig eller övergiva dig.
Var frimodig och oförfärad; ty du skall utskifta åt detta folk såsom arv det land som jag med ed har lovat deras fäder att giva dem.
Allenast må du vara helt frimodig och oförfärad till att i alla stycken hålla den lag som min tjänare Mose har givit dig och göra efter den; vik icke av därifrån vare sig till höger eller till vänster; på det att du må hava framgång i allt vad du företager dig.
Låt icke denna lagbok vara skild från din mun; tänk på den både dag och natt, så att du i alla stycken håller det som är skrivet i den och gör därefter; ty då skola dina vägar vara lyckosamma, och då skall du hava framgång.
Se, jag har bjudit dig att vara frimodig och oförfärad; så var nu icke förskräckt eller försagd.
Ty HERREN, din Gud, är med dig i allt vad du företager dig.»
Då bjöd Josua folkets tillsyningsmän och sade:
»Gån igenom lägret och bjuden folket och sägen: 'Reden till reskost åt eder; ty om tre dagar skolen I gå över denna Jordan, för att komma in i och taga i besittning det land som HERREN, eder Gud, vill giva eder till besittning.'»
Men till rubeniterna och gaditerna och ena hälften av Manasse stam sade Josua:
»Tänken på det som HERRENS tjänare Mose bjöd eder, när han sade: 'HERREN, eder Gud, vill låta eder komma till ro och giva eder detta land.'
Edra hustrur, edra barn och eder boskap må nu stanna kvar i det land som Mose har givit eder här på andra sidan Jordan; men I själva, så många av eder som äro tappra stridsmän, skolen draga väpnade åstad i spetsen för edra bröder och hjälpa dem,
till dess att HERREN har låtit edra bröder komma till ro såväl som eder, när också de hava tagit i besittning det land som HERREN, eder Gud, vill giva dem.
Sedan mån I vända tillbaka till det land som skall vara eder besittning; det mån I då taga i besittning, det land som HERRENS tjänare Mose har givit eder här på andra sidan Jordan, på östra sidan.»
Då svarade de Josua och sade: »Allt vad du har bjudit oss vilja vi göra, och varthelst du sänder oss, dit vilja vi gå.
Såsom vi i allt hava lytt Mose, så vilja vi ock lyda dig; allenast må HERREN, din Gud, vara med dig, såsom han var med Mose.
Var och en som är gensträvig mot dina befallningar och icke lyssnar till dina ord, vadhelst du bjuder honom, han skall bliva dödad.
Allenast må du vara frimodig och oförfärad.»
Josua, Nuns son, sände hemligen ut två spejare från Sittim och sade: »Gån och besen landet och Jeriko.»
De gingo åstad och kommo in i ett hus där en sköka bodde, vid namn Rahab, och där lade de sig till vila.
Men för konungen i Jeriko blev inberättat: »I natt hava några män kommit hit från Israels barn för att utforska landet.»
Då sände konungen i Jeriko till Rahab och lät säga: »Lämna ut de män som hava kommit till dig och tagit in i ditt hus, ty de hava kommit hit för att utforska hela landet.»
Men kvinnan tog de båda männen och dolde dem; sedan svarade hon: »Ja, männen kommo till mig, men jag visste icke varifrån de voro;
och när porten skulle stängas, sedan det hade blivit mörkt, gingo männen ut, och jag vet icke vart de togo vägen; skynden eder att sätta efter dem, så fån I nog fatt i dem.»
Men hon hade fört dem upp på taket och gömt dem under linstjälkar, som hon hade där, utbredda på taket.
Så satte nu männen efter dem åt Jordan till, bort emot vadställena; och man stängde stadsporten så snart förföljarna hade begivit sig åstad.
Men innan de främmande männen hade lagt sig, steg hon upp till dem på taket
och sade till dem: »Jag vet att HERREN har givit eder detta land, och att förskräckelse för eder har fallit över oss, ja, att alla landets inbyggare äro i ångest för eder.
Ty vi hava hört huru HERREN lät vattnet i Röda havet torka ut framför eder, när I drogen ut ur Egypten, och vad I haven gjort med amoréernas konungar, de två på andra sidan Jordan, Sihon och Og, huru I gåven dem till spillo.
Då vi hörde detta, blevo våra hjärtan förfärade, och numera har ingen mod att stå eder emot; ty HERREN, eder Gud, är Gud, uppe i himmelen och nere på jorden.
Så loven mig nu med ed vid HERREN, att eftersom jag har gjort barmhärtighet med min faders hus och giva mig ett säkert tecken därpå,
och låta min fader och min moder, mina bröder och mina systrar leva, så ock alla som tillhöra dem, och rädda oss från döden.»
Männen sade till henne: »Med vårt eget liv svara vi för edert, såframt I icke förråden vårt förehavande; när HERREN giver oss landet, skola vi bevisa dig barmhärtighet och trofasthet.»
Då släppte hon ned dem genom fönstret med ett tåg; ty hennes hus låg invid stadsmuren, så att hon bodde invid själva muren.
Och hon sade till dem: »Gån upp i bergsbygden, så att edra förföljare icke träffa på eder; och hållen eder gömda där i tre dagar, till dess edra förföljare hava kommit tillbaka, så kunnen I sedan fortsätta eder färd.»
Och männen sade till henne: »Vi vilja likväl vara fria ifrån den ed som du nu har tagit av oss,
om du, när vi komma in i landet, underlåter att binda detta röda snöre i det fönster genom vilket du har släppt ned oss, och likaledes om du icke har din fader och din moder och dina bröder, alla av din faders hus, samlade hemma hos dig.
Dock, om någon går åstad, utom dörrarna till ditt hus, så komme hans blod över hans huvud, och vi äro utan skuld; om däremot någons hand kommer vid en av dem som äro inne i ditt hus, så må dennes blod komma över vårt huvud.
Och om du förråder vårt förehavande, så äro vi likaledes fria ifrån den ed som du har tagit av oss.»
Hon svarade: »Vare det såsom I haven sagt.»
Och så lät hon dem gå, och de drogo åstad.
Men hon band det röda snöret i fönstret.
Så drogo de nu åstad och kommo upp i bergsbygden och stannade där i tre dagar, till dess att deras förföljare hade vänt tillbaka; ty dessa hade sökt efter dem överallt på vägarna, men hade icke funnit dem.
Sedan vände de båda männen tillbaka och kommo ned från bergsbygden och gingo över floden och kommo så till Josua, Nuns son; och de förtäljde för honom allt vad som hade vederfarits dem.
Och de sade till Josua: »HERREN har givit hela landet i vår hand; alla landets inbyggare äro i ångest för oss.»
Bittida följande morgon bröt Josua med alla Israels barn upp från Sittim och kom till Jordan; där stannade de om natten, innan de gingo över.
Men efter tre dagar gingo tillsyningsmännen genom lägret
och bjödo folket och sade: »Så snart I fån se HERRENS, eder Guds, förbundsark, och att de levitiska prästerna bära den, skolen ock I bryta upp från eder plats och följa efter den
-- låten dock mellan den och eder vara ett avstånd av vid pass två tusen alnar; närmare mån I icke komma den -- på det att I mån kunna veta vilken väg I skolen gå, ty I haven icke förut dragit den vägen fram.»
Och Josua sade till folket: »Helgen eder, ty i morgon skall HERREN göra under bland eder.»
Därefter sade Josua till prästerna: »Tagen förbundsarken och dragen åstad framför folket.»
Då togo de förbundsarken och gingo framför folket.
Och HERREN sade till Josua: »I dag skall jag begynna att göra dig stor i hela Israels ögon, på det att de må förnimma, att såsom jag har varit med Mose, så vill jag ock vara med dig.
Bjud du nu prästerna som bära förbundsarken och säg: 'Så snart I kommen till den yttersta randen av Jordans vatten, skolen I stanna där, vid Jordan.'»
Då sade Josua till Israels barn: »Träden fram hit och hören HERRENS, eder Guds, ord.»
Och Josua sade: »Härav skolen I förnimma att en levande Gud är mitt ibland eder, och att han förvisso vill fördriva för eder kananéerna, hetiterna, hivéerna, perisséerna, girgaséerna, amoréerna och jebuséerna:
förbundsarken, hela jordens Herres förbundsark, drager nu framför eder över Jordan.
Väljen alltså ut tolv män ur Israels stammar, en man för var stam.
Så snart då prästerna som bära HERRENS, hela jordens Herres, ark stå stilla med sina fötter i Jordans vatten, det vatten som kommer uppifrån, bliva avskuret i sitt lopp, och det skall stå såsom en samlad hög.»
Folket bröt då upp från sina tält för att gå över Jordan, och prästerna som buro förbundsarken gingo framför folket.
När nu de som buro arken kommo till Jordan, så att prästerna, som buro arken, med sina fötter vidrörde yttersta randen av vattnet i Jordan, vilken under hela skördetiden är full över alla sina bräddar,
då stannade det vatten som kom uppifrån, och blev stående såsom en samlad hög långt borta, uppe vid Adam, staden som ligger bredvid Saretan; och det vatten som flöt ned mot Hedmarkshavet, Salthavet, blev sålunda helt och hållet avskuret.
Och folket gick över mitt emot Jeriko.
Men prästerna som buro HERRENS förbundsark stodo orörliga på torr mark mitt i Jordan; och hela Israel gick över på torr mark, till dess att allt folket helt och hållet hade kommit över Jordan.
Då nu allt folket helt och hållet hade kommit över Jordan, sade HERREN till Josua:
»Väljen ut bland folket tolv män, en man ur var stam,
och bjuden dem och sägen: 'Tagen här ur Jordan, från den plats där prästerna stodo med sina fötter, tolv stenar, och lyften upp dem och fören dem över med eder, och läggen ned dem på det ställe, där I skolen lägra eder i natt.'»
Då kallade Josua till sig de tolv män som han hade utsett bland Israels barn, en man ur var stam.
Och Josua sade till dem: »Dragen åstad framför HERRENS, eder Guds, ark, och gån ut mitt i Jordan; och var och en av eder må där lyfta upp en sten på axeln, efter antalet av Israels barns stammar.
Detta skall nämligen bliva ett minnesmärke bland eder.
När då edra barn i framtiden fråga: 'Vad betyda dessa stenar?',
skolen I svara dem så: 'De betyda att Jordans vatten här blev avskuret i sitt lopp, framför HERRENS förbundsark; ja, när den gick över Jordan, blev Jordans vatten avskuret i sitt lopp.
Därför skola dessa stenar vara ett åminnelsemärke för Israels barn till evärdlig tid.'»
Då gjorde Israels barn såsom Josua bjöd dem; de togo upp tolv stenar ur Jordan, såsom HERREN hade tillsagt Josua, efter antalet av Israels barns stammar; och de förde dem över med sig till lägerstället och lade ned dem där.
Tillika reste Josua tolv stenar mitt i Jordan, på samma plats där prästerna som buro förbundsarken hade stått med sina fötter; och de finnas kvar där ännu i dag.
Och prästerna som buro arken blevo stående mitt i Jordan, till dess att allt det var fullgjort, som HERREN hade bjudit Josua att tillsäga folket, alldeles i enlighet med vad Mose förut hade bjudit Josua; och folket gick över med hast.
Men när allt folket helt och hållet hade kommit över, gick ock HERRENS ark över, jämte prästerna, och tog plats framför folket.
Och Rubens barn och Gads barn och ena hälften av Manasse stam drogo väpnade åstad i spetsen för Israels barn, såsom Mose hade tillsagt dem.
Det var vid pass fyrtio tusen män som så drogo åstad, väpnade till strid, för att kämpa inför HERREN på Jerikos hedmarker.
På den dagen gjorde HERREN Josua stor i hela Israels ögon, och de fruktade honom, såsom de fruktat Mose, så länge denne levde.
Och HERREN sade till Josua:
»Bjud prästerna som bära vittnesbördets ark att stiga upp ur Jordan.»
Och Josua bjöd prästerna och sade: »Stigen upp ur Jordan.»
När då prästerna som buro HERRENS förbundsark stego upp ur Jordan, hade deras fötter knappt hunnit upp på torra landet, förrän Jordans vatten vände tillbaka till sin plats och nådde, såsom förut, upp över alla sina bräddar.
Det var på tionde dagen i första månaden som folket steg upp ur Jordan; och de lägrade sig i Gilgal, på gränsen av östra Jerikoområdet.
Och de tolv stenarna som de hade tagit ur Jordan reste Josua i Gilgal.
Och han sade till Israels barn: »När nu edra barn i framtiden fråga sina fäder: 'Vad betyda dessa stenar?',
då skolen I göra det kunnigt för edra barn och säga: 'Israel gick på torr mark över denna Jordan,
i det att HERREN, eder Gud, lät vattnet i Jordan torka ut framför eder, till dess I haden gått över den, likasom HERREN, eder Gud, gjorde med Röda havet, som han lät torka ut framför oss, till dess vi hade gått över det;
på det att alla folk på jorden må förnimma huru stark HERRENS hand är, så att I frukten HERREN, eder Gud, alltid.'»
Då nu alla amoréernas konungar på andra sidan Jordan, på västra sidan, och alla kananéernas konungar vid havet hörde huru HERREN hade låtit vattnet i Jordan torka ut framför Israels barn, medan vi gingo över den, blevo deras hjärtan förfärade, och de hade icke längre mod att stå emot Israels barn.
Vid den tiden sade HERREN till Josua: »Gör dig stenknivar och omskär åter Israels barn, för andra gången.»
Då gjorde Josua sig stenknivar och omskar Israels barn vid Förhudshöjden.
Och orsaken varför Josua omskar dem var denna: allt det folk av mankön, som hade dragit ut ur Egypten, alla stridbara män, hade dött i öknen under vägen, efter uttåget ur Egypten.
Ty väl hade bland folket alla de som voro med under uttåget blivit omskurna, men de bland folket, som voro födda i öknen under vägen, efter uttåget ur Egypten, de voro alla oomskurna.
Ty Israels barn vandrade i öknen i fyrtio år, under vilken tid alla stridbara män i folket, som hade dragit ut ur Egypten, förgingos, eftersom de icke hörde HERRENS röst, varför ock HERREN svor att han icke skulle låta dem se det land som han med ed hade lovat deras fäder att giva oss, ett land som flyter av mjölk och honung.
Men deras barn, som han hade låtit uppstå i deras ställe, dem omskar nu Josua, ty de hade förhud, eftersom de icke hade blivit omskurna under vägen.
Och när allt folket hade blivit omskuret, stannade de kvar där de voro i lägret, till dess de hade blivit läkta.
Och HERREN sade till Josua: »I dag har jag avvältrat från eder Egyptens smälek.»
Och detta ställe fick namnet Gilgal, såsom det heter ännu i dag.
Medan nu Israels barn voro lägrade i Gilgal, höllo de påskhögtid den fjortonde dagen i månaden, om aftonen, på Jerikos hedmarker.
Och dagen efter påskhögtiden åto de osyrat bröd och rostade ax av landets säd, just på den dagen.
Och mannat upphörde dagen därefter, då de nu åto av landets säd, och Israels barn fingo icke manna mer, utan de åto det året av landet Kanaans avkastning.
Och medan Josua var vid Jeriko, hände sig att han, i det han lyfte upp sina ögon, fick se en man stå där framför sig med ett draget svärd i sin hand.
Då gick Josua fram till honom och frågade honom: »Tillhör du oss eller våra ovänner?»
Han svarade: »Nej, jag är hövitsman över HERRENS här, och jag har just nu kommit hit.»
Då föll Josua ned till jorden på sitt ansikte och bugade sig; sedan sade han till honom: »Vad har min herre att säga till sin tjänare?»
Hövitsmannen över HERRENS här sade då till Josua: »Drag dina skor av dina fötter, ty platsen där du står är helig.»
Och Josua gjorde så.
Och Jeriko hade sina portar stängda, det höll sig tillstängt för Israels barn; ingen gick ut eller in.
Men HERREN sade till Josua: »Se, jag har givit Jeriko med dess konung, med dess tappra stridsmän, i din hand.
Tågen nu omkring staden, så många stridbara män I ären, runt omkring staden en gång; så skall du göra i sex dagar.
Och sju präster skola bära de sju jubelbasunerna framför arken; men på sjunde dagen skolen I tåga omkring staden sju gånger; och prästerna skola stöta i basunerna.
Och när det blåses i jubelhornet med utdragen ton, och I hören basunljudet, skall allt folket upphäva ett stort härskri; då skola stadsmurarna falla på stället, och folket skall draga in över dem, var och en rätt fram.»
Då kallade Josua, Nuns son, till sig prästerna och sade till dem: »Tagen förbundsarken, och sju präster skola bära sju jubelbasuner framför HERRENS ark.»
Och till folket blev sagt: »Dragen ut och tågen omkring staden; och den väpnade skaran skall draga framför HERRENS ark.»
Då nu Josua hade sagt detta till folket, drogo de sju präster som buro jubelbasunerna framför HERREN åstad och stötte i basunerna; och HERRENS förbundsark följde efter dem.
Och den väpnade skaran gick framför prästerna som stötte i basunerna, och den övriga hopen slutade tåget och följde efter arken, under det att man alltjämt stötte i basunerna.
Men Josua hade bjudit folket och sagt: »I skolen icke upphäva något härskri eller låta höra eder röst eller ens låta något ord utgå av eder mun, förrän den dag då jag säger till eder: 'Häven upp ett härskri'; då skolen I upphäva ett härskri.»
Och när han så hade låtit bära HERRENS ark omkring staden, runt omkring den en gång, gingo de in i lägret och stannade i lägret över natten.
Och följande morgon stod Josua bittida upp, och prästerna togo HERRENS ark.
Och de sju präster som buro de sju jubelbasunerna framför HERRENS ark gingo alltjämt och stötte i basunerna; och den väpnade skaran gick framför dem, och den övriga hopen slutade tåget och följde efter HERRENS ark, under det att man alltjämt stötte i basunerna.
De tågade också nu på andra dagen en gång omkring staden och återvände sedan till lägret; så gjorde de i sex dagar.
Men på sjunde dagen stodo de bittida upp vid morgonrodnadens uppgång och tågade då sju gånger omkring staden på samma sätt; endast denna dag tågade de sju gånger omkring staden.
Och när prästerna sjunde gången stötte i basunerna, sade Josua till folket: »Häven upp ett härskri, ty HERREN har givit eder staden.
Men staden med allt vad däri är skall givas till spillo åt HERREN; allenast skökan Rahab skall få leva, jämte alla som äro inne i hennes hus, därför att hon gömde de utskickade som vi hade sänt åstad.
Men tagen eder väl till vara för det tillspillogivna, så att I icke, sedan I haven givit det till spillo, ändå tagen något av det tillspillogivna och därigenom kommen Israels läger att hemfalla åt tillspillogivning, och så dragen olycka över det.
Allt silver och guld och allt som är av koppar eller järn skall vara helgat åt HERREN och ingå till HERRENS skatt.»
Då hov folket upp ett härskri, och man stötte i basunerna.
Ja, när folket hörde basunljudet, hov det upp ett stort härskri; då föllo murarna på stället, och folket drog över dem in i staden, var och en rätt fram; så intogo de staden.
Och de gåvo till spillo allt vad som fanns i staden, både män och kvinnor, både unga och gamla, så ock oxar, får och åsnor, och slogo dem med svärdsegg.
Men till de båda män som hade bespejat landet sade Josua: »Gån in i skökans hus och fören kvinnan, jämte alla som tillhöra henne, ut därifrån, såsom I med ed haven lovat henne.»
Då gingo de unga män som hade varit där såsom spejare ditin och förde ut Rahab, jämte hennes fader och moder och hennes bröder och alla som tillhörde henne; hela hennes släkt förde de ut.
Och de släppte dem utanför Israels läger.
Men staden med allt vad som fanns däri brände de upp i eld; allenast silvret och guldet och det som var av koppar eller järn lade de till skatten i HERRENS hus.
Men skökan Rahab och hennes faders hus och alla som tillhörde henne lät Josua leva, och hon fick bo bland Israels folk, intill denna dag; detta därför att hon gömde de utskickade som Josua hade sänt åstad för att bespeja Jeriko.
På den tiden lät Josua folket svärja denna ed: »Förbannad vare inför HERREN den man som tager sig före att åter bygga upp denna stad, Jeriko.
När han lägger dess grund, må detta kosta honom hans äldste son, och när han sätter upp dess portar, må detta kosta honom hans yngste son.»
Och HERREN var med Josua, så att ryktet om honom gick ut över hela landet.
Men Israels barn förgrepo sig trolöst på det tillspillogivna; ty Akan, son till Karmi, son till Sabdi, son till Sera, av Juda stam, tog något av det tillspillogivna.
Då upptändes HERRENS vrede mot Israels barn.
Och Josua sände från Jeriko några män åstad till Ai, som ligger vid Bet-Aven, öster om Betel, och sade till dem: »Dragen ditupp och bespejen landet.»
Så drogo då männen upp och bespejade Ai.
Och när de kommo tillbaka till Josua, sade de till honom: »Allt folket behöver icke draga ditupp; om vid pass två eller tre tusen man draga upp, skola de nog intaga Ai.
Du behöver icke låta allt folket göra sig mödan att tåga dit, ty dess invånare äro få.»
Alltså fingo vid pass tre tusen man av folket draga ditupp; men dessa måste fly för ajiterna.
Och sedan ajiterna hade slagit vid pass trettiosex man av dem, förföljde de de övriga utanför stadsporten ända till Sebarim och slogo dem på sluttningen där.
Då blev folkets hjärta förfärat, det blev såsom vatten.
Och Josua med de äldste i Israel rev sönder sina kläder, och föll ned på sitt ansikte till jorden framför HERRENS ark och låg där ända till aftonen, och de strödde stoft på sina huvuden.
Och Josua sade: »Ack, Herre, HERRE, varför har du då fört detta folk över Jordan, om du vill giva i amoréernas hand och så förgöra oss?
O att vi hade beslutit oss för att stanna på andra sidan Jordan!
Ack Herre, vad skall jag nu säga, sedan Israel har tagit till flykten för sina fiender?
När kananéerna och landets alla övriga inbyggare få höra detta, skola de omringa oss och utrota till och med vårt namn från jorden.
Vad vill du då göra för ditt stora namns ära?»
Men HERREN svarade Josua: »Stå upp.
Varför ligger du så på ditt ansikte?
Israel har syndat, de hava överträtt det förbund som jag stadgade för dem; de hava tagit av det tillspillogivna, de hava stulit, de hava ljugit, de hava gömt det bland sitt eget gods.
Därför kunna Israels barn icke stå emot sina fiender, utan de måste taga till flykten för sina fiender, ty de äro nu själva hemfallna åt tillspillogivning.
Jag vill icke mer vara med eder, om I icke alldeles skaffen bort ifrån eder det tillspillogivna.
Stå nu upp och helga folket och säg: Helgen eder till i morgon.
Ty så säger HERREN, Israels Gud: Något tillspillogivet finnes hos dig, Israel; du skall icke kunna stå emot dina fiender, förrän I skiljen det tillspillogivna från eder.
I morgon skolen I träda fram, den ena stammen efter den andra; i den stam som HERREN då låter träffas av lotten skall den ena släkten efter den andra träda fram; och i den släkt som HERREN låter träffas av lotten skall den ena familjen efter den andra träda fram; och i den familj som HERREN låter träffas av lotten skall den ena mannen efter den andra träda fram.
Och den som då träffas av lotten såsom skyldig till förgripelse på det tillspillogivna, han skall brännas upp i eld med allt vad han har, därför att han överträdde HERRENS förbund och gjorde vad som var en galenskap i Israel.»
Så lät nu Josua bittida följande morgon Israel träda fram, den ena stammen efter den andra; då träffades Juda stam av lotten.
När han då lät Juda släkter träda fram, träffade lotten seraiternas släkt; och när han lät seraiternas släkt träda fram, den ena mannen efter den andra, träffades Sabdi av lotten.
När han då lät hans familj träda fram, den ena mannen efter den andra, träffade lotten Akan, son till Karmi, son till Sabdi, son till Sera av Juda stam.
Då sade Josua till Akan: »Min son, giv ära åt HERREN, Israels Gud, och bekänn, honom till pris: säg mig vad du gjort och dölj intet för mig.»
Akan svarade Josua och sade: »Det är sant, jag har syndat mot HERREN, Israels Gud, ty så har jag gjort:
jag såg ibland bytet en dyrbar mantel från Sinear och två hundra siklar silver och en guldplatta, femtio siklar i vikt, och till detta fick begärelse och tog det; se, det är gömt i jorden, i mitten av mitt tält, och silvret underst.»
Då sände Josua några män dit för att se efter, och de skyndade till tältet; och de funno det gömt där i hans tält, och silvret underst.
Och de togo det ur tältet och buro det till Josua och Israels barns menighet och lade det ned inför HERREN.
Då tog Josua och Israels menighet med honom Akan, Seras son, och silvret och manteln och guldplattan, och hans söner och döttrar, hans oxar, åsnor och får, och hans tält, och allt övrigt som han hade, och förde alltsammans upp till Akors dal.
Och Josua sade: »Varför drog du olycka över oss?
Nu skall ock HERREN i dag låta olycka komma över dig.»
Och Israels menighet stenade honom; de brände upp dem i eld och kastade stenar på dem.
Och de uppkastade över honom ett stort stenröse, som finnes kvar ännu i dag; och så vände sig HERREN ifrån sin vredes glöd.
Därav fick det stället namnet Akors dal, såsom det heter ännu i dag.
Och HERREN sade till Josua: »Frukta icke och var icke förfärad; tag med dig allt krigsfolket och stå upp och drag åstad mot Ai.
Se, i din hand har jag givit konungen i Ai med hans folk, hans stad och hans land.
Och du skall göra med Ai och dess konung på samma sätt som du gjorde med Jeriko och dess konung; dock mån I behålla rovet därifrån och boskapen, såsom edert byte.
Lägg nu ett bakhåll mot staden, på andra sidan därom.»
Då bröt Josua upp med allt krigsfolket för att draga åstad mot Ai.
Och Josua utvalde trettio tusen man, de tappraste stridsmännen, och sände dem ut om natten.
Och han bjöd dem och sade: »Given akt: I skolen lägga eder i bakhåll mot staden, på andra sidan därom, men läggen eder icke alltför långt ifrån staden; och hållen eder alla redo.
Själv skall jag, med allt det folk som är kvar hos mig, rycka fram mot staden.
När de då draga ut mot oss såsom förra gången, vilja vi fly för dem.
Då skola de draga efter oss, till dess vi hava lockat dem långt bort ifrån staden; ty de skola tänka: 'De flyr för oss, nu såsom förra gången.'
Men under det att vi fly för dem, skolen I bryta fram ifrån bakhållet och intaga staden, ty HERREN, eder Gud, har givit den i eder hand.
Och så snart I haven fått staden i edert våld, skolen I tända eld på den; efter HERRENS ord skolen I så göra.
Given akt på vad jag nu har bjudit eder.»
Så sände Josua dem åstad, och de gingo och lade sig i bakhåll mellan Betel och Ai, väster om Ai.
Men Josua stannade över natten bland folket.
Och bittida följande morgon mönstrade Josua folket och drog så, med de äldste i Israel i spetsen för folket, upp till Ai.
Och allt det krigsfolk som var kvar hos honom drog med ditupp och ryckte allt närmare, till dess de kommo mitt emot staden; där lägrade de sig norr om Ai, med dalen mellan sig och Ai.
Men han tog vid pass fem tusen man och lade dem i bakhåll mellan Betel och Ai, väster om staden.
Och sedan folket hade blivit uppställt, såväl hela lägret, norr om staden, gick Josua den natten fram till mitten av dalen.
När konungen i Ai såg detta, skyndade sig männen i staden, han själv med allt sitt folk, och drogo bittida om morgonen ut till strid mot Israel, bort till den utsedda platsen, framför hedmarken; han själv visste nämligen icke att ett bakhåll var lagt mot honom på andra sidan om staden.
Och Josua och hela Israel läto slå sig av dem och flydde åt öknen till.
Då uppbådades allt folket i staden till att förfölja dem; och under det att de förföljde Josua, blevo de lockade långt bort ifrån staden.
Icke en enda man blev kvar i Ai eller i Betel, utan alla drogo ut efter Israel och lämnade staden öppen, i det att de förföljde Israel.
Och HERREN sade till Josua: »Räck ut lansen, som du har i din hand, mot Ai, ty jag skall giva det i din hand.»
Då räckte Josua ut lansen, som han hade i sin hand, mot staden.
Och de som lågo i bakhåll bröto med hast upp från sin plats och skyndade åstad, så snart han räckte ut sin hand, och kommo in i staden och intogo den; och de tände strax eld på staden.
När då männen från Ai vände sig om, fingo de se röken från staden stiga upp mot himmelen; och de hade ingen utväg att fly, vare sig hit eller dit, då nu det folk som flydde åt öknen vände sig mot sina förföljare.
Ty när Josua och hela Israel sågo att de som lågo i bakhåll hade intagit staden, och att röken steg upp från staden, vände de om och angrepo ajiterna.
De andra drogo nu också ut från staden emot dem, så att de kommo mitt emellan israeliterna och fingo dem på båda sidor om sig, och dessa nedgjorde dem då och läto ingen av dem slippa undan och rädda sig.
Men konungen i Ai blev levande tagen till fånga och förd till Josua.
Och när Israel hade dräpt alla Ais invånare ute på fältet, i öknen, dit de hade förföljt dem, och dessa allasammans så hade fallit för svärdsegg och blivit nedgjorda, då vände hela Israel tillbaka till Ai och slog med svärdsegg också dem som voro där.
Och de som föllo på den dagen, män och kvinnor, utgjorde tillsammans tolv tusen personer, allt folket i Ai.
Ty Josua drog icke tillbaka sin hand, med vilken han hade räckt ut lansen, förrän alla Ais invånare hade blivit givna till spillo.
Allenast boskapen och rovet från denna stad togo israeliterna såsom sitt byte, efter den befallning som HERREN hade givit Josua.
Och Josua brände upp Ai och gjorde det till en grushög för evärdlig tid, till en ödemark, såsom det är ännu i dag.
Och konungen i Ai lät han hänga upp på en påle, där han fick hänga ända till aftonen.
Men när solen gick ned, tog man på Josuas befallning hans döda kropp ned från pålen och kastade den vid ingången till stadsporten; och man uppkastade över den ett stort stenröse, som finnes kvar ännu i dag.
Då byggde Josua åt HERREN, Israels Gud, ett altare på berget Ebal,
såsom HERRENS tjänare Mose hade bjudit Israels barn, och såsom det var föreskrivet i Moses lagbok: ett altare av ohuggna stenar, vid vilka man icke hade kommit med något järn; och på det offrade de brännoffer åt HERREN och slaktade tackoffer.
Och han lät där på stenarna sätta en avskrift av Moses lag, den lag som Mose hade skrivit och förelagt Israels barn.
Och Israels menighet, med dess äldste och tillsyningsmän och domare, stod på båda sidor om arken, så att de hade framför sig de levitiska prästerna som buro HERRENS förbundsark, menigheten, främlingar såväl som infödingar, den ena hälften vänd mot berget Gerissim och den andra hälften mot berget Ebal, i enlighet med vad HERRENS tjänare Mose hade bjudit, nämligen att man först skulle välsigna Israels folk.
Därefter läste han upp alla lagens ord, välsignelsen och förbannelsen, alldeles såsom det var skrivet i lagboken.
Icke ett ord av allt det som Mose hade bjudit underlät Josua att uppläsa inför Israels hela församling, med kvinnor och barn, och inför de främlingar som följde med dem.
Då nu alla de konungar som bodde på andra sidan Jordan, i Bergsbygden, i Låglandet och i hela kustlandet vid Stora havet upp emot Libanon, hörde vad som hade skett -- hetiterna, amoréerna, kananéerna, perisséerna, hivéerna och jebuséerna --
slöto de sig endräktigt tillhopa för att strida mot Josua och Israel.
Men när invånarna i Gibeon hörde vad Josua hade gjort med Jeriko och Ai,
togo också de sin tillflykt till list: de gingo åstad och föregåvo sig vara sändebud; de lade utslitna packsäckar på sina åsnor, så ock utslitna, sönderspruckna och hopflickade vinläglar av skinn,
och togo utslitna, lappade skor på sina fötter och klädde sig i utslitna kläder, varjämte allt det bröd de togo med sig till reskost var torrt och söndersmulat.
Så gingo de till Josua i lägret vid Gilgal och sade till honom och Israels män: »Vi hava kommit hit från ett avlägset land; sluten nu förbund med oss.»
Men Israels män svarade hivéerna: »Kanhända bon I här mitt ibland oss; huru skulle vi då kunna sluta förbund med eder?»
Då sade de till Josua: »Vi vilja bliva dig underdåniga.»
Josua frågade dem: »Vilka ären I då, och varifrån kommen I?»
De svarade honom: »Dina tjänare hava kommit från ett mycket avlägset land för HERRENS, din Guds, namns skull; ty vi hava hört ryktet om honom och allt vad han har gjort i Egypten
och allt vad han har gjort med amoréernas konungar, de två på andra sidan Jordan, Sihon, konungen i Hesbon, och Og, konungen i Basan, som bodde i Astarot.
Därför sade våra äldste och alla vårt lands inbyggare till oss: 'Tagen reskost med eder och gån dem till mötes och sägen till dem: Vi vilja bliva eder underdåniga, sluten nu förbund med oss.'
Detta vårt bröd var nybakat, när vi togo det med oss till reskost hemifrån, den dag vi gåvo oss i väg för att gå till eder; men se, nu är det torrt och söndersmulat.
Dessa vinläglar, som voro nya, när vi fyllde dem, se, de äro nu sönderspruckna.
Och dessa kläder och skor som vi hava på oss hava blivit utslitna under vår mycket långa resa.»
Då togo männen av deras reskost, men rådfrågade icke HERRENS mun.
Och Josua tillförsäkrade dem fred och slöt ett förbund med dem, att de skulle få leva; och menighetens hövdingar gåvo dem sin ed.
Men när tre dagar voro förlidna, sedan de hade slutit förbund med dem, fingo de höra att de voro från grannskapet, ja, att de bodde mitt ibland dem.
Då bröto Israels barn upp och kommo på tredje dagen till deras städer; och deras städer voro: Gibeon, Kefira, Beerot och Kirjat-Jearim.
Likväl angrepo Israels barn dem icke, eftersom menighetens hövdingar hade givit dem sin ed vid HERREN, Israels Gud.
Men hela menigheten knorrade mot hövdingarna.
Då sade alla hövdingarna till menigheten: »Vi hava givit dem vår ed vid HERREN, Israels Gud; därför kunna vi nu icke komma vid dem.
Detta är vad vi vilja göra med dem, i det att vi låta dem leva, på det att icke förtörnelse må komma över oss, för edens skull som vi hava svurit dem.»
Och hövdingarna sade till dem att de skulle få leva; men de måste bliva vedhuggare och vattenbärare åt hela menigheten, såsom hövdingarna hade sagt till dem.
Och Josua kallade dem till sig och talade till dem och sade: »Varför haven I bedragit oss och sagt: 'Vi bo mycket långt borta från eder', fastän I bon mitt ibland oss?
Så varen I därför nu förbannade; I skolen aldrig upphöra att vara trälar, vedhuggare och vattenbärare vid min Guds hus.»
De svarade Josua och sade: »Det hade blivit berättat för dina tjänare huru HERREN, din Gud, hade tillsagt sin tjänare Mose att han ville giva eder hela detta land och förgöra alla landets inbyggare för eder; därför fruktade vi storligen för våra liv, när I kommen, och så gjorde vi detta.
Och se, nu äro vi i din hand.
Vad dig synes gott och rätt att göra med oss, det må du göra.»
Och han gjorde så med dem; han friade dem från Israels barns hand, så att de icke dräpte dem;
men tillika bestämde Josua på den dagen att de skulle bliva vedhuggare och vattenbärare och vid HERRENS altare -- såsom de äro ännu i dag -- på den plats som han skulle utvälja.
Då nu Adoni-Sedek, konungen i Jerusalem, hörde att Josua hade intagit Ai och givit det till spillo, och att han hade gjort med Ai och dess konung på samma sätt som han hade gjort med Jeriko och dess konung, och att invånarna i Gibeon hade ingått fred med Israel och fingo bo mitt ibland dem,
fruktade han och hans folk storligen, ty Gibeon var en stor stad, såsom en av konungastäderna, ja, det var större än Ai, och dess män voro alla tappra.
Och Adoni-Sedek, konungen i Jerusalem, sände till Hoham, konungen i Hebron, till Piram, konungen i Jarmut, till Jafia, konungen i Lakis, och till Debir, konungen i Eglon, och lät säga:
»Kommen hitupp till mig och hjälpen mig, så att vi kunna slå gibeoniterna, ty de hava ingått fred med Josua och Israels barn.»
Så församlade sig då de fem amoreiska konungarna, konungen i Jerusalem, konungen i Hebron, konungen i Jarmut, konungen i Lakis, konungen i Eglon, och drogo ditupp med alla sina härar; och de belägrade Gibeon och angrepo det.
Men gibeoniterna sände till Josua i lägret vid Gilgal och läto säga: »Drag icke din hand från dina tjänare, utan kom hitupp till oss med hast och undsätt oss och hjälp oss, ty konungarna över amoréerna, som bo i bergsbygden, hava församlat sig mot oss.»
Då drog Josua ditupp från Gilgal med allt sitt krigsfolk och alla sina tappraste stridsmän.
Och HERREN sade till Josua: »Frukta icke för dem, ty jag har givit dem i dina händer; ingen av dem skall kunna stå dig emot.»
Och Josua kom plötsligt över dem, ty han tågade hela natten, sedan han hade brutit upp från Gilgal.
Och HERREN sände en sådan förvirring bland dem, när de fingo se israeliterna, att dessa tillfogade dem ett stort nederlag vid Gibeon; därefter förföljde de dem på vägen upp till Bet-Horon och nedgjorde dem, och drevo dem ända till Aseka och Mackeda.
Och när de så, under sin flykt för Israel, hade kommit till den sluttning som går ned från Bet-Horon, lät HERREN stora stenar falla över dem från himmelen, hela vägen ända till Aseka, så att de blevo dödade; de som dödades genom hagelstenarna voro till och med flera än de som Israels barn dräpte med svärd.
Och Josua talade till HERREN på den dag då HERREN gav amoréerna i Israels barns våld; han sade inför Israel: »Du sol, stå stilla i Gibeon, du måne, i Ajalons dal!»
Då stod solen stilla, och månen blev stående, till dess folket hade tagit hämnd på sina fiender.
Detta finnes ju upptecknat i »Den redliges bok».
Solen blev stående mitt på himmelen nästan en hel dag och hastade icke att gå ned.
Aldrig har någon dag, varken förr eller senare, varit lik denna, i det att HERREN då lydde en mans ord; ty HERREN stridde för Israel.
Och Josua med hela Israel vände tillbaka till lägret vid Gilgal.
Men de fem konungarna flydde och gömde sig i grottan vid Mackeda.
Då blev det inberättat för Josua: »Man har funnit de fem konungarna gömda i grottan till Mackeda.»
Josua sade: »Vältren stora stenar framför ingången till grottan, och sätten dit folk för att bevaka den.
Men I andra, stannen icke, utan förföljen edra fiender, och nedgören dem som bliva efter; låten dem icke komma in i sina städer, ty HERREN, eder Gud har givit dem i eder hand.»
Då nu Josua och Israels barn hade tillfogat dem ett mycket stort nederlag och nedgjort dem -- varvid dock några av dem lyckades rädda sig och komma in i de befästa städerna --
vände allt folket välbehållet tillbaka till Josua i lägret vid Mackeda, ty ingen vågade mer ens röra sin tunga mot någon av Israels barn.
Då sade Josua: »Öppnen grottan och fören de fem konungarna till mig, ut ur grottan.»
De gjorde så och förde de fem konungarna ut till honom ur grottan: konungen i Jerusalem, konungen i Hebron, konungen i Jarmut, konungen i Lakis, och konungen i Eglon.
När dessa konungar hade blivit förda ut till Josua, kallade Josua till sig alla Israels män och sade till anförarna för krigsfolket som hade dragit med honom: »Träden fram och sätt edra fötter på dessa konungars halsar.»
Och de trädde fram och satte sina fötter på deras halsar.
Sedan sade Josua till dem: »Frukten icke och varen icke försagda, utan varen frimodiga och oförfärade, ty så skall HERREN göra med alla sina fiender som I kommen i strid med.»
Därefter lät Josua slå dem till döds och hänga upp dem på fem pålar; och de fingo på pålarna ända till aftonen.
Men vid solnedgången togos de på Josuas befallning ned från pålarna och kastades in i grottan där de hade varit gömda; och framför ingången till grottan lade man stora stenar, som ligga kvar där ännu i denna dag.
Och Josua intog Mackeda på den dagen och slog dess invånare och dess konung med svärdsegg; han gav det till spillo med alla dem som voro därinne och lät ingen slippa undan.
Och han gjorde med konungen i Mackeda på samma sätt som han hade gjort med konungen i Jeriko.
Därefter drog Josua med hela Israel från Mackeda till Libna och belägrade Libna.
Och HERREN gav också det och dess konung i Israels hand; och de slogo dess invånare med svärdsegg, alla dem som voro därinne, och läto ingen därinne slippa undan.
Och han gjorde med dess konung på samma sätt som han hade gjort med konungen i Jeriko.
Sedan drog Josua med hela Israel från Libna till Lakis och belägrade och angrep det.
Och HERREN gav Lakis i Israels hand, så att de intogo det på andra dagen; och de slogo dess invånare med svärdsegg, alla dem som voro därinne -- alldeles såsom de hade gjort med Libna.
Då drog Horam, konungen i Geser, upp för att hjälpa Lakis; men Josua slog honom och hans folk och lät ingen av dem slippa undan.
Och från Lakis drog Josua med hela Israel till Eglon, och de belägrade och angrepo det.
Och de intogo det samma dag och slogo dess invånare med svärdsegg, och han gav på den dagen till spillo alla dem som voro därinne -- alldeles såsom han hade gjort med Lakis.
Sedan drog Josua med hela Israel från Eglon upp till Hebron och belägrade det.
Och de intogo det och slogo dess invånare och dess konung med svärdsegg, så ock alla dess lydstäder och alla dem som voro därinne, och han lät ingen slippa undan -- alldeles såsom han hade gjort med Eglon.
Han gav det till spillo med alla dem som voro därinne.
Därefter vände Josua med hela Israel tillbaka till Debir och belägrade det.
Och han underkuvade det med dess konung och alla dess lydstäder, och de slogo deras invånare med svärdsegg; de gåvo till spillo alla dem som voro därinne, och han lät ingen slippa undan.
Han gjorde med Debir och dess konung på samma sätt som han hade gjort med Hebron, och såsom han hade gjort med Libna och dess konung.
Så intog Josua hela landet, Bergsbygden, Sydlandet, Låglandet och Bergssluttningarna, och slog alla konungar där och lät ingen slippa undan; han gav till spillo allt vad andra hade, såsom HERREN, Israels Gud, hade bjudit.
Josua intog allt som fanns mellan Kades-Barnea och Gasa, så ock hela landet Gosen ända till Gibeon.
Alla dessa konungar och deras land underkuvade Josua på en gång, ty HERREN, Israels Gud, stridde för Israel.
Därefter vände Josua med hela Israel tillbaka till lägret vid Gilgal.
Då nu Jabin, konungen i Hasor, hörde detta, sände han bud till Jobab, konungen i Madon, och till konungen i Simron och konungen i Aksaf
och till de konungar som bodde norrut, i Bergsbygden och på Hedmarken, söder om Kinarot, och i Låglandet, så ock i Nafot-Dor, västerut,
vidare till kananéerna österut och västerut och till amoréerna, hetiterna, perisséerna och jebuséerna i Bergsbygden, så och till hivéerna nedanför Hermon, i Mispalandet.
Dessa drogo nu ut med alla sina härar, en folkskara så talrik som sanden på havets strand, jämte hästar och vagnar i stor myckenhet.
Alla dessa konungar rotade sig samman; och de kommo och lägrade sig tillhopa vid Meroms vatten, för att strida mot Israel.
Men HERREN sade till Josua: »Frukta icke för dem, ty i morgon vid denna tid vill jag själv giva dem allasammans slagna i Israels våld.
På deras hästar skall du avskära fotsenorna, och deras vagnar skall du bränna upp i eld.»
Och Josua kom med allt sitt krigsfolk plötsligt över dem vid Meroms vatten och anföll dem.
Och HERREN gav dem i Israels hand, och de slogo dem och förföljde dem ända till Stora Sidon, till Misrefot-Maim och till Mispedalen, österut; de slogo dem och läto ingen slippa undan.
Och Josua gjorde med dem såsom HERREN hade befallt honom: på deras hästar lät han avskära fotsenorna, och deras vagnar lät han bränna upp i eld.
Därefter, vid samma tid, vände Josua tillbaka och intog Hasor och slog dess konung med svärd; ty Hasor var fordom huvudstaden för alla dessa riken.
Alla de som voro därinne blevo slagna med svärdsegg och givna till spillo, så att intet som anda hade lämnades kvar; och själva Hasor brände han upp i eld.
Likaledes underkuvade Josua alla de andra konungastäderna med alla deras konungar, och han slog deras invånare med svärdsegg och gav dem till spillo, såsom HERRENS tjänare Mose hade bjudit.
Dock brände Israel icke upp någon av de städer som lågo på höjder, utom Hasor allena, ty det uppbrändes av Josua.
Och allt rovet från dessa städer, så ock boskapen, togo Israels barn såsom sitt byte; men alla människor i dem slogo de med svärdsegg, till dess att de hade förgjort dem; de läto intet som anda hade bliva kvar.
Såsom HERREN hade bjudit sin tjänare Mose, så hade Mose bjudit Josua, och så gjorde Josua; han underlät icke något av allt det som HERREN hade bjudit Mose.
Så intog Josua hela detta land: Bergsbygden, hela Sydlandet och hela landet Gosen, Låglandet och Hedmarken, så ock Israels bergsbygd och dess lågland,
landet från Halakberget, som höjer sig mot Seir, ända till Baal-Gad i Libanonsdalen nedanför berget Hermon; och alla konungar där tog han till fånga och slog dem till döds.
I lång tid förde Josua krig mot alla dessa konungar.
Om man undantager de hivéer som bodde i Gibeon, fanns ingen stad som ingick fred med Israels barn, utan dessa intogo dem alla med strid.
Ty från HERREN kom det att de förstockade sina hjärtan och mötte Israel med krig, för att de skulle givas till spillo, och för att nåd icke skulle vederfaras dem; i stället skulle de förgöras, såsom HERREN hade bjudit Mose.
Under denna tid drog Josua åstad och utrotade anakiterna i Bergsbygden, i Hebron, Debir och Anab, i hela Juda bergsbygd och i hela Israels bergsbygd; Josua gav dem med deras städer till spillo.
I Israels barns land lämnades inga anakiter kvar; allenast i Gasa, Gat och Asdod blevo några kvar.
Så intog Josua hela landet, alldeles såsom HERREN hade lovat Mose; och Josua gav det till arvedel åt Israel, efter deras avdelningar och stammar.
Och landet hade nu ro från krig.
Dessa voro de konungar i landet, som Israels barn slogo, och vilkas land de togo i besittning på andra sidan Jordan, på östra sidan, landet från bäcken Arnon ända till berget Hermon, så ock hela Hedmarken på östra sidan:
Sihon, amoréernas konung, som bodde i Hesbon och rådde över landet Aroer vid bäcken Arnons strand och från dalens mitt, samt över ena hälften av Gilead ända till bäcken Jabbok, som är Ammons barns gräns,
ävensom över Hedmarken ända upp till Kinarotsjön, på östra sidan, och ända ned till Hedmarkshavet, Salthavet, på östra sidan, åt Bet-Hajesimot till, och längre söderut till trakten nedanför Pisgas sluttningar.
Vidare intogo de Ogs område, konungens i Basan, vilken var en av de sista rafaéerna och bodde i Astarot och Edrei.
Han rådde över Hermons bergsbygd och över Salka och hela Basan ända till gesuréernas och maakatéernas område, så ock över andra hälften av Gilead, till Sihons område, konungens i Hesbon.
HERRENS tjänare Mose och Israels barn hade slagit dessa; och HERRENS tjänare Mose hade givit landet till besittning åt rubeniterna, gaditerna och ena hälften av Manasse stam.
Och följande voro de konungar i landet, som Josua och Israels barn slogo på andra sidan Jordan, på västra sidan, från Baal-Gad i Libanonsdalen ända till Halakberget, som höjer sig mot Seir.
(Josua gav sedan landet till besittning åt Israels stammar, efter deras avdelningar,
såväl Bergsbygden, Låglandet, Hedmarken och Bergssluttningarna som ock Öknen och Sydlandet, hetiternas, amoréernas, kananéernas, perisséernas, hivéernas och jebuséernas land.)
De voro: konungen i Jeriko en, konungen i Ai, som ligger bredvid Betel, en,
konungen i Jerusalem en, konungen i Hebron en,
konungen i Jarmut en, konungen i Lakis en,
konungen i Eglon en, konungen i Geser en,
konungen i Debir en, konungen i Geder en,
konungen i Horma en, konungen i Arad en,
konungen i Libna en, konungen i Adullam en,
konungen i Mackeda en, konungen i Betel en,
konungen i Tappua en, konungen i Hefer en,
konungen i Afek en, konungen i Lassaron en,
konungen i Madon en, konungen i Hasor en,
konungen i Simron-Meron en, konungen i Aksaf en,
konungen i Taanak en, konungen i Megiddo en,
konungen i Kedes en, konungen i Jokneam vid Karmel en,
konungen över Dor i Nafat-Dor en, konungen över Goim vid Gilgal en,
konungen i Tirsa en -- tillsammans trettioen konungar.
Då nu Josua var gammal och kommen till hög ålder, sade HERREN till honom: »Du är gammal och kommen till hög ålder, men ännu återstår av landet en mycket stor del som skall intagas.
Detta är nämligen vad som återstår av landet: alla filistéernas kretsar och hela gesuréernas land.
Ty allt som finnes mellan Sihor, öster om Egypten, och Ekrons område norrut räknas till Kananéernas land, nämligen vad filistéernas fem hövdingar innehava -- den i Gasa, den i Asdod, den i Askelon, den i Gat och den i Ekron -- så ock avéernas område,
hela kananéernas land söderut, vidare Meara, som tillhör sidonierna, ända till Afek, ända till amoréernas område.
och gebaléernas land samt hela Libanonstrakten österut, från Baal-Gad, nedanför berget Hermon, ända dit där vägen går till Hamat --
alla inbyggarna i bergsbygden, från Libanon ända till Misrefot-Maim, alla sidonier: dessa skall jag själv fördriva för Israels barn.
Men fördela du genom lottkastning landet åt Israel till arvedel, såsom jag har bjudit dig.
Ja, redan nu må du utskifta detta land till arvedel åt de nio stammarna och åt ena hälften av Manasse stam.»
Jämte Manasse hade ock rubeniterna och gaditerna fått sin arvedel, den som Mose gav dem på andra sidan Jordan, på östra sidan, just såsom HERRENS tjänare Mose gav den åt dem:
landet från Aroer, vid bäcken Arnons strand, och från staden i dalens mitt, så ock hela Medebaslätten ända till Dibon,
jämte alla övriga städer som hade tillhört Sihon, amoréernas konung, vilken regerade i Hesbon, ända till Ammons barns område,
vidare Gilead och gesuréernas och maakatéernas område och hela Hermons bergsbygd och hela Basan ända till Salka,
hela Ogs rike i Basan, hans som regerade i Astarot och Edrei, och som levde kvar såsom en av de sista rafaéerna, sedan Mose hade slagit och fördrivit dem.
Dock fördrevo Israels barn icke gesuréerna och maakatéerna; därför bodde ock gesuréer och maakatéer kvar bland Israels folk, såsom de göra ännu i dag.
(Men åt Levi stam gav han icke någon arvedel.
HERRENS, Israels Guds, eldsoffer äro hans arvedel, såsom han har sagt honom.)
Mose gav alltså land åt Rubens barns stam, efter deras släkter.
De fingo området från Aroer, vid bäcken Arnons strand, och från staden i dalens mitt, så ock hela slätten vid Medeba,
Hesbon med alla dess lydstäder på slätten, Dibon, Bamot-Baal, Bet-Baal-Meon,
Jahas, Kedemot, Mefaat,
Kirjataim, Sibma, Seret-Hassahar på Dalberget,
Bet-Peor samt Pisgas sluttningar och Bet-Hajesimot,
alla städerna på slätten, hela Sihons rike, amoréernas konungs, hans som regerade i Hesbon, och som hade blivit slagen av Mose jämte de midjanitiska hövdingarna Evi, Rekem, Sur, Hur och Reba, Sihons lydfurstar, som bodde där i landet.
Bileam, Beors son, spåmannen, dräptes ock av Israels barn med svärd, jämte andra som då blevo slagna av dem.
Och gränsen för Rubens barn var Jordan; den utgjorde gränsen.
Detta är Rubens barns arvedel, efter deras släkter, städerna med sina byar.
Likaledes gav Mose land åt Gads stam, åt Gads barn, efter deras släkter.
De fingo till sitt område Jaeser och alla städer i Gilead och hälften av Ammons barns land, ända till det Aroer som ligger gent emot Rabba,
vidare landet från Hesbon ända till Ramat-Hammispe och Betonim, och från Mahanaim ända till Lidebirs område,
samt i dalen: Bet-Haram, Bet-Nimra, Suckot och Safon, det övriga av Sihons rike, konungens i Hesbon, intill Jordan, som utgjorde gränsen, upp till ändan av Kinneretsjön, landet på andra sidan Jordan, på östra sidan.
Detta är Gads barns arvedel, efter deras släkter, städerna med sina byar.
Och Mose gav också land åt ena hälften av Manasse stam, så att denna hälft av Manasse barns stam fick land, efter sina släkter.
Deras område utgjordes av landet från Mahanaim, av hela Basan, hela Ogs rike, konungens i Basan, med alla Jairs byar i Basan, sextio städer,
alltså ock av halva Gilead jämte Astarot och Edrei, Ogs huvudstäder i Basan; detta gavs åt Makirs, Manasses sons, barn, nämligen åt ena hälften av Makirs barn, efter deras släkter.
Dessa voro de arvslotter som Mose utskiftade på Moabs hedar, på andra sidan Jordan mitt emot Jeriko, på östra sidan.
Men åt Levi stam gav Mose icke någon arvedel.
HERREN, Israels Gud, är deras arvedel, såsom han har sagt dem.
Och dessa äro de arvslotter som Israels barn fingo i Kanaans land, de som prästen Eleasar och Josua, Nuns son, och huvudmännen för familjerna inom Israels barns stammar utskiftade åt dem,
nämligen genom lottkastning om vars och ens arvedel, såsom HERREN hade bjudit genom Mose angående de nio stammarna och den ena halva stammen.
Ty de två övriga stammarna och den andra halva stammen hade av Mose fått sin arvedel på andra sidan Jordan, men leviterna hade han icke givit någon arvedel bland dem.
Ty Josefs barn utgjorde två stammar, Manasse och Efraim; och åt leviterna gav man icke någon särskild del av landet, utan allenast några städer att bo i, med tillhörande utmarker för deras boskap och deras övriga egendom.
Såsom HERREN hade bjudit Mose, så gjorde Israels barn, när de utskiftade landet
Men Juda barn trädde fram inför Josua i Gilgal, och kenaséen Kaleb, Jefunnes son, sade till honom: »Du vet själv vad HERREN sade till gudsmannen Mose angående mig och dig i Kades-Barnea.
Jag var fyrtio år gammal, när HERRENS tjänare Mose sände mig åstad från Kades-Barnea för att bespeja landet, och jag avgav sedan min berättelse därom inför honom efter bästa förstånd.
Mina bröder, som hade varit däruppe med mig, gjorde folkets hjärtan försagda, men jag efterföljde i allt HERREN, min Gud.
Då betygade Mose på den dagen med ed och sade: 'Sannerligen, det land som din fot har beträtt skall vara din och dina barns arvedel för evärdlig tid, därför att du i allt har efterföljt HERREN, min Gud.'
Och se, nu har HERREN låtit mig leva, såsom han lovade, i ytterligare fyrtiofem år, sedan HERREN talade så till Mose -- de år Israel vandrade i öknen; se, jag är nu åttiofem år gammal.
Ännu i dag är jag lika stark som jag var den dag då Mose sände mig åstad, ja, sådan min kraft då var, sådan är den ännu, vare sig det gäller att strida eller att vara ledare och anförare.
Så giv mig nu denna bergsbygd om vilken HERREN talade på den dagen.
Du hörde ju själv då att anakiterna bo där, och att där finnas stora befästa städer; måhända är HERREN med mig, så att jag kan fördriva dem, såsom HERREN har lovat.»
Då välsignade Josua Kaleb, Jefunnes son, och gav honom Hebron till arvedel.
Alltså fick då kenaséen Kaleb, Jefunnes son, Hebron till arvedel, såsom det är ännu i dag, därför att han i allt hade efterföljt HERREN, Israels Gud.
Men Hebron hette fordom Kirjat-Arba efter den störste mannen bland anakiterna.
Och landet hade nu ro från krig.
Juda barns stam fick, efter sina släkter, sin lott söderut intill Edoms gräns, intill öknen Sin, längst ned i söder.
Och deras södra gräns begynte vid ändan av Salthavet, vid dess sydligaste vik,
gick vidare söder om Skorpionhöjden och fram till Sin, drog sig så upp söder om Kades-Barnea, gick därefter framom Hesron och drog sig upp till Addar samt böjde sig sedan mot Karka.
Vidare gick den fram till Asmon och därifrån ut till Egyptens bäck; sedan gick gränsen ut vid havet. »Detta», sade han, »skall vara eder gräns i söder.»
Gränsen i öster var Salthavet ända till Jordans utlopp.
Och gränsen på norra sidan begynte vid den vik av detta hav, där Jordan har sitt utlopp.
Därifrån drog sig gränsen upp mot Bet-Hogla och gick fram norr om Bet-Haaraba; vidare drog sig gränsen upp till Bohans, Rubens sons, sten.
Därefter drog sig gränsen upp till Debir från Akors dal i nordlig riktning mot det Gilgal som ligger mitt emot Adummimshöjden, söder om bäcken; sedan gick gränsen fram till Semeskällans vatten och så ut till Rogelskällan.
Vidare drog sig gränsen uppåt Hinnoms sons dal, söder om Jebus' höjd, det är Jerusalem; därefter drog sig gränsen upp till toppen av det berg som ligger gent emot Hinnomsdalen, västerut, i norra ändan av Refaimsdalen.
Och från toppen av detta berg drog sig gränsen fram till Neftoavattnets källa och vidare till städerna i Efrons bergsbygd; sedan drog sig gränsen till Baala, det är Kirjat-Jearim.
Och från Baala böjde sig gränsen åt väster mot Seirs bergsbygd och gick fram till Jearims bergshöjd, det är Kesalon, norr om denna, och gick så ned till Bet-Semes och framom Timna.
Vidare gick gränsen till Ekrons höjd, norrut; därefter drog sig gränsen till Sickeron, gick så framom berget Baala och därifrån ut till Jabneel; sedan gick gränsen ut vid havet.
Och gränsen i väster följde Stora havet; det utgjorde gränsen.
Dessa voro Juda barns gränser runt omkring, efter deras släkter.
Men åt Kaleb, Jefunnes son, gavs, efter HERRENS befallning till Josua, en särskild del bland Juda barn, nämligen Arbas, Anaks faders, stad, det är Hebron.
Och Kaleb fördrev därifrån Anaks tre söner, Sesai, Ahiman och Talmai, Anaks avkomlingar.
Därifrån drog han upp mot Debirs invånare.
Men Debir hette fordom Kirjat-Sefer.
Och Kaleb sade: »Åt den som angriper Kirjat-Sefer och intager det vill jag giva min dotter Aksa till hustru.»
När då Otniel, son till Kenas, Kalebs broder, intog det, gav han honom sin dotter Aksa till hustru.
Och när hon kom till honom, intalade hon honom att begära ett stycke åkermark av hennes fader; och hon steg hastigt ned från åsnan.
Då sade Kaleb till henne: »Vad önskar du?»
Hon sade: »Giv mig en avskedsskänk; eftersom du har gift bort mig till det torra Sydlandet, må du giva mig vattenkällor.»
Då gav han henne Illiotkällorna och Tatiotkällorna.
Detta var nu Juda barns stams arvedel, efter deras släkter.
Och de städer som lågo ytterst i Juda barns stam, mot Edoms gräns, i Sydlandet, voro: Kabseel, Eder, Jagur,
Kina, Dimona, Adada,
Kedes, Hasor och Jitnan,
Sif, Telem, Bealot,
Hasor-Hadatta, Keriot, Hesron, det är Hasor,
Amam, Sema, Molada,
Hasar-Gadda, Hesmon, Bet-Pelet,
Hasar-Sual, Beer-Seba och Bisjotja,
Baala, Ijim, Esem,
Eltolad, Kesil, Horma,
Siklag, Madmanna, Sansanna,
Lebaot, Silhim, Ain och Rimmon -- tillsammans tjugunio städer med sina byar.
I Låglandet: Estaol, Sorga, Asna,
Sanoa och En-Gannim, Tappua och Enam,
Jarmut och Adullam, Soko och Aseka,
Saaraim, Aditaim, Gedera och Gederotaim -- fjorton städer med sina byar;
Senan, Hadasa, Migdal-Gad,
Dilean, Mispe, Jokteel,
Lakis, Boskat, Eglon,
Kabbon, Lamas, Kitlis,
Gederot, Bet-Dagon, Naama och Mackeda -- sexton städer med sina byar;
Libna, Eter, Asan,
Jifta, Asna, Nesib,
Kegila, Aksib och Maresa -- nio städer med sina byar;
Ekron med underlydande städer och byar;
från Ekron till havet allt vad som ligger på sidan om Asdod samt dithörande byar;
vidare Asdod med underlydande städer och byar, Gasa med underlydande städer och byar ända till Egyptens bäck och fram till Stora havet, som utgjorde gränsen.
Och i Bergsbygden: Samir, Jattir, Soko,
Danna, Kirjat-Sanna, det är Debir,
Anab, Estemo, Anim,
Gosen, Holon och Gilo -- elva städer med sina byar;
Arab, Ruma, Esean,
Janum, Bet-Tappua, Afeka,
Humta, Kirjat-Arba, det är Hebron, och Sior -- nio städer med sina byar;
Maon, Karmel, Sif, Juta,
Jisreel, Jokdeam och Sanoa,
Kain, Gibea och Timna -- tio städer med sina byar;
Halhul, Bet-Sur, Gedor,
Maarat, Bet-Anot och Eltekon -- sex städer med sina byar;
Kirjat-Baal, det är Kirjat-Jearim, och Rabba -- två städer med sina byar;
I Öknen: Bet-Haaraba, Middin, Sekaka,
Nibsan, Ir-Hammela och En-Gedi -- sex städer med sina byar.
Men jebuséerna, som bodde i Jerusalem, kunde Juda barn icke fördriva; därför bodde ock jebuséerna kvar bland Juda barn i Jerusalem, såsom de göra ännu i dag.
Och lotten föll ut för Josefs barn sålunda: Landet från Jordan vid Jeriko till Jerikos vatten österut, öknen, som från Jeriko höjer sig uppåt Bergsbygden mot Betel.
Och gränsen gick vidare från Betel till Lus och så fram till arkiternas område, mot Atarot.
Därefter gick den västerut ned till jafletiternas område, ända till Nedre Bet-Horons område och till Geser; sedan gick den ut vid havet.
Detta fingo nu Josefs barn, Manasse och Efraim, till arvedel.
Efraims barn fingo, efter sina släkter, sina gränser sålunda: Gränsen för deras arvedel i öster gick från Atrot-Addar ända till Övre Bet-Horon.
Sedan gick gränsen ut vid havet.
I norr var Mikmetat gräns.
Därifrån böjde sig gränsen österut till Taanat-Silo.
Därefter gick den fram där i öster till Janoa.
Från Janoa gick den ned till Atarot och Naara, träffade så Jeriko och gick ut vid Jordan.
Från Tappua gick gränsen västerut till Kanabäcken och gick sedan ut vid havet.
Detta var Efraims barns stams arvedel, efter deras släkter.
Dit hörde ock de städer som avsöndrades åt Efraims barn inom Manasse barns arvedel, alla dessa städer med sina byar.
Men de fördrevo icke kananéerna som bodde i Geser; därför bodde ock kananéerna kvar bland Efraims barn, såsom de göra ännu i dag, men de blevo arbetspliktiga tjänare under dem.
Och Manasse stam fick sin lott sålunda, ty han var Josefs förstfödde: Makir, Manasses förstfödde, Gileads fader, fick Gilead och Basan, ty han var en stridsman.
Manasses övriga barn fingo ock land, efter sina släkter: Abiesers barn, Heleks barn, Asriels barn, Sikems barn, Hefers barn, och Semidas barn.
Dessa voro Manasses, Josefs sons, manliga avkomlingar, efter deras släkter.
Men Selofhad, son till Hefer, son till Gilead, son till Makir, son till Manasse, hade inga söner, utan allenast döttrar; och hans döttrar hette Mahela, Noa, Hogla, Milka och Tirsa.
Dessa trädde fram inför prästen Eleasar och Josua, Nuns son, och stamhövdingarna och sade: »HERREN bjöd Mose att giva oss en arvedel bland våra bröder.»
Då gav man dem, efter HERRENS befallning, en arvedel bland deras faders bröder.
Alltså blevo de lotter som tillföllo Manasse tio -- förutom Gileads land och Basan på andra sidan Jordan --
eftersom Manasses döttrar fingo en arvedel bland hans söner.
Men Gileads land hade Manasses övriga barn fått.
Och Manasse fick sin gräns bestämd sålunda: Den gick från Aser till Mikmetat, som ligger gent emot Sikem; därefter gick gränsen åt höger, till En-Tappuas inbyggare.
(Tappuas land tillföll nämligen Manasse, men själva Tappua, inemot Manasse gräns, tillföll Efraims barn.)
Och gränsen gick vidare ned till Kanabäcken, söder om bäcken; men städerna där tillföllo Efraim, fastän de lågo bland Manasse städer.
Manasse gräns gick vidare norr om bäcken och gick sedan ut vid havet.
Det som låg söder om den tillföll Efraim, men det som låg norr om den tillföll Manasse, och deras gräns var havet; och i norr nådde de till Aser och i öster till Isaskar.
Och inom Isaskar och Aser fick Manasse Bet-Sean med underlydande orter, Jibleam med underlydande orter, invånarna i Dor och underlydande orter, invånarna i En-Dor och underlydande orter, invånarna i Taanak och underlydande orter, invånarna i Megiddo och underlydande orter, de tre höjdernas land.
Men Manasse barn kunde icke intaga dessa städer, utan kananéerna förmådde hålla sig kvar där i landet.
När sedan Israels barn blevo de starkare, gjorde de kananéerna arbetspliktiga under sig; de fördrevo dem icke heller då.
Och Josefs barn talade till Josua och sade: »Varför har du givit oss till arvedel allenast en lott och ett skifte, fastän vi äro ett talrikt folk, då ju HERREN hitintills har välsignat oss?»
Då svarade Josua dem: »Om du är ett för talrikt folk, så drag upp till skogsbygden och röj dig där mark i perisséernas och rafaéernas land, eftersom Efraims bergsbygd är dig för trång.»
Men Josefs barn sade: »I bergsbygden finnes icke rum nog för oss; och de kananéer som bo i dalbygden hava allasammans stridsvagnar av järn, både de som bo i Bet-Sean och underlydande orter och de som bo i Jisreels dal.»
Josua sade till Josefs hus, till Efraim och Manasse: »Du är ett talrikt folk och har stor kraft, därför skall du icke hava allenast en lott;
utan du skall få en bergsbygd, som ju ock är en skogsbygd, men som du skall röja upp, så att till och med utkanterna därav skola tillhöra dig.
Ty du måste fördriva kananéerna, eftersom de hava stridsvagnar av järn och äro så starka.»
Och Israels barns hela menighet församlade sig i Silo och uppsatte där uppenbarelsetältet, då nu landet var dem underdånigt.
Men ännu återstodo av Israels barn sju stammar som icke hade fått sin arvedel sig tillskiftad.
Därför sade Josua till Israels barn: »Huru länge viljen I försumma att gå åstad och taga i besittning det land som HERREN, edra fäders Gud, har givit eder?
Utsen åt eder tre män för var stam, så skall jag sända dem åstad, för att de må stå upp och draga omkring i landet och sätta upp en beskrivning däröver, efter som vars och ens arvedel skall bliva, och så komma tillbaka till mig.
De skola nämligen uppdela det åt sig i sju delar, varvid Juda skall förbliva vid sitt område i söder och Josefs hus förbliva vid sitt område i norr.
Och sedan skolen I sätta upp beskrivningen över landet, efter dessa sju delar, och bära den hit till mig, så vill jag kasta lott för eder här inför HERREN, vår Gud.
Ty leviterna få ingen särskild del bland eder, utan HERRENS prästadöme är deras arvedel; och Gad och Ruben och ena hälften av Manasse stam hava redan fått sin arvedel på andra sidan Jordan, på östra sidan, den arvedel som HERRENS tjänare Mose gav dem.»
Och männen stodo upp och gingo åstad; och när de gingo åstad bjöd Josua dem att de skulle sätta upp en beskrivning över landet, i det han sade: »Gån åstad och dragen omkring i landet och sätten upp en beskrivning däröver, och vänden sedan tillbaka till mig, så vill jag kasta lott för eder här inför HERREN i Silo.»
Så gingo då männen åstad och drogo genom landet och satte upp en beskrivning över det, efter dess sju delar, med dess städer, och kommo så tillbaka till Josua i lägret vid Silo.
Sedan kastade Josua lott för dem i Silo inför HERREN, och Josua utskiftade där landet åt Israels barn, efter deras avdelningar.
Då nu lotten drogs för Benjamins barns stam, efter deras släkter, föll den ut så, att det område som lotten gav dem låg mellan Juda barns och Josefs barns områden.
Deras gräns på norra sidan begynte vid Jordan, och gränsen drog sig så upp mot Jerikos höjd i norr och uppåt bergsbygden västerut och gick så ut i öknen vid Bet-Aven.
Därifrån gick gränsen fram till Lus, till höjden söder om Lus, det är Betel; sedan gick gränsen ned till Atrot-Addar över berget söder om Nedre Bet-Horon.
Och gränsen drog sig vidare framåt och böjde sig på västra sidan söderut från berget som ligger gent emot Bet-Horon, söder därom, och gick så ut till Kirjat-Baal, det är staden Kirjat-Jearim inom Juda barns område.
Detta var västra sidan.
Och södra sidan begynte vid ändan av Kirjat-Jearims område, och gränsen gick så åt väster fram till Neftoavattnets källa.
Sedan gick gränsen ned till ändan av det berg som ligger gent emot Hinnoms sons dal, norrut i Refaimsdalen, och därefter ned i Hinnomsdalen, på södra sidan om Jebus' höjd, och gick så ned till Rogelskällan.
Därefter drog den sig norrut och gick fram till Semeskällan och vidare till Gelilot, som ligger mitt emot Adummimshöjden, och gick så ned till Bohans, Rubens sons, sten.
Vidare gick den fram till den höjd som ligger framför Hedmarken, norrut, och så ned till Hedmarken.
Sedan gick gränsen fram till Bet-Hoglas höjd, norrut, och så gick gränsen ut till Salthavets norra vik, vid Jordans södra ända.
Detta var södra gränsen.
Men på östra sidan var Jordan gränsen.
Detta var Benjamins barns arvedel med dess gränser runt omkring, efter deras släkter.
Och de städer som tillföllo Benjamins barns stam, efter deras släkter, voro: Jeriko, Bet-Hogla, Emek-Kesis,
Bet-Haaraba, Semaraim, Betel,
Avim, Para, Ofra,
Kefar-Haammoni, Ofni och Geba -- tolv städer med sina byar;
Gibeon, Rama, Beerot,
Mispe, Kefira, Mosa,
Rekem, Jirpeel, Tarala,
Sela, Elef, Jebus, det är Jerusalem, Gibeat och Kirjat -- fjorton städer med sina byar.
Detta var nu Benjamins barns arvedel, efter deras släkter.
Och den andra lotten föll ut för Simeon, för Simeons barns stam, efter deras släkter; och de fingo sin arvedel inom Juda barns arvedel.
De fingo inom dessas arvedel Beer-Seba, Seba, Molada,
Hasar-Sual, Bala, Esem,
Eltolad, Betul, Horma,
Siklag, Bet-Hammarkabot, Hasar-Susa,
Bet-Lebaot och Saruhen -- tretton städer med deras byar;
Ain, Rimmon, Eter och Asan -- fyra städer med deras byar;
därtill alla de byar som lågo runt omkring dessa städer, ända till Baalat-Beer, det sydliga Rama.
Detta var Simeons barns arvedel, efter deras släkter.
Ur Juda barns skifte fingo Simeons barn sin arvedel, ty Juda barns lott var för stor för dem; därför fingo Simeons barn sin arvedel inom deras arvedel.
Den tredje lotten drogs ut för Sebulons barn, efter deras släkter; och gränsen för deras arvedel gick ända till Sarid.
Därifrån drog sig deras gräns västerut uppåt till Mareala och träffade Dabbeset och träffade vidare dalen som ligger gent emot Jokneam.
På andra sidan från Sarid, österut mot solens uppgång, vände den sig åt Kislot-Tabors område och gick vidare till Dobrat och upp till Jafia.
Därifrån gick den fram österut mot solens uppgång till Gat-Hefer och Et-Kasin och vidare till det Rimmon som sträcker sig till Nea.
Härförbi böjde sig gränsen i norr till Hannaton och gick så ut vid Jifta-Els dal.
Och den omfattade Kattat, Nahalal, Simron, Jidala och Bet-Lehem -- tolv städer med deras byar.
Detta var Sebulons barns arvedel, efter deras släkter, de nämnda städerna med sina byar.
För Isaskar föll den fjärde lotten ut, för Isaskars barn, efter deras släkter.
Och deras gräns omfattade Jisreel, Kesullot, Sunem,
Hafaraim, Sion, Anaharat,
Rabbit, Kisjon, Ebes,
Remet, En-Gannim, En-Hadda och Bet-Passes;
och gränsen träffade Tabor, Sahasuma och Bet-Semes; och deras gräns gick ut vid Jordan -- sexton städer med deras byar.
Detta var Isaskars barns stams arvedel, efter deras släkter, städerna med sina byar.
Den femte lotten föll ut för Asers barns stam, efter deras släkter.
Och deras gräns omfattade Helkat, Hali, Beten, Aksaf,
Alammelek, Amead och Miseal; och vid havet träffade den Karmel och Sihor-Libnat.
Därefter vände den sig åt öster till Bet-Dagon och träffade Sebulon och Jifta-Els dal i norr, vidare Bet-Haemek och Negiel och gick så ut till Kabul i norr.
Och den omfattade Ebron, Rehob, Hammon och Kana, ända upp till Stora Sidon.
Och gränsen vände sig till Rama och gick fram till den befästa staden Tyrus; sedan vände sig gränsen till Hosa och gick så ut vid havet där landsträckan vid Aksib begynner.
Och den omfattade Umma, Afek och Rehob -- tjugutvå städer med deras byar.
Detta var Asers barns stams arvedel, efter deras släkter, de nämnda städerna med sina byar.
För Naftali barn föll den sjätte lotten ut, för Naftali barn, efter deras släkter.
Och deras gräns gick från Helef, från terebinten i Saanannim till Adami-Hannekeb och Jabneel, ända till Lackum, och gick så ut vid Jordan.
Och gränsen vände sig västerut till Asnot-Tabor och gick vidare därifrån till Huckok; den träffade Sebulon i söder, och Aser träffade den i väster och Juda med Jordan i öster.
Och den omfattade de befästa städerna Siddim, Ser och Hammat, Rackat och Kinneret,
Adama, Rama, Hasor,
Kedes, Edrei, En-Hasor,
Jireon och Migdal-El, Horem, Bet-Anat och Bet-Semes -- nitton städer med deras byar.
Detta var Naftali barns stams arvedel efter deras släkter, städerna med sina byar.
För Dans barns stam, efter deras släkter, föll den sjunde lotten ut.
Och gränsen för deras arvedel omfattade Sorga, Estaol, Ir-Semes,
Saalabbin, Ajalon, Jitla,
Elon, Timna, Ekron,
Elteke, Gibbeton, Baalat,
Jehud, Bene-Berak, Gat-Rimmon,
Me-Hajarkon och Harackon, tillika med området framför Jafo.
(Men när sedan Dans barns område gick förlorat för dem, drogo Dans barn upp och belägrade Lesem och intogo det och slogo dess invånare med svärdsegg; och sedan de så hade tagit det i besittning, bosatte de sig där och kallade Lesem för Dan, efter Dans, sin faders, namn.)
Detta var Dans barns stams arvedel, efter deras släkter, de nämnda städerna med sina byar.
När Israels barn så hade utskiftat landet efter dess gränser, gåvo de åt Josua, Nuns son, en särskild arvedel ibland sig.
Efter HERRENS befallning gåvo de honom nämligen den stad som han begärde, Timnat-Sera i Efraims bergsbygd; och han bebyggde staden och bosatte sig där.
Dessa voro de arvslotter som prästen Eleasar och Josua, Nuns son, och huvudmännen för familjerna inom Israels barns stammar utskiftade genom lottkastning i Silo inför HERRENS ansikte, vid ingången till uppenbarelsetältet.
Så avslutade de nu fördelningen av landet.
Och HERREN talade till Josua och sade:
»Tala till Israels barn och säg: Utsen åt eder de fristäder om vilka jag har talat till eder genom Mose,
de städer till vilka en dråpare som ouppsåtligen, utan vett och vilja, har dödat någon må kunna fly; och I skolen hava dem såsom tillflyktsorter undan blodshämnaren.
Och när någon flyr till en av dessa städer, skall han stanna vid ingången till stadsporten och omtala sin sak för de äldste i den staden; därefter må de taga honom in i staden till sig och giva honom en plats där han får bo ibland dem.
Och om blodshämnaren förföljer honom, skola de icke överlämna dråparen i hans hand, eftersom han utan vett och vilja har dödat sin nästa, och utan att förut hava burit hat till honom.
Och han skall stanna kvar där i staden, till dess han har stått till rätta inför menigheten, och till dess den dåvarande översteprästen har dött; sedan må dråparen vända tillbaka och komma till sin stad från vilken han har flytt.»
Så helgade de då därtill Kedes i Galileen, i Naftali bergsbygd, Sikem i Efraims bergsbygd och Kirjat-Arba, det är Hebron, i Juda bergsbygd.
Och på andra sidan Jordan mitt emot Jeriko, på östra sidan, utsågo de därtill inom Rubens stam Beser i öknen på slätten, inom Gads stam Ramot i Gilead, och inom Manasse stam Golan i Basan.
Dessa voro de städer som för alla Israels barn, och för de främlingar som bodde ibland dem, bestämdes att vara orter till vilka var och en som ouppsåtligen hade dödat någon finge fly, så att han skulle slippa dö för blodshämnarens hand, innan han hade stått till rätta inför menigheten.
Och huvudmännen för leviternas familjer trädde fram inför prästen Eleasar och Josua, Nuns son, och huvudmännen för familjerna inom Israels barns stammar
och talade till dem i Silo i Kanaans land, och sade: »HERREN bjöd genom Mose att man skulle giva oss städer att bo i, med tillhörande utmarker för vår boskap.»
Så gåvo då Israels barn, efter HERRES befallning, av sina arvslotter åt leviterna följande städer med tillhörande utmarker.
För kehatiternas släkter föll lotten ut så, att bland dessa leviter prästen Arons söner genom lotten fingo ur Juda stam, ur simeoniternas stam och ur Benjamins stam tretton städer.
Och Kehats övriga barn fingo genom lotten ur Efraims stams släkter, ur Dans stam och ur ena hälften av Manasse stam tio städer.
Gersons barn åter fingo genom lotten ur Isaskars stams släkter, ur Asers stam, ur Naftali stam och ur andra hälften av Manasse stam, i Basan, tretton städer.
Meraris barn fingo, efter sina släkter, ur Rubens stam, ur Gads stam och ur Sebulons stam tolv städer.
Israels barn gåvo nu åt leviterna dessa städer med tillhörande utmarker, genom lottkastning, såsom HERREN hade bjudit genom Mose.
Ur Juda barns stam och ur Simeons barns stam gav man följande här namngivna städer:
Bland kehatiternas släkter bland Levi barn fingo Arons söner följande, ty dem träffade lotten först:
Man gav dem Arbas, Anoks faders, stad, det är Hebron, i Juda bergsbygd, med dess utmarker runt omkring.
Men åkerjorden och byarna som hörde till staden gav man till besittning åt Kaleb, Jefunnes son.
Åt prästen Arons söner gav man alltså dråparfristaden Hebron med dess utmarker, vidare Libna med dess utmarker,
Jattir med dess utmarker, Estemoa med dess utmarker,
Holon med dess utmarker, Debir med dess utmarker,
Ain med dess utmarker, Jutta med dess utmarker och Bet-Semes med dess utmarker -- nio städer ur dessa två stammar;
och ur Benjamins stam Gibeon med dess utmarker, Geba med dess utmarker,
Anatot med dess utmarker och Almon med dess utmarker -- fyra städer.
De städer som Arons söner, prästerna, fingo utgjorde alltså tillsammans tretton städer, med tillhörande utmarker.
Och Kehats barns släkter av leviterna, nämligen de övriga Kehats barn, fingo ur Efraims stam följande städer, som lotten bestämde åt dem:
Man gav dem dråparfristaden Sikem med dess utmarker i Efraims bergsbygd, Geser med dess utmarker,
Kibsaim med dess utmarker och Bet-Horon med dess utmarker -- fyra städer;
och ur Dans stam Elteke med dess utmarker, Gibbeton med dess utmarker,
Ajalon med dess utmarker och Gat-Rimmon med dess utmarker -- fyra städer;
och ur ena hälften av Manasse stam Taanak med dess utmarker och Gat-Rimmon med dess utmarker -- två städer.
De städer som de övriga Kehats barns släkter fingo utgjorde alltså tillsammans tio, med tillhörande utmarker.
Bland leviternas släkter fingo vidare Gersons barn ur ena hälften av Manasse stam dråparfristaden Golan i Basan med dess utmarker och Beestera med dess utmarker -- två städer;
och ur Isaskars stam Kisjon med dess utmarker, Dobrat med dess utmarker,
Jarmut med dess utmarker och En-Gannim med dess utmarker -- fyra städer;
och ur Asers stam Miseal med dess utmarker, Abdon med dess utmarker,
Helkat med dess utmarker och Rehob med dess utmarker -- fyra städer;
och ur Naftali stam dråparfristaden Kedes i Galileen med dess utmarker, Hammot-Dor med dess utmarker och Kartan med dess utmarker -- tre städer.
Gersoniternas städer, efter deras släkter, utgjorde alltså tillsammans tretton städer, med tillhörande utmarker.
Och de övriga leviterna, Meraris barns släkter, fingo ur Sebulons stam Jokneam med dess utmarker, Karta med dess utmarker,
Dimna med dess utmarker och Nahalal med dess utmarker -- fyra städer.
64180
64190
och ur Gads stam dråparfristaden Ramot i Gilead med dess utmarker, Mahanaim med dess utmarker,
Hesbon med dess utmarker och Jaeser med dess utmarker -- tillsammans fyra städer.
De städer som dessa de övriga leviternas släkter, Meraris barn, fingo på sin lott, efter sina släkter, utgjorde alltså tillsammans tolv städer.
Tillsammans utgjorde levitstäderna inom Israels barns besittningsområde fyrtioåtta städer med tillhörande utmarker.
Var och en av dessa städer skulle bestå av själva staden och tillhörande utmarker runt omkring.
Så var det med alla dessa städer.
Så gav då HERREN åt Israel hela det land som han med ed hade lovat giva åt deras fäder; och de togo det i besittning och bosatte sig där.
Och HERREN lät dem hava ro på alla sidor, alldeles såsom han med ed hade lovat deras fäder; och ingen av deras fiender kunde stå dem emot, utan HERREN gav alla deras fiender i deras hand.
Intet uteblev av allt det goda som HERREN hade lovat Israels hus; det gick allt i fullbordan.
Då kallade Josua till sig rubeniterna och gaditerna och ena hälften av Manasse stam
och sade till dem: »I haven hållit allt vad HERRENS tjänare Mose har bjudit eder; I haven ock lyssnat till mina ord, vadhelst jag har befallt eder.
I haven under denna långa tid, ända till denna dag, icke övergivit edra bröder, och I haven hållit vad HERRENS, eder Guds, bud har befallt eder hålla.
Och nu har HERREN, eder Gud, låtit edra bröder komma till ro, såsom han lovade dem; så vänden nu om och gån hem till edra hyddor i det land I haven fått till besittning, det som HERRENS tjänare Mose har givit eder på andra sidan Jordan.
Allenast mån I noga hålla och göra efter de bud och den lag som HERRENS tjänare Mose har givit eder, så att I älsken HERREN, eder Gud, och alltid vandren på hans vägar och iakttagen hans bud och hållen eder till honom och tjänen honom av allt edert hjärta och av all eder själ.»
Och Josua välsignade dem och lät dem gå, och så gingo de hem till sina hyddor.
Ty åt ena hälften av Manasse stam hade Mose givit land i Basan, och åt andra hälften hade Josua givit land jämte deras bröder på andra sidan Jordan, på västra sidan.
Då nu Josua lät dem gå hem till sina hyddor, välsignade han dem
och sade till dem: »Vänden tillbaka till edra hyddor med de stora skatter I haven fått, med boskap i stor myckenhet, med silver, guld, koppar och järn och kläder i stor myckenhet; skiften så med edra bröder bytet från edra fiender.»
Så vände då Rubens barn och Gads barn och ena hälften av Manasse stam tillbaka, och gingo bort ifrån de övriga israeliterna, bort ifrån Silo i Kanaans land, för att begiva sig till Gileads land, det land de hade fått till besittning, och där de skulle hava sina besittningar, efter HERRENS befallning genom Mose.
När så Rubens barn och Gads barn och ena hälften av Manasse stam kommo till stenkretsarna vid Jordan i Kanaans land, byggde de där ett altare vid Jordan, ett ansenligt altare.
Och de övriga israeliterna fingo höra sägas: »Se, Rubens barn och Gads barn och ena hälften av Manasse stam hava byggt ett altare mitt emot Kanaans land, i stenkretsarna vid Jordan, på andra sidan om de övriga israeliternas område.»
När Israels barn hörde detta, församlade sig deras hela menighet i Silo för att draga upp till strid mot dem.
Därefter sände Israels barn Pinehas till Rubens barn och Gads barn och ena hälften av Manasse stam, i Gileads land, Pinehas, prästen Eleasars son,
och med honom tio hövdingar, en hövding för var stamfamilj inom Israels alla stammar; var och en av dem var huvudman för sin familj inom Israels ätter.
Och när dessa kommo till Rubens barn och Gads barn och ena hälften av Manasse stam, i Gileads land, talade de till dem och sade:
»Så säger hela HERRENS menighet: Vad är detta för en otrohet som I haven begått mot Israels Gud, då I haven vänt eder bort ifrån HERREN, därigenom att I haven byggt eder ett altare och sålunda nu satt eder upp mot HERREN?
Är det icke nog att vi hava begått missgärningen med Peor, från vilken vi ännu i dag icke hava blivit renade, och för vilken en hemsökelse drabbade HERRENS menighet?
Viljen I nu ytterligare vända eder bort ifrån HERREN?
Om I i dag sätten eder upp mot HERREN, så skall förvisso i morgon hans förtörnelse drabba Israels hela menighet.
Men om det land I haven fått till besittning tyckes eder vara orent, så dragen över till det land HERREN har tagit till besittning, där HERRENS tabernakel har sin plats, och haven edra besittningar där bland oss.
Sätten eder icke upp mot HERREN och sätten eder icke upp mot oss genom att bygga eder ett altare, ett annat än HERRENS, vår Guds, altare.
När Akan, Seras son, hade trolöst förgripit sig på det tillspillogivna, kom icke då förtörnelse över Israels hela menighet, så att han själv icke blev den ende som förgicks genom den missgärningen?
Då svarade Rubens barn och Gads barn och ena hälften av Manasse stam och talade till huvudmännen för Israels ätter:
»Gud, HERREN Gud, ja, Gud, HERREN Gud, han vet det, och Israel må ock veta det: Sannerligen, om detta har skett i upproriskhet och otrohet mot HERREN -- du må då i dag undandraga oss din hjälp! --
om vi hava byggt altaret åt oss, därför att vi vilja vända oss bort ifrån HERREN, och om vi vilja offra därpå brännoffer eller spisoffer eller frambära tackoffer därpå, då må HERREN själv utkräva vad vi hava förskyllt.
Nej, vi hava sannerligen gjort så av fruktan för vad som kunde hända, i det att vi tänkte att edra barn i framtiden skulle kunna säga till våra barn: 'Vad haven I att göra med HERREN, Israels Gud?
HERREN har ju satt Jordan till gräns mellan oss och eder, I Rubens barn och Gads barn; alltså haven I ingen del i HERREN.'
Och så skulle edra barn kunna hindra våra barn från att frukta HERREN.
Därför sade vi: Må vi gripa oss an och bygga detta altare, men icke till brännoffer eller till slaktoffer,
utan till att vara ett vittne mellan oss och eder, och mellan bådas efterkommande efter oss, att vi vilja förrätta HERRENS tjänst inför hans ansikte med våra brännoffer och slaktoffer och tackoffer, så att edra barn i framtiden icke kunna säga till våra barn: 'I haven ingen del i HERREN.'
Och vi tänkte: Om det i framtiden händer att de så säga till oss och våra efterkommande, då kunna vi svara: 'Sen på den bild av HERRENS altare, som våra fäder hava gjort, men icke till brännoffer eller till slaktoffer, utan till att vara ett vittne mellan oss och eder.'
Bort det, att vi skulle sätta oss upp mot HERREN och nu vända oss bort ifrån HERREN genom att bygga ett altare till brännoffer eller till spisoffer eller slaktoffer, ett annat än HERRENS, vår Guds, altare, som står framför hans tabernakel.»
Då nu prästen Pinehas och menighetens hövdingar, nämligen huvudmännen för Israels ätter, som voro med honom, hörde vad Rubens barn, Gads barn och Manasse barn talade, behagade det dem.
Och Pinehas, prästen Eleasars son, sade till Rubens barn, Gads barn och Manasse barn: »Nu hava vi förnummit att HERREN är mitt ibland oss, därav nämligen, att I icke haven velat begå en sådan otrohet mot HERREN.
Därmed haven I ock räddat Israels barn undan HERRENS hand.»
Därefter vände Pinehas, prästen Eleasars son, jämte hövdingarna tillbaka från Rubens barn och Gads barn, i Gileads land, in i Kanaans land till de övriga israeliterna och avgåvo sin berättelse härom inför dem.
Denna behagade Israels barn, och Israels barn lovade Gud; och de tänkte icke mer på att draga upp till strid mot dem, för att fördärva det land där Rubens barn och Gads barn bodde.
Och Rubens barn och Gads barn gåvo namn åt altaret; de sade: »Ett vittne är det mellan oss, att HERREN är Gud.»
En lång tid härefter, när HERREN hade låtit Israel få ro för alla dess fiender runt omkring, och då Josua var gammal och kommen till hög ålder,
kallade han till sig hela Israel, dess äldste, dess huvudmän, dess domare och tillsyningsmän och sade till dem: »Jag är nu gammal och kommen till hög ålder.
Och I haven själva sett allt vad HERREN, eder Gud, gjorde med alla dessa folk, när I drogen härin, ty HERREN eder Gud, stridde själv för eder.
Se, dessa folk som ännu äro kvar har jag genom lottkastning fördelat åt eder till arvedel, efter edra stammar, allt ifrån Jordan intill Stora havet västerut, för att icke nämna alla de folk jag har utrotat.
Och HERREN, eder Gud, skall själv driva dem undan för eder och förjaga dem för eder, så att I skolen taga deras land i besittning, såsom HERREN, eder Gud, har lovat eder.
Men varen I nu ståndaktiga i att hålla och göra allt vad som är föreskrivet i Moses lagbok, så att I icke viken av därifrån vare sig till höger eller till vänster,
och icke träden i gemenskap med dessa folk som ännu äro kvar här jämte eder, ej heller nämnen deras gudars namn eller svärjen vid dem eller tjänen och tillbedjen dem.
Nej, till HERREN, eder Gud, skolen I hålla eder, såsom I haven gjort ända till denna dag,
varför ock HERREN har fördrivit för eder stora och mäktiga folk, så att ingen har kunnat stå eder emot ända till denna dag.
En enda man bland eder jagade tusen framför sig, ty HERREN, eder Gud, stridde själv för eder, såsom han hade lovat eder.
Så haven nu noga akt på eder själva, så att I älsken HERREN, eder Gud.
Ty om I vänden eder bort ifrån honom, och hållen eder till återstoden av dessa folk som ännu äro kvar här jämte eder, och befrynden eder med dem, så att I träden i gemenskap med dem och de med eder,
då mån I förvisso veta att HERREN, eder Gud, icke mer skall fördriva dessa folk undan för eder, utan de skola bliva eder till en snara och ett giller och bliva ett gissel för edra sidor och taggar i edra ögon, till dess I bliven utrotade ur detta goda land, som HERREN, eder Gud, har givit eder.
Se, jag går nu all världens väg.
Så besinnen då av allt edert hjärta och av all eder själ att intet har uteblivit av allt det goda som HERREN, eder Gud, har lovat angående eder; det har allt gått i fullbordan för eder, intet därav har uteblivit.
Men likasom allt det goda som HERREN, eder Gud, lovade eder har kommit över eder, så skall ock HERREN låta allt det onda komma över eder, till dess han har förgjort eder ur detta goda land, som HERREN, eder Gud, har givit eder.
Om I nämligen överträden HERRENS, eder Guds, förbund, det som han har stadgat för eder, och gån åstad och tjänen andra gudar och tillbedjen dem, så skall HERRENS vrede upptändas mot eder, och I skolen med hast bliva utrotade ur det goda land som han har givit eder.»
Och Josua församlade alla Israels stammar till Sikem; och han kallade till sig de äldste i Israel, dess huvudmän, dess domare och dess tillsyningsmän, och de trädde fram inför Gud.
Och Josua sade till allt folket: »Så säger HERREN, Israels Gud: På andra sidan floden bodde edra fäder i forna tider; så gjorde ock Tera, Abrahams och Nahors fader.
Och de tjänade där andra gudar.
Men jag hämtade eder fader Abraham från andra sidan floden och lät honom vandra omkring i hela Kanaans land.
Och jag gjorde hans säd talrik; jag gav honom Isak,
och åt Isak gav jag Jakob och Esau.
Och jag gav Seirs bergsbygd till besittning åt Esau; men Jakob och hans söner drogo ned till Egypten.
Sedan sände jag Mose och Aron och hemsökte Egypten med de gärningar jag där gjorde, och därefter förde jag eder ut.
Och när jag förde edra fäder ut ur Egypten och I haden kommit till havet, förföljde egyptierna edra fäder med vagnar och ryttare ned i Röda havet.
Då ropade de till HERREN, och han satte ett tjockt mörker mellan eder och egyptierna och lät havet komma över dem, så att det övertäckte dem; ja, I sågen med egna ögon vad jag gjorde med egyptierna.
Sedan bodden I i öknen en lång tid.
Därefter förde jag eder in i amoréernas land, vilka bodde på andra sidan Jordan, och de inläto sig i strid med eder; men jag gav dem i eder hand, så att I intogen deras land, och jag förgjorde dem för eder.
Då uppreste sig Balak, Sippors son, konungen i Moab, och gav sig i strid med Israel.
Och han sände och lät kalla till sig Bileam, Beors son, för att denne skulle förbanna eder.
Men jag ville icke höra på Bileam, utan han måste välsigna eder, och jag räddade eder ur hans hand.
Och när I haden gått över Jordan och kommit till Jeriko, gåvo sig Jerikos borgare i strid med eder, så och amoréerna, perisséerna, kananéerna, hetiterna och girgaséerna, hivéerna och jebuséerna; men jag gav dem i eder hand.
Och jag sände getingar framför eder, och genom dessa förjagades amoréernas två konungar för eder, icke genom ditt svärd eller din båge.
Och jag gav eder ett land varpå du icke hade nedlagt något arbete, så ock städer som I icke haden byggt, och i dem fingen I bo; och av vingårdar och olivplanteringar som I icke haden planterat fingen I äta.
Så frukten nu HERREN och tjänen honom ostraffligt och troget; skaffen bort de gudar som edra fäder tjänade på andra sidan floden och i Egypten, och tjänen HERREN.
Men om det misshagar eder att tjäna HERREN, så utväljen åt eder i dag vem I viljen tjäna, antingen de gudar som edra fäder tjänade, när de bodde på andra sidan floden, eller de gudar som dyrkas av amoréerna, i vilkas land I själva bon.
Men jag och mitt hus, vi vilja tjäna HERREN.»
Då svarade folket och sade: »Bort det, att vi skulle övergiva HERREN och tjäna andra gudar!
Nej, HERREN är vår Gud, han är den som har fört oss och våra fäder upp ur Egyptens land, ur träldomshuset, och som inför våra ögon har gjort dessa stora under, och bevarat oss på hela den väg vi hava vandrat och bland alla de folk genom vilkas land vi hava dragit fram.
HERREN har förjagat för oss alla dessa folk, så ock amoréerna som bodde i landet.
Därför vilja vi ock tjäna HERREN; ty an är vår Gud.»
Josua sade till folket: »I kunnen icke tjäna HERREN, ty han är en helig Gud; han är en nitälskande Gud, han skall icke hava fördrag med edra överträdelser och synder.
Om I övergiven HERREN och tjänen främmande gudar, så skall han vända sig bort och låta det gå eder illa och förgöra eder, i stället för att han hittills har låtit det gå eder väl.»
Men folket sade till Josua: »Icke så, utan vi vilja tjäna HERREN.»
Då sade Josua till folket: »I ären nu själva vittnen mot eder, att I haven utvalt HERREN åt eder, för att tjäna honom.»
De svarade: »Ja.»
Han sade: »Så skaffen nu bort de främmande gudar som I haven bland eder, och böjen edra hjärtan till HERREN, Israels Gud.»
Folket svarade Josua: »HERREN, vår Gud, vilja vi tjäna, och hans röst vilja vi höra.»
Så slöt då Josua på den dagen ett förbund med folket och förelade dem lag och rätt i Sikem.
Och Josua tecknade upp allt detta i Guds lagbok.
Och han tog en stor sten och reste den där, under eken som stod vid HERRENS helgedom.
Och Josua sade till allt folket: »Se, denna sten skall vara vittne mot oss, ty den har hört alla de ord som HERREN har talat med oss; den skall vara vittne mot eder, så att I icke förneken eder Gud.»
Sedan lät Josua folket gå, var och en till sin arvedel.
En tid härefter dog HERRENS tjänare Josua, Nuns son, ett hundra tio år gammal.
Och man begrov honom på hans arvedels område, i Timnat-Sera i Efraims bergsbygd, norr om berget Gaas.
Och Israel tjänade HERREN, så länge Josua levde, och så länge de äldste levde, de som voro kvar efter Josua, och som visste av alla de gärningar HERREN hade gjort för Israel.
Och Josefs ben, som Israels barn hade fört upp ur Egypten, begrovo de i Sikem, på det jordstycke som Jakob hade köpt av Hamors, Sikems faders, barn för hundra kesitor; Josefs barn fingo detta till arvedel.
Och Eleasar, Arons son, dog, och man begrov honom i hans son Pinehas' stad, Gibea, som hade blivit denne given i Efraims bergsbygd.
Efter Josuas död frågade Israels barn HERREN och sade: »Vem bland oss skall först draga upp mot kananéerna och strida mot dem?»
HERREN sade: »Juda skall göra det; se, jag har givit landet i hans hand.»
Då sade Juda till sin broder Simeon: »Drag upp med mig in i min arvslott, och låt oss strida mot kananéerna, så skall jag sedan tåga med dig in i din arvslott.»
Så tågade då Simeon med honom.
När nu Juda drog ditupp, gav HERREN kananéerna och perisséerna i deras hand, så att de slogo dem vid Besek, tio tusen man.
Ty vid Besek träffade de på Adoni-Besek och stridde mot honom och slogo så kananéerna och perisséerna.
Och Adoni-Besek flydde, men de förföljde honom och grepo honom och höggo av honom hans tummar och stortår.
Då sade Adoni-Besek: »Sjuttio konungar med avhuggna tummar och stortår hämtade upp smulorna under mitt bord; efter mina gärningar har Gud nu vedergällt mig.»
Sedan förde de honom till Jerusalem, och där dog han.
Men Juda barn belägrade Jerusalem och intogo det och slogo dess invånare med svärdsegg; därefter satte de eld på staden.
Sedan drogo Juda barn ned för att strida mot de kananéer som bodde i Bergsbygden, i Sydlandet och i Låglandet.
Och Juda tågade åstad mot de kananéer som bodde i Hebron -- vilket fordom hette Kirjat-Arba -- och de slogo Sesai, Ahiman och Talmai.
Därifrån tågade de åstad mot Debirs invånare.
Men Debir hette fordom Kirjat-Sefer.
Och Kaleb sade: »Åt den som angriper Kirjat-Sefer och intager det vill jag giva min dotter Aksa till hustru.»
När då Otniel, son till Kenas, Kalebs yngre broder, intog det, gav han honom sin dotter Aksa till hustru.
Och när hon kom till honom, intalade hon honom att begära ett stycke åkermark av hennes fader; och hon steg hastigt ned från åsnan.
Då sade Kaleb till henne: »Vad önskar du?»
Hon sade till honom: »Låt mig få en avskedsskänk; eftersom du har gift bort mig till det torra Sydlandet, må du giva mig vattenkällor.»
Då gav Kaleb henne Illitkällorna och Tatitkällorna.
Och kainéens, Moses svärfaders, barn hade dragit upp från Palmstaden med Juda barn till Juda öken, söder om Arad; de gingo åstad och bosatte sig bland folket där.
Men Juda tågade åstad med sin broder Simeon, och de slogo de kananéer som bodde i Sefat; och de gåvo staden till spillo; så fick den namnet Horma.
Därefter intog Juda Gasa med dess område, Askelon med dess område och Ekron med dess område.
Och HERREN var med Juda, så att de intogo bergsbygden; men de kunde icke fördriva dem som bodde i dalbygden, därför att dessa hade stridsvagnar av järn.
Och de gåvo Hebron åt Kaleb, såsom Mose hade föreskrivit; och han fördrev därifrån Anaks tre söner.
Men jebuséerna, som bodde i Jerusalem, blevo icke fördrivna av Benjamins barn; därför bodde ock jebuséerna kvar bland Benjamins barn i Jerusalem, såsom de göra ännu dag.
Så drogo ock männen av Josefs hus upp till Betel, och HERREN var med dem.
Och männen av Josefs hus läto bespeja Betel, samma stad som fordom hette Lus.
Då fingo deras kunskapare se en man gå ut ur staden, och de sade till honom: »Visa oss var vi kunna komma in i staden, så vilja vi sedan göra barmhärtighet med dig.»
När han sedan hade visat dem var de kunde komma in i staden, slog de stadens invånare med svärdsegg; men den mannen och hela hans släkt läto de gå.
Och mannen begav sig till hetiternas land; där byggde han en stad och gav den namnet Lus, såsom den heter ännu i dag.
Men Manasse intog icke Bet-Sean med underlydande orter, ej heller Taanak med underlydande orter; och ej heller fördrevo de invånarna i Dor och underlydande orter, ej heller invånarna i Jibleam och underlydande orter, ej heller invånarna i Megiddo och underlydande orter, utan kananéerna förmådde hålla sig kvar där i landet.
När sedan israeliterna blevo de starkare, läto de kananéerna bliva arbetspliktiga under sig; de fördrevo dem icke heller då.
Icke heller fördrev Efraim de kananéer som bodde i Geser, utan kananéerna bodde kvar bland dem där i Geser.
Sebulon fördrev icke invånarna i Kitron och invånarna i Nahalol, utan kananéerna bodde kvar bland dem, men blevo arbetspliktiga under dem.
Aser fördrev icke invånarna i Acko eller invånarna i Sidon, ej heller dem i Alab, Aksib, Helba, Afik och Rehob.
Alltså bodde aseriterna bland kananéerna, landets gamla inbyggare; ty de fördrevo dem icke.
Naftali fördrev icke invånarna i Bet-Semes, ej heller invånarna i Bet-Anat, utan bodde ibland kananéerna, landets gamla inbyggare; men invånarna i Bet-Semes och Bet-Anat blevo arbetspliktiga åt dem.
Men amoréerna trängde undan Dans barn till bergsbygden, ty de tillstadde dem icke att komma ned till dalbygden.
Och amoréerna förmådde hålla sig kvar i Har-Heres, Ajalon och Saalbim; men Josefs barns hand blev tung över dem, så att de blevo arbetspliktiga under dessa.
Och amoréernas område sträckte sig från Skorpionhöjden, från Sela vidare uppåt.
Och HERRENS ängel kom från Gilgal upp till Bokim.
Och han sade: »Jag förde eder upp ur Egypten och lät eder komma in i det land som jag med ed hade lovat åt edra fäder; och jag sade: 'Jag skall icke bryta mitt förbund med eder till evig tid.
I åter skolen icke sluta förbund med detta lands inbyggare; I skolen bryta ned deras altaren.'
Men I haven icke velat höra min röst.
Vad haven I gjort! --
Därför säger jag nu ock: 'Jag vill icke förjaga dem för eder, utan de skola tränga eder i sidorna, och deras gudar skola bliva eder till en snara.'»
När HERRENS ängel hade talat dessa ord till alla Israels barn, brast folket ut i gråt.
Och de gåvo den platsen namnet Bokim; och de offrade där åt HERREN.
Sedan Josua hade låtit folket gå, drogo Israels barn åstad var och en till sin arvedel, för att taga landet i besittning.
Och folket tjänade HERREN, så länge Josua levde, och så länge de äldste levde, de som voro kvar efter Josua, dessa som hade sett alla de stora gärningar HERREN hade gjort för Israel.
Men HERRENS tjänare Josua, Nuns son, dog, när han var ett hundra tio år gammal.
Och man begrov honom på hans arvedels område i Timna-Heres i Efraims bergsbygd, norr om berget Gaas.
När sedan också hela det släktet hade blivit samlat till sina fäder, kom ett annat släkte upp efter dem, ett som icke visste av HERREN eller de gärningar som han hade gjort för Israel.
Då gjorde Israels barn vad ont var i HERRENS ögon och tjänade Baalerna.
De övergåvo HERREN, sina fäders Gud, som hade fört dem ut ur Egyptens land, och följde efter andra gudar, de folks gudar, som bodde omkring dem, och dessa tillbådo de; därmed förtörnade de HERREN.
Ty när de övergåvo HERREN och tjänade Baal och Astarterna,
upptändes HERRENS vrede mot i Israel, och han gav dem i plundrares hand, och dessa utplundrade dem; han sålde dem i deras fienders hand där runt omkring, så att de icke mer kunde stå emot sina fiender.
Varthelst de drogo ut var HERRENS hand emot dem, så att de kommo i olycka, såsom HERREN hade hotat, och såsom HERREN hade svurit att det skulle gå dem, och de kommo i stor nöd.
Då lät HERREN domare uppstå, som frälste dem ur deras plundrares hand.
Men de hörde icke heller på sina domare, utan lupo i trolös avfällighet efter andra gudar och tillbådo dem; de veko med hast av ifrån den väg som deras fäder hade vandrat, i lydnad för HERRENS bud, och gjorde icke såsom de.
När HERREN alltså lät någon domare uppstå bland dem, var han med domaren och frälste dem ur deras fienders hand, så länge domaren levde; ty då de jämrade sig över sina förtryckare och plågare, förbarmade sig HERREN.
Men när domaren dog, vände de tillbaka och togo sig till vad fördärvligt var, ännu mer än deras fäder, så att de följde efter andra gudar och tjänade och tillbådo dem; de avstodo icke från sina gärningar och sin hårdnackenhet.
Därför upptändes HERRENS vrede mot Israel, så att han sade: »Eftersom detta folk har överträtt det förbund som jag stadgade för deras fäder, och icke har velat höra min röst,
därför skall icke heller jag hädanefter fördriva för dem en enda man av de folk som Josua lämnade efter sig, när han dog;
ty jag skall med dem sätta Israel på prov, om de vilja hålla HERRENS väg och vandra därpå, såsom deras fäder hava hållit den, eller om de icke vilja det.»
Alltså lät HERREN dessa folk bliva kvar och fördrev dem icke med hast; han gav dem icke i Josuas hand.
Dessa voro de folk som HERREN lät bliva kvar, för att genom dem sätta Israel på prov, alla de israeliter nämligen, som icke hade varit med om alla krigen i Kanaan
-- allenast på det att dessa Israels barns efterkommande skulle få vara med om sådana, för att han så skulle lära dem att föra krig, dock allenast dem som förut icke hade varit med om sådana --:
filistéernas fem hövdingar och alla kananéer och sidonier, samt de hivéer som bodde i Libanons bergsbygd, från berget Baal-Hermon ända dit där vägen går till Hamat.
Med dessa ville HERREN sätta Israel på prov, för att förnimma om de ville hörsamma de bud som han hade givit deras fäder.
Då nu Israels barn bodde: ibland kananéerna, hetiterna, amoréerna, perisséerna, hivéerna och jebuséerna,
togo de deras döttrar till hustrur åt sig och gåvo sina döttrar åt deras söner och tjänade deras gudar.
Så gjorde Israels barn vad ont var i HERRENS ögon och glömde HERREN, sin Gud, och tjänade Baalerna och Aserorna.
Då upptändes HERRENS vrede mot Israel, och han sålde dem i Kusan-Risataims hand, konungens i Aram-Naharaim; och Israels barn måste tjäna Kusan-Risataim i åtta år.
Men Israels barn ropade till HERREN, och HERREN lät då bland Israels barn en frälsare uppstå, som frälste dem, nämligen Otniel, son till Kenas, Kalebs yngre broder.
HERRENS Ande kom över honom, och han blev domare i Israel, och när han drog ut till strid, gav HERREN Kusan-Risataim, konungen i Aram, i hans hand, så att hans hand blev Kusan-Risataim övermäktig.
Och landet hade nu ro i fyrtio år; så dog Otniel, Kenas' son.
Men Israels barn gjorde åter vad ont var i HERRENS ögon, då gav HERREN Eglon, konungen i Moab, makt över Israel, eftersom de gjorde vad ont var i HERRENS ögon.
Denne förenade med sig Ammons barn och Amalek; sedan tågade han åstad och slog Israel, varefter de intogo Palmstaden.
Och Israels barn måste nu tjäna: Eglon, konungen i Moab, i aderton år.
Men Israels barn ropade till HERREN, och HERREN lät då bland dem en frälsare uppstå, benjaminiten Ehud, Geras son, en vänsterhänt man.
När Israels barn genom honom skulle sända sina skänker till Eglon, konungen i Moab,
gjorde sig Ehud ett tveeggat svärd, en fot långt; och han band detta under sina kläder vid sin högra länd.
Så överlämnade han skänkerna till Eglon, konungen i Moab.
Men Eglon var en mycket fet man.
När han nu hade överlämnat skänkerna, lät han folket som hade burit dem gå sin väg.
Men själv vände han tillbaka från Belätesplatsen vid Gilgal och lät säga: »Jag har ett hemligt ärende till dig, o konung.»
När denne då sade: »Lämnen oss i ro», gingo alla de som stodo omkring honom ut därifrån.
Men sedan Ehud hade kommit in till honom, där han satt i sommarsalen, som han hade för sig allena, sade Ehud: »Jag har ett ord från Gud att säga dig.»
Då stod han upp från sin stol.
Men Ehud räckte ut sin vänstra hand och tog svärdet från sin högra länd och stötte det i hans buk,
så att ock fästet följde med in efter klingan, och klingan omslöts av fettet, ty han drog icke ut svärdet ur hans buk.
Därefter gick Ehud ut i försalen;
och när han hade kommit ditut, i förhallen, stängde han igen dörrarna till salen efter sig och riglade dem.
Sedan, då han hade gått sin väg, kommo Eglons tjänare, och när de fingo se att dörrarna till salen voro riglade, tänkte de: »Förvisso har han något avsides bestyr i sin sommarkammare.»
Men sedan de hade väntat länge och väl, och han ändå icke öppnade dörrarna till salen, togo de nyckeln och öppnade själva, och se, då låg deras herre död där på golvet.
Men Ehud hade flytt undan, medan de dröjde; han hade redan hunnit förbi Belätesplatsen och flydde sedan undan till Seira.
Och så snart han hade kommit hem, lät han stöta i basun Efraims bergsbygd; då drogo Israels barn ned från bergsbygden med honom i spetsen för sig.
Och han sade till dem: »Följen efter mig, ty HERREN har givit edra fiender, moabiterna, i eder hand.»
Då drogo de efter honom längre ned och besatte vadställena över Jordan för moabiterna och läto ingen komma över.
Där slogo de då moabiterna, vid pass tio tusen man, allasammans ansenligt och tappert folk; icke en enda kom undan.
Så blev Moab då kuvat under Israels hand.
Och landet hade nu ro i åttio år.
Efter honom kom Samgar, Anats son; han slog filistéerna, sex hundra man, med en oxpik.
Också han frälste Israel.
Men Israels barn gjorde åter vad ont var i HERRENS ögon, när Ehud var död.
Då sålde HERREN dem i Jabins hand, den kananeiske konungens, som regerade i Hasor.
Hans härhövitsman var Sisera, och denne bodde i Haroset-Haggoim.
Och Israels barn ropade till HERREN; ty han hade nio hundra stridsvagnar av järn, och han förtryckte Israels barn våldsamt i tjugu år.
Men Debora, en profetissa, Lappidots hustru, var på den tiden domarinna i Israel.
Hon plägade sitta under Deborapalmen, mellan Rama och Betel i Efraims bergsbygd, och Israels barn drogo ditupp till henne, for att hon skulle skipa rätt.
Hon sände nu och lät kalla till sig Barak, Abinoams son, från Kedes i Naftali, och sade till honom: »Se, HERREN, Israels Gud, bjuder: Drag åstad upp på berget Tabor och tag med dig tio tusen man av Naftali barn och Sebulons barn.
Ty jag vill draga Sisera, Jabins härhövitsman, med hans vagnar och skaror, till dig vid bäcken Kison och giva honom i din hand.»
Barak sade till henne: »Om du går med mig, så går jag, men om du icke går med mig, så går icke heller jag.»
Då svarade hon: »Ja, jag skall gå med dig; dock skall äran då icke bliva din på den väg du nu går, utan HERREN skall sälja Sisera i en kvinnas hand.»
Så stod Debora upp och gick med Barak till Kedes.
Då bådade Barak upp Sebulon och Naftali till Kedes, och tio tusen man följde honom ditupp; Debora gick ock ditupp med honom.
Men kainéen Heber hade skilt sig från de övriga kainéerna, Hobabs, Moses svärfaders, barn; och han hade sina tältplatser ända till terebinten i Saannim vid Kedes.
Och man berättade för Sisera att Barak, Abinoams son, hade dragit upp på berget Tabor.
Då bådade Sisera upp alla sina stridsvagnar, nio hundra vagnar av järn, därtill ock allt folk han hade, att draga från Haroset-Haggoim till bäcken Kison.
Men Debora sade till Barak: »Stå upp, ty detta är den dag på vilken HERREN har givit Sisera i din hand; se, HERREN har dragit ut framför dig.»
Så drog då Barak ned från berget Tabor, och tio tusen man följde honom.
Och HERREN sände förvirring över Sisera och alla hans vagnar och hela hans här, så att de veko tillbaka för Baraks svärd; och Sisera steg ned från sin vagn och flydde till fots.
Och Barak jagade efter vagnarna och hären ända till Haroset-Haggoim.
Och hela Siseras här föll för svärdsegg; icke en enda kom undan.
Men Sisera hade under flykten styrt sina steg till Jaels, kainéen Hebers hustrus, tält; ty vänskap rådde mellan Jabin, konungen i Hasor, och kainéen Hebers hus.
Då gick Jael ut emot Sisera och sade till honom: »Kom in, min herre, kom in till mig, frukta intet.»
Så gick han då in till henne i tältet, och hon höljde över honom med ett täcke.
Och han sade till henne: »Giv mig litet vatten att dricka, ty jag är törstig.»
Då öppnade hon mjölk- kärlet och gav honom att dricka och höljde sedan åter över honom.
Och han sade till henne: »Ställ dig vid ingången till tältet; och kommer någon och frågar dig om någon är här, så svara nej.»
Men Jael, Hebers hustru, grep en tältplugg och tog en hammare i sin hand, gick därefter sakta in till honom och slog pluggen genom tinningen på honom, så att den gick ned i marken.
Så dödades han, där han låg försänkt i tung sömn, medtagen av trötthet.
I samma stund kom Barak jagande efter Sisera; då gick Jael ut emot honom och sade till honom: »Kom hit, så skall jag visa dig den man som du söker.»
När han då gick in till henne, fick han se Sisera ligga död där, med tältpluggen genom tinningen.
Så lät Gud på den dagen Jabin, konungen i Kanaan, bliva kuvad av Israels barn.
Och Israels barns hand vilade allt tyngre på Jabin, konungen i Kanaan; och till slut förgjorde de Jabin, konungen i Kanaan.
De sjöngo Debora och Barak, Abinoams son, denna sång:
Att härförare förde an i Israel, att folket villigt följde dem -- loven HERREN därför!
Hören, I konungar; lyssnen, I furstar.
Till HERRENS ära vill jag, vill jag sjunga, lovsäga HERREN, Israels Gud.
HERRE, när du drog ut från Seir, när du gick fram ifrån Edoms mark, då bävade jorden, då strömmade det från himmelen, då strömmade vatten ned ifrån molnen;
bergen skälvde inför HERRENS ansikte, ja, Sinai inför HERRENS, Israels Guds, ansikte.
I Samgars dagar, Anats sons, i Jaels dagar lågo vägarna öde; vandrarna måste färdas svåra omvägar.
Inga styresmän funnos, inga funnos mer i Israel, förrän du stod upp, Debora, stod upp såsom en moder i Israel.
Man valde sig nya gudar; då nådde striden fram till portarna.
Men ingen sköld, intet spjut var att se hos de fyrtio tusen i Israel.
Mitt hjärta tillhör Israels hövdingar och dem bland folket, som villigt följde;
ja, loven HERREN.
I som riden på vita åsninnor, I som sitten hemma på mattor, och I som vandren på vägen, talen härom.
När man under rop skiftar byte mellan vattenhoarna, då lovprisar man där HERRENS rättfärdiga gärningar, att han i rättfärdighet regerar i Israel.
Då drog HERRENS folk ned till portarna.
Upp, upp, Debora!
Upp, upp, sjung din sång!
Stå upp, Barak; tag dig fångar, du Abinoams son.
Då satte folkets kvarleva de tappre till anförare, HERREN satte mig till anförare över hjältarna.
Från Efraim kommo män som hade rotfäst sig i Amalek; Benjamin följde dig och blandade sig med dina skaror.
Ned ifrån Makir drogo hövdingar åstad, och från Sebulon män som buro anförarstav.
Furstarna i Isaskar slöto sig till Debora; och likasom Isaskar, så gjorde ock Barak; ned i dalen skyndade man i dennes spår.
Bland Rubens ätter höllos stora rådslag.
Men varför satt du kvar ibland dina fållor och lyssnade till flöjtspel vid hjordarna?
Ja, av Rubens ätter fördes stora överläggningar.
Gilead stannade på andra sidan Jordan.
Och Dan varför -- dröjer han ännu vid skeppen?
Aser satt kvar vid havets strand, vid sina vikar stannade han.
Men Sebulon var ett folk som prisgav sitt liv åt döden, Naftali likaså, på stridsfältets höjder.
Konungar drogo fram och stridde ja, då stridde Kanaans konungar vid Taanak, invid Megiddos vatten; men byte av silver vunno de icke.
Från himmelen fördes strid, stjärnorna stridde från sina banor mot Sisera.
Bäcken Kison ryckte dem bort, urtidsbäcken, bäcken Kison.
Gå fram, min själ, med makt!
Då stampade hästarnas hovar, när deras tappra ryttare jagade framåt, framåt.
Förbannen Meros, säger HERRENS ängel, ja, förbannen dess inbyggare, därför att de ej kommo HERREN till hjälp, HERREN till hjälp bland hjältarna.
Välsignad vare Jael framför andra kvinnor, Hebers hustru, kainéens, välsignad framför alla kvinnor som bo i tält!
Vatten begärde han; då gav hon honom mjölk, gräddmjölk bar hon fram i högtidsskålen.
Sin hand räckte hon ut efter tältpluggen, sin högra hand efter arbetshammaren med den slog hon Sisera och krossade hans huvud, spräckte hans tinning och genomborrade den.
Vid hennes fötter sjönk han ihop, föll omkull och blev liggande; ja, vid hennes fötter sjönk han ihop och föll omkull; där han sjönk ihop, där föll han dödsslagen.
Ut genom fönstret skådade hon och ropade, Siseras moder, ut genom gallret: »Varför dröjer väl hans vagn att komma?
Varför äro de så senfärdiga, hans vagnshästars fötter?»
Då svara de klokaste av hennes hovtärnor, och själv giver hon sig detsamma svaret:
»Förvisso vunno de byte, som de nu utskifta: en flicka, ja, två åt envar av männen, byte av praktvävnader för Siseras räkning, byte av praktvävnader, brokiga tyger; en präktig duk, ja, två brokiga dukar för de fångnas halsar.»
Så må alla dina fiender förgås, o HERRE.
Men de som älska honom må likna solen, när den går upp i hjältekraft.
Och landet hade nu ro i fyrtio år.
Men när Israels barn gjorde vad ont var i HERRENS ögon, gav HERREN dem i Midjans hand, i sju år.
Och Midjans hand blev Israel så övermäktig, att Israels barn till skydd mot Midjan gjorde sig de hålor som nu äro att se i bergen, så ock grottorna och bergfästena.
Så ofta israeliterna hade sått, drogo midjaniterna, amalekiterna och österlänningarna upp emot dem
och lägrade sig där och överföllo dem och fördärvade landets gröda ända fram emot Gasa; de lämnade inga livsmedel kvar i Israel, inga får, oxar eller åsnor.
Ty de drogo ditupp med sin boskap och sina tält och kommo så talrika som gräshoppor; de själva och deras kameler voro oräkneliga.
Och de föllo in i landet för att fördärva det.
Så kom Israel i stort elände genom Midjan; då ropade Israels barn till HERREN.
Och när Israels barn ropade till HERREN för Midjans skull,
sände HERREN en profet till Israels barn.
Denne sade till dem: »Så säger HERREN, Israels Gud: Jag själv har fört eder upp ur Egypten och hämtat eder ut ur träldomshuset.
Jag har räddat eder från egyptiernas hand och från alla edra förtryckares hand; jag har förjagat dem för eder och givit eder deras land.
Och jag sade till eder: Jag är HERREN, eder Gud; I skolen icke frukta de gudar som dyrkas av amoréerna, i vilkas land I bon.
Men I villen icke höra min röst.
Och HERRENS ängel kom och satte sig under terebinten vid Ofra, som tillhörde abiesriten Joas; dennes son Gideon höll då på att klappa ut vete i vinpressen, för att bärga det undan Midjan.
För honom uppenbarade sig nu HERRENS ängel och sade till honom: »HERREN är med dig, du tappre stridsman.»
Gideon svarade honom: »Ack min herre, om HERREN är med oss, varför har då allt detta kommit över oss?
Och var äro alla hans under, om vilka våra fäder hava förtäljt för oss och sagt: 'Se, HERREN har fört oss upp ur Egypten'?
Nu har ju HERREN förskjutit oss och givit oss i Midjans våld.»
Då vände sig HERREN till honom och sade: »Gå åstad i denna din kraft och fräls Israel ur Midjans våld; se, jag har sänt dig.»
Han svarade honom: »Ack Herre, varmed kan jag frälsa Israel?
Min ätt är ju den oansenligaste i Manasse, och jag själv den ringaste i min faders hus.»
HERREN sade till honom: »Jag vill vara med dig, så att du skall slå Midjan, såsom voro det en enda man.»
Men han svarade honom: »Om jag har funnit nåd för dina ögon, så låt mig få ett tecken att det är du som talar med mig.
Gå icke bort härifrån, förrän jag har kommit tillbaka till dig och hämtat ut min offergåva och lagt fram den för dig.»
Han sade: »Jag vill stanna, till dess du kommer igen.»
Då gick Gideon in och tillredde en killing, så ock osyrat bröd av en efa mjöl; därefter lade han köttet i en korg och hällde spadet i en kruka; sedan bar han ut det till honom under terebinten och satte fram det.
Men Guds ängel sade till honom: Tag köttet och det osyrade brödet, och lägg det på berghällen där, och gjut spadet däröver.»
Och han gjorde så.
Och HERRENS ängel räckte ut staven som han hade i sin hand och rörde med dess ända vid köttet och det osyrade brödet; då kom eld ut ur klippan och förtärde köttet och det osyrade brödet; och därvid försvann HERRENS ängel ur hans åsyn.
Då såg Gideon att det var HERRENS ängel.
Och Gideon sade: »Ve mig, Herre, HERRE, eftersom jag nu har sett HERRENS ängel ansikte mot ansikte!»
Men HERREN sade till honom: »Frid vare med dig, frukta icke; du skall icke dö.»
Då byggde Gideon där ett altare åt HERREN och kallade det HERREN är frid; det finnes kvar ännu i dag i det abiesritiska Ofra.
Den natten sade HERREN till honom: »Tag den tjur som tillhör din fader och den andra sjuåriga tjuren.
Riv sedan ned det Baalsaltare som tillhör din fader, och hugg sönder Aseran som står därinvid.
Bygg därefter upp ett altare åt HERREN, din Gud, överst på denna fasta plats, och uppför det på övligt sätt; tag så den andra tjuren och offra den till brännoffer på styckena av Aseran som du har huggit sönder.»
Då tog Gideon tio av sina tjänare med sig och gjorde såsom HERREN sade sagt till honom.
Men eftersom han fruktade att göra det om dagen, av rädsla för sin faders hus och för männen i staden, gjorde han det om natten.
Bittida följande morgon fingo mannen i staden se att Baals altare låg nedbrutet, att Aseran därinvid var sönderhuggen, och att den andra tjuren hade blivit offrad såsom brännoffer på det nyuppbyggda altaret.
Då sade de till varandra: »Vem har gjort detta?»
Och när de frågade och gjorde efterforskningar, fingo de veta att Gideon, Joas' son, hade gjort det.
Då sade männen i staden till Joas: »För din son hitut, han måste dö; ty han har brutit ned Baals altare, och han har ock huggit sönder Aseran som stod därinvid.»
Men Joas svarade alla som stodo omkring honom: »Viljen I utföra Baals sak, viljen I komma honom till hjälp?
Den som vill utföra hans sak, han skall bliva dödad innan nästa morgon.
Är han Gud, så utföre han själv sin sak, eftersom denne har brutit ned hans altare.
Härav kallade man honom då Jerubbaal, i det man sade: »Baal utföre sin sak mot honom, eftersom han har brutit ned hans altare.»
Och midjaniterna, amalekiterna och österlänningarna hade alla tillhopa församlat sig och gått över floden och lägrat sig i Jisreels dal.
Men Gideon hade blivit beklädd med HERRENS Andes kraft; han stötte i basun, och abiesriterna församlade sig och följde efter honom.
Och han sände omkring budbärare i hela Manasse, så att ock de övriga församlade sig och följde efter honom; likaledes sände han budbärare till Aser, Sebulon och Naftali, och dessa drogo då också upp, de andra till mötes.
Och Gideon sade till Gud: »Om du verkligen vill genom min hand frälsa Israel, såsom du har lovat,
så se nu här: jag lägger denna avklippta ull på tröskplatsen; ifall dagg kommer allenast på ullen, under det att marken eljest överallt förbliver torr, då vet jag att du genom min hand skall frälsa Israel, såsom du har lovat.»
Och det skedde så, ty när han bittida dagen därefter kramade ur ullen, kunde han av den pressa ut så mycket dagg, att en hel skål blev full med vatten.
Men Gideon sade till Gud: »Må din vrede icke upptändas mot mig, därför att jag talar ännu en enda gång.
Låt mig få försöka blott en gång till med ullen: gör nu så, att allenast ullen förbliver torr, under det att dagg kommer eljest överallt på marken.»
Och Gud gjorde så den natten; allenast ullen var torr, men eljest hade dagg kommit överallt på marken.
Bittida följande morgon drog Jerubbaal, det är Gideon, åstad med allt folket som följde honom, och de lägrade sig vid Harodskällan; han hade då midjaniternas läger norr om sig, från Morehöjden ned i dalen.
Men HERREN sade till Gideon: »Folket som har följt dig är för talrikt för att jag skulle vilja giva Midjan i deras hand; ty Israel kunde då berömma sig mot mig och säga: 'Min egen hand har frälst mig.'
Låt därför nu utropa för folket och säga: Om någon fruktar och är rädd, så må han vända tillbaka hem och skynda bort ifrån Gileads berg.»
Då vände tjugutvå tusen man av folket tillbaka, så att allenast tio tusen man stannade kvar.
Men HERREN sade till Gideon: »Folket är ännu för talrikt; för dem ned till vattnet, så skall jag där göra ett urval av dem åt dig.
Den om vilken jag då säger till dig: 'Denne skall gå med dig', han får gå med dig, men var och en om vilken jag säger till dig: 'Denne skall icke gå med dig', han får icke gå med.»
Så förde han då folket ned till vattnet.
Och HERREN sade till Gideon: »Alla som läppja av vattnet, såsom hunden gör, dem skall du ställa för sig, och likaså alla som falla ned på knä för att dricka.»
Då befanns antalet av dem som hade läppjat av vattnet, genom att med handen föra det till munnen, vara tre hundra man; allt det övriga folket hade fallit ned på knä för att dricka vatten.
Och HERREN sade till Gideon: »Med de tre hundra män som hava läppjat av vattnet skall jag frälsa eder och giva Midjan i din hand; allt det andra folket må begiva sig hem, var och en till sitt.»
Då tog hans folk till sig sitt munförråd och sina basuner, därefter lät han alla de andra israeliterna gå hem, var och en till sin hydda; han behöll allenast de tre hundra männen.
Och midjaniternas läger hade han nedanför sig i dalen.
Och HERREN sade den natten till honom: »Stå upp och drag ned i lägret, ty jag har givit det i din hand.
Men om du fruktar för att draga ditned, så må du gå förut med din tjänare Pura ned till lägret
och höra efter, vad man där talar; sedan skall du få mod till att draga ditned och bryta in i lägret.»
Så gick han då med sin tjänare Pura ned till förposterna i lägret.
Och midjaniterna, amalekiterna och alla österlänningarna lågo där i dalen, talrika såsom gräshoppor; och deras kameler voro oräkneliga, talrika såsom sanden på havets strand.
Då nu Gideon kom dit, höll en man just på att förtälja en dröm för en annan.
Han sade: »Jag har nyss haft en dröm.
Jag tyckte att en kornbrödskaka kom rullande in i midjaniternas läger.
Den kom ända fram till tältet och slog emot det, så att det föll, och vände upp och ned på det, och tältet blev så liggande.»
Då svarade den andre och sade: »Detta betyder intet annat än israeliten Gideons, Joas' sons, svärd; Gud har givit Midjan och hela lägret i hans hand.»
När Gideon hörde denna dröm förtäljas och hörde dess uttydning, föll han ned och tillbad.
Därefter vände han tillbaka till Israels läger och sade: »Stån upp, ty HERREN har givit midjaniternas läger i eder hand.
Och han delade sina tre hundra män i tre hopar och gav allasammans basuner i händerna, så ock tomma krukor, med facklor inne i krukorna.
Och han sade till dem: »Sen på mig och gören såsom jag; så snart jag har kommit till utkanten av lägret, skolen I göra såsom jag gör.
När nämligen jag och alla som jag har med mig stöta i basunerna, skolen ock I stöta i basunerna runt omkring hela lägret och ropa: 'För HERREN och för Gideon!'»
Så kommo nu Gideon och de hundra män, som han hade med sig, till utkanten av lägret, när den mellersta nattväkten ingick; och man hade just ställt ut vakterna.
Då stötte de i basunerna och krossade krukorna som de hade i sina händer.
De tre hoparna stötte i basunerna och slogo sönder krukorna; de fattade med vänstra handen i facklorna och med högra handen i basunerna och stötte i dem; och de ropade: »HERRENS och Gideons svärd!»
Men de stodo stilla, var och en på sin plats, runt omkring lägret.
Då begynte alla i lägret att löpa hit och dit och skria och fly.
Och när de stötte i de tre hundra basunerna, vände HERREN den enes svärd mot den andre i hela lägret; och de som voro i lägret flydde ända till Bet-Hasitta, åt Serera till, ända till stranden vid Abel-Mehola, förbi Tabbat.
Och åter församlade sig israeliterna, från Naftali och Aser och från hela Manasse, och förföljde midjaniterna.
Och Gideon hade sänt omkring budbärare i hela Efraims bergsbygd och låtit säga: »Dragen ned mot Midjan och besätten i deras väg vattendragen ända till Bet-Bara, ävensom Jordan.»
Så församlade sig alla Efraims män och besatte vattendragen ända till Bet-Bara, ävensom Jordan.
Och de togo två midjanitiska hövdingar, Oreb och Seeb, till fånga, och dräpte Oreb vid Orebsklippan, och Seeb dräpte de vid Seebspressen, och förföljde så midjaniterna.
Men Orebs och Seebs huvuden förde de över till Gideon på andra sidan Jordan.
Men Efraims män sade till honom: »Huru har du kunnat handla så mot oss?
Varför bådade du icke upp oss, när du drog ut till strid mot Midjan?»
Och de foro häftigt ut mot honom.
Han svarade dem: »Vad har jag då uträttat i jämförelse med eder?
Är icke Efraims efterskörd bättre än Abiesers vinbärgning?
I eder hand var det som Gud gav de midjanitiska hövdingarna Oreb och Seeb.
Vad har jag kunnat uträtta i jämförelse med eder?»
Då han så talade, stillades deras vrede mot honom.
När sedan Gideon kom till Jordan, gick han över jämte de tre hundra män som han hade med sig; och de voro trötta av förföljandet.
Han sade därför till männen i Suckot: »Given några kakor bröd åt folket som följer mig, ty de äro trötta; se, jag är nu i färd med att förfölja Seba och Salmunna, de midjanitiska konungarna.»
Men de överste i Suckot svarade: »Har du då redan Seba och Salmunna i ditt våld, eftersom du fordrar att vi skola giva bröd åt din här?»
Gideon sade »Nåväl; när HERREN, giver Seba och Salmunna i min hand, skall jag söndertröska edert kött med ökentörnen och tistlar.»
Så drog han vidare därifrån upp till Penuel och talade på samma sätt till dem som voro där; och männen i Penuel gåvo honom samma svar som männen i Suckot hade givit.
Då sade han ock till männen i Penuel: »När jag kommer välbehållen tillbaka, skall jag riva ned detta torn.»
Men Seba och Salmunna befunno sig i Karkor och hade sin här hos sig, vid pass femton tusen man, allt som var kvar av österlänningarnas hela här; ty de stupade utgjorde ett hundra tjugu tusen svärdbeväpnade män.
Och Gideon drog upp på karavanvägen, öster om Noba och Jogbeha, och överföll hären, där den låg sorglös i sitt läger.
Och Seba och Salmunna flydde, men han satte efter dem; och han tog de två midjanitiska konungarna Seba och Salmunna till fånga och skingrade hela hären.
När därefter Gideon, Joas' son, vände tillbaka från striden, ned från Hereshöjden,
fick han fatt på en ung man, en av invånarna i Suckot, och utfrågade denne, och han måste skriva upp åt honom de överste i Suckot och de äldste där, sjuttiosju män.
När han sedan kom till männen i Suckot, sade han: »Se här äro nu Seba och Salmunna, om vilka I hånfullt saden till mig: 'Har du redan Seba och Salmunna i ditt våld, eftersom du fordrar att vi skola giva bröd åt dina trötta män?'»
Därefter lät han gripa de äldste i staden och tog ökentörnen och tistlar och lät männen i Suckot få känna dem.
Och tornet i Penuel rev han ned och dräpte männen i staden.
Och till Seba och Salmunna sade han: »Hurudana voro de män som I dräpten på Tabor?»
De svarade: »De voro lika dig; var och en såg ut såsom en konungason.»
Han sade: »Då var det mina bröder, min moders söner.
Så sant HERREN lever: om I haden låtit dem leva, skulle jag icke hava dräpt eder.»
Sedan sade han till Jeter, sin förstfödde: »Stå upp och dräp dem.»
Men gossen drog icke ut sitt svärd, ty han var försagd, eftersom han ännu var allenast en gosse.
Då sade Seba och Salmunna: »Stå upp, du själv, och stöt ned oss; ty sådan mannen är, sådan är ock hans styrka.»
Så stod då Gideon upp och dräpte Seba och Salmunna.
Och han tog för sin räkning de prydnader som sutto på deras kamelers halsar.
Och israeliterna sade till Gideon: »Råd du över oss, och såsom du så ock sedan din son och din sonson; ty du har frälst oss ur Midjans hand.»
Men Gideon svarade dem: »Jag vill icke råda över eder, och min son skall icke heller råda över eder, utan HERREN skall råda över eder.»
Och Gideon sade ytterligare till dem: »Ett vill jag dock begära av eder: var och en av eder må giva mig den näsring han har fått såsom byte.»
Ty midjaniterna buro näsringar av guld, eftersom de voro ismaeliter.
De svarade: »Ja, vi vilja giva dig dem.»
Och de bredde ut ett kläde, och var och en kastade på detta den näsring han hade fått såsom byte.
Och guldringarna, som han hade begärt, befunnos väga ett tusen sju hundra siklar i guld -- detta förutom de halsprydnader, de örhängen och de purpurröda kläder som de midjanitiska konungarna hade burit, och förutom de kedjor som hade suttit på deras kamelers halsar.
Och Gideon lät därav göra en efod och satte upp den i sin stad, Ofra; och hela Israel lopp där i trolös avfällighet efter den.
Och den blev för Gideon och hans hus till en snara.
Så blev nu Midjan kuvat under Israels barn och upplyfte icke mer sitt huvud.
Och landet hade ro i fyrtio år, så länge Gideon levde.
Men Jerubbaal, Joas' son, gick hem och stannade sedan i sitt hus.
Och Gideon hade sjuttio söner, som hade utgått från hans länd, ty han ägde många hustrur.
En bihustru som han hade i Sikem födde honom ock en son; denne gav han namnet Abimelek.
Och Gideon, Joas' son, dog i en god ålder och blev begraven i sin fader Joas' grav i det abiesritiska Ofra
Men när Gideon var död, begynte Israels barn åter i trolös avfällighet löpa efter Baalerna; och de gjorde Baal-Berit till gud åt sig.
Israels barn tänkte icke på HERREN, sin Gud, som hade räddat dem från alla deras fienders hand runt omkring.
Ej heller visade de Jerubbaals, Gideons, hus någon kärlek, till gengäld för allt det goda som han hade gjort mot Israel.
Men Abimelek, Jerubbaals son, gick bort till sin moders bröder i Sikem och talade till dem och till alla som voro besläktade med hans morfaders hus, och sade:
»Talen så till alla Sikems borgare: Vilket är bäst för eder: att sjuttio män, alla Jerubbaals söner, råda över eder, eller att en enda man råder över eder?
Kommen därjämte ihåg att jag är edert kött och ben.»
Då talade hans moders bröder till hans förmån allt detta inför alla Sikems borgare.
Och dessa blevo vunna för Abimelek, ty de tänkte: »Han är ju vår broder.»
Och de gåvo honom sjuttio siklar silver ur Baal-Berits tempel; för dessa lejde Abimelek löst folk och äventyrare, vilkas anförare han blev.
Därefter begav han sig till sin faders hus i Ofra och dräpte där sina bröder, Jerubbaals söner, sjuttio män, och detta på en och samma sten; dock blev Jotam, Jerubbaals yngste son, vid liv, ty han hade gömt sig.
Sedan församlade sig alla Sikems borgare och alla som bodde i Millo och gingo åstad och gjorde Abimelek till konung vid Vård-terebinten invid Sikem.
När man berättade detta far Jotam, gick han åstad och ställde sig på toppen av berget Gerissim och hov upp sin röst och ropade och sade till dem: »Hören mig, I Sikems borgare, för att Gud ock må höra eder.
Träden gingo en gång åstad för att smörja en konung över sig.
Och de sade till olivträdet: 'Bliv du konung över oss'
Men olivträdet svarade dem: 'Skulle jag avstå från min fetma, som både gudar och människor ära mig för, och gå bort för att svaja över de andra träden?'
Då sade träden till fikonträdet: 'Kom du och bliv konung över oss.'
Men fikonträdet svarade dem: 'Skulle jag avstå från min sötma och min goda frukt och gå bort för att svaja över de andra träden?'
Då sade träden till vinträdet: 'Kom du och bliv konung över oss.'
Men vinträdet svarade dem: 'Skulle jag avstå från min vinmust, som gör både gudar och människor glada, och gå bort för att svaja över de andra träden?'
Då sade alla träden till törnbusken: 'Kom du och bliv konung över oss.'
Törnbusken svarade träden: 'Om det är eder uppriktiga mening att smörja mig till konung över eder, så kommen och tagen eder tillflykt under min skugga; varom icke, så skall eld gå ut ur törnbusken och förtära cedrarna på Libanon.'
Så hören nu: om I haven förfarit riktigt och redligt däri att I haven gjort Abimelek till konung, och om I haven förfarit väl mot Jerubbaal och hans hus, och haven vedergällt honom efter hans gärningar --
ty I veten att min fader stridde för eder och vågade sitt liv för att rädda eder från Midjans hand,
under det att I däremot i dag haven rest eder upp mot min faders hus och dräpt hans söner, sjuttio män, på en och samma sten, och gjort Abimelek, hans tjänstekvinnas son, till konung över Sikems borgare, eftersom han är eder broder --
om I alltså denna dag haven förfarit riktigt och redligt mot Jerubbaal och hans hus, då mån I glädja eder över Abimelek, och han må ock glädja sig över eder;
varom icke, så må eld gå ut från Abimelek och förtära Sikems borgare och dem som bo i Millo, och från Sikems borgare och från dem som bo i Millo må eld gå ut och förtära Abimelek.»
Och Jotam skyndade sig undan och flydde bort till Beer, och där bosatte han sig för att vara i säkerhet för sin broder Abimelek.
När Abimelek hade härskat över Israel i tre år,
sände Gud en tvedräktsande mellan Abimelek och Sikems borgare, så att Sikems borgare avföllo från Abimelek.
Detta skedde, för att våldet mot Jerubbaals sjuttio söner skulle bliva hämnat, och för att deras blod skulle komma över deras broder Abimelek som dräpte dem, så ock över Sikems borgare, som lämnade honom understöd, så att han kunde dräpa sina bröder.
För att skada honom lade Sikems borgare nu folk i försåt på bergshöjderna, och dessa plundrade alla som drogo vägen fram därförbi.
Detta blev berättat för Abimelek.
Men Gaal, Ebeds son, kom nu dit med sina bröder, och de drogo in i Sikem.
Och Sikems borgare fattade förtroende för honom.
Så hände sig en gång att de gingo ut på fältet och avbärgade sina vingårdar och pressade druvorna och höllo en glädjefest, och de gingo därvid in i sin guds hus och åto och drucko, och uttalade förbannelser över Abimelek.
Och Gaal, Ebeds son, sade: »Vad är Abimelek, och vad är Sikem, eftersom vi skola tjäna honom?
Han är ju Jerubbaals son, och Sebul är hans tillsyningsman.
Nej, tjänen män som härstamma från Hamor, Sikems fader.
Varför skulle vi tjäna denne?
Ack om jag hade detta folk under min vård!
Då skulle jag driva bort Abimelek.»
Och i fråga om Abimelek sade han: »Föröka din här och drag ut.»
Men när Sebul, hövitsmannen i staden, fick höra vad Gaal, Ebeds son, hade sagt, upptändes hans vrede.
Och han sände listeligen bud till Abimelek och lät säga: »Se, Gaal, Ebeds son, och hans bröder hava kommit till Sikem, och de hålla just nu på att uppvigla staden mot dig.
Bryt därför nu upp om natten, du med ditt folk, och lägg dig i bakhåll på fältet.
Sedan må du i morgon bittida, när solen går upp, störta fram mot staden.
När han då med sitt folk drager ut mot dig, må du göra med honom vad tillfället giver vid handen.»
Då bröt Abimelek med allt sitt folk upp om natten, och de lade sig i bakhåll mot Sikem, i fyra hopar.
Och Gaal, Ebeds son, kom ut och ställde sig vid ingången till stadsporten; och i detsamma bröt Abimelek med sitt folk fram ifrån bakhållet.
När då Gaal såg folket, sade han till Sebul: »Se, där kommer folk ned från bergshöjderna.»
Men Sebul svarade honom: »Det är skuggan av bergen, som för dina ögon ser ut såsom människor.»
Gaal tog åter till orda och sade: »Jo, där kommer folk ned från Mittelhöjden, och en annan hop kommer på vägen från Teckentydarterebinten.»
Då sade Sebul till honom: »Var är nu din stortalighet, du som sade: 'Vad är Abimelek, eftersom vi skola tjäna honom?'
Se, här kommer det folk som du så föraktade.
Drag nu ut och strid mot dem.
Så drog då Gaal ut i spetsen för Sikems borgare och gav sig i strid med Abimelek.
Men Abimelek jagade honom på flykten, och han flydde undan för honom; och många föllo slagna ända fram till stadsporten.
Och Abimelek stannade i Aruma; men Sebul drev bort Gaal och hans bröder och lät dem icke längre stanna i Sikem.
Dagen därefter gick folket ut på fältet; och man berättade detta för Abimelek.
Då tog han sitt folk och delade dem i tre hopar och lade sig i bakhåll på fältet.
Och när han fick se att folket gick ut ur staden, bröt han upp och anföll dem och nedgjorde dem.
Abimelek och de hopar han hade med sig störtade nämligen fram och ställde sig vid ingången till stadsporten; men de båda andra hoparna störtade fram mot alla som voro på fältet och nedgjorde dem.
När så Abimelek hade ansatt staden hela den dagen, intog han den och dräpte det folk som fanns därinne Sedan rev han ned staden och beströdde platsen med salt.
När besättningen i Sikems torn hörde detta, begåvo de sig alla till det fasta valvet i El-Berits tempelbyggnad.
Och när det blev berättat for Abimelek att hela besättningen i Sikems torn hade församlat sig där,
gick han med allt sitt folk upp till berget Salmon; och Abimelek tog en yxa i sin hand och högg av en trädgren och lyfte upp den och lade den på axeln; och han sade till sitt folk: »Gören med hast detsamma som I haven sett mig göra.»
Då högg också allt folket av var sin gren och följde efter Abimelek, och de lade grenarna intill det fasta valvet och tände upp eld till att förbränna valvet jämte dem som voro där.
Så omkommo ock alla de människor som bodde i Sikems torn, vid pass tusen män och kvinnor.
Och Abimelek drog åstad till Tebes och belägrade Tebes och intog det.
Men mitt i staden var ett starkt torn, och dit flydde alla män och kvinnor, alla borgare i staden, och stängde igen om sig; sedan stego de upp på tornets tak.
Och Abimelek kom till tornet och angrep det; och han gick fram till porten på tornet för att bränna upp den i eld.
Men en kvinna kastade en kvarnsten ned på Abimeleks huvud och bräckte så hans huvudskål.
Då ropade han med hast på sin vapendragare och sade till honom: »Drag ut ditt svärd och döda mig, för att man icke må säga om mig: En kvinna dräpte honom.»
Då genomborrade hans tjänare honom, så att han dog.
När nu israeliterna sågo att Abimelek var död, gingo de hem, var och en till sitt.
Alltså lät Gud det onda som Abimelek hade gjort mot sin fader, då han dräpte sina sjuttio bröder, komma tillbaka över honom.
Och allt det onda som Sikems män hade gjort lät Gud ock komma tillbaka över deras huvuden.
Så gick Jotams, Jerubbaals sons, förbannelse i fullbordan på dem.
Efter Abimelek uppstod till Israels frälsning Tola, son till Pua, son till Dodo, en man från Isaskar; och han bodde i Samir, i Efraims bergsbygd.
Han var domare i Israel i tjugutre år; sedan dog han och blev begraven i Samir.
Efter honom uppstod gileaditen Jair.
Han var domare i Israel i tjugutvå år.
Han hade trettio söner, som plägade rida på trettio åsnor; och de hade trettio städer.
Dessa kallar man ännu i dag Jairs byar, och de ligga i Gileads land.
Och Jair dog och blev begraven i Kamon.
Men Israels barn gjorde åter vad ont var i HERRENS ögon och tjänade Baalerna och Astarterna, så ock Arams, Sidons, Moabs, Ammons barns och filistéernas gudar och övergåvo HERREN och tjänade honom icke.
Då upptändes HERRENS vrede mot Israel, och han sålde dem i filistéernas och Ammons barns hand.
Och dessa plågade Israels barn och förforo våldsamt mot dem det året; i aderton år gjorde de så mot alla de israeliter som bodde på andra sidan Jordan, i amoréernas land, i Gilead.
Därtill gingo Ammons barn över Jordan och gåvo sig i strid också med Juda, Benjamin och Efraims hus, så att Israel kom i stor nöd.
Då ropade Israels barn till HERREN och sade: »Vi hava syndat mot dig, ty vi hava övergivit vår Gud och tjänat Baalerna.»
Men HERREN sade till Israels barn: »Har jag icke frälst eder från egyptierna, amoréerna, Ammons barn och filistéerna?
Likaledes bleven I förtryckta av sidonierna, amalekiterna och maoniterna; och när I ropaden till mig, frälste jag eder från deras hand.
Men I haven nu övergivit mig och tjänat andra gudar; därför vill jag icke mer frälsa eder.
Gån bort och ropen till de gudar som I haven utvalt; må de frälsa eder, om I nu ären i nöd.
Då sade Israels barn till HERREN: »Vi hava syndat; gör du med oss alldeles såsom dig täckes.
Allenast rädda oss nu denna gång.»
Därefter skaffade de bort ifrån sig de främmande gudarna och tjänade HERREN.
Då kunde han icke längre lida att se Israels vedermöda.
Och Ammons barn blevo uppbådade och lägrade sig i Gilead; men Israels barn församlade sig och lägrade sig i Mispa.
Då sade folket, nämligen de överste i Gilead, till varandra: »Vem vill begynna striden mot Ammons barn?
Den som det vill skall bliva hövding över alla Gileads inbyggare.»
Gileaditen Jefta var en tapper stridsman, men han var son till en sköka; och Jeftas fader var Gilead.
Nu födde ock Gileads hustru honom söner; och när dessa hans hustrus söner hade växt upp, drevo de ut Jefta och sade till honom: »Du skall icke taga arv i vår faders hus, ty du är son till en kvinna som icke är hans hustru.»
Då flydde Jefta bort ifrån sina bröder och bosatte sig i landet Tob; där sällade sig löst folk till Jefta och gjorde strövtåg med honom.
Någon tid därefter gåvo Ammons barn sig i strid med Israel.
Men när Ammons barn gåvo sig i strid med Israel, gingo de äldste i Gilead åstad för att hämta Jefta från landet Tob.
Och de sade till Jefta: »Kom och bliv vår anförare, så vilja vi strida mot Ammons barn.»
Men Jefta svarade de äldste i Gilead: »I haven ju hatat mig och drivit mig ut ur min faders hus.
Huru kunnen I då nu, när I ären i nöd, komma till mig?»
De äldste i Gilead sade till Jefta: »Just därför hava vi nu kommit tillbaka till dig, och du måste gå med oss och strida mot Ammons barn; ty du skall bliva hövding över oss, alla Gileads inbyggare.»
Jefta svarade de äldste i Gilead: »Om I nu fören mig tillbaka för att strida mot Ammons barn och HERREN giver dem i mitt våld, så vill jag ock sedan vara eder hövding.»
Då sade de äldste i Gilead till Jefta: »HERREN höre vårt avtal.
Förvisso skola vi låta det bliva så om du har sagt.»
Så gick då Jefta med de äldste i Gilead, och folket satte honom till hövding och anförare över sig.
Och Jefta uttalade inför HERREN i Mispa allt vad han hade sagt.
Och Jefta skickade sändebud till Ammons barns konung och lät säga: »Vad har du med mig att göra, eftersom du har kommit emot mig och angripit mitt land?»
Då svarade Ammons barns konung Jeftas sändebud: »När Israel drog upp från Egypten, togo de ju mitt land från Arnon ända till Jabbok och till Jordan; så giv mig nu detta tillbaka i godo.»
Åter skickade Jefta sändebud till Ammons barns konung
och lät säga till honom: »Så säger Jefta: Israel har icke tagit något land vare sig från Moab eller från Ammons barn.
Ty när de drogo upp från Egypten och Israel hade tågat genom öknen ända till Röda havet och sedan kommit till Kades,
skickade Israel sändebud till konungen i Edom och lät säga: 'Låt mig tåga genom ditt land.'
Men konungen i Edom hörde icke därpå.
De skickade ock till konungen i Moab, men denne ville icke heller Då stannade Israel i Kades.
Därefter tågade de genom öknen och gingo omkring Edoms land och Moabs land och kommo öster om Moabs land och lägrade sig på andra sidan Arnon; de kommo icke in på Moabs område, ty Arnon är Moabs gräns.
Sedan skickade Israel sändebud till Sihon, amoréernas konung, konungen i Hesbon; och Israel lät säga till honom: 'Låt oss genom ditt land tåga dit vi skola.'
Men Sihon litade icke på Israel och lät dem icke tåga genom sitt land, utan församlade allt sitt folk, och de lägrade sig i Jahas; där in- lät han sig i strid med Israel.
Men HERREN, Israels Gud, gav Sihon och allt hans folk i Israels hand, så att de slogo dem; och Israel intog hela amoréernas land, ty dessa bodde då i detta land.
De intogo hela amoréernas område, från Arnon ända till Jabbok, och från öknen ända till Jordan.
Och nu, då HERREN, Israels Gud, har fördrivit amoréerna för sitt folk Israel, skulle du taga deras land i besittning!
Är det icke så: vad din gud Kemos giver dig till besittning, det tager du i besittning?
Så taga ock vi, närhelst HERREN, vår Gud, fördriver ett folk för oss, deras land i besittning.
Menar du att du är så mycket förmer än Balak, Sippors sons konungen i Moab?
Han dristade ju icke att inlåta sig i tvist med Israel eller giva sig i strid med dem.
När Israel nu i tre hundra år har bott i Hesbon och underlydande orter, i Aror och underlydande orter och i alla städer på båda sidor om Arnon, varför haven I då under hela den tiden icke tagit detta ifrån oss?
Jag har icke försyndat mig mot dig, men du gör illa mot mig, då du nu överfaller mig.
HERREN, domaren, må i dag döma mellan Israels barn och Ammons barn.»
Men Ammons barns konung hörde icke på vad Jefta lät säga honom genom sändebuden.
Då kom HERRENS Ande över Jefta; och han tågade genom Gilead och Manasse och tågade så genom Mispe i Gilead, och från Mispe i Gilead tågade han fram mot Ammons barn.
Och Jefta gjorde ett löfte åt HERREN och sade: »Om du giver Ammons barn i min hand,
så lovar jag att vadhelst som ur dörrarna till mitt hus går ut emot mig, när jag välbehållen kommer tillbaka från Ammons barn, det skall höra HERREN till, och det skall jag offra till brännoffer.»
Så drog nu Jefta åstad mot Ammons barn för att strida mot dem; och HERREN gav dem i hans hand.
Och han tillfogade dem ett mycket stort nederlag och intog landet från Aroer ända till fram emot Minnit, tjugu städer, och ända till Abel-Keramim.
Alltså blevo Ammons barn kuvade under Israels barn.
När sedan Jefta kom hem till sitt hus i Mispa, då gick hans dotter ut emot honom med pukor och dans.
Och hon var hans enda barn, han hade utom henne varken son eller dotter.
I detsamma han nu fick se henne, rev han sönder sina kläder och ropade: »Ve mig, min dotter, du kommer mig att sjunka till jorden, du drager olycka över mig!
Ty jag har öppnat min mun inför HERREN till ett löfte och kan icke taga mitt ord tillbaka.»
Hon svarade honom: »Min fader, har du öppnat din mun inför HERREN, så gör med mig enligt din muns tal, eftersom HERREN nu har skaffat dig hämnd på dina fiender, Ammons barn.»
Och hon sade ytterligare till sin fader: »Uppfyll dock denna min begäran: unna mig två månader, så att jag får gå åstad ned på bergen och begråta min jungfrudom med mina väninnor.
Han svarade: »Du får gå åstad.»
Och han tillstadde henne att vara borta i två månader.
Då gick hon åstad med sina väninnor och begrät sin jungfrudom på bergen.
Men efter två månader vände hon tillbaka till sin fader, och han förfor då med henne efter det löfte han hade gjort.
Och hon hade icke känt någon man.
Sedan blev det en sedvänja i Israel att Israels döttrar år efter år gingo åstad för att lovprisa gileaditen Jeftas dotter, under fyra dagar vart år.
Men Efraims män församlade sig och drogo till Safon; och de sade till Jefta: »Varför drog du åstad till strid mot Ammons barn utan att kalla på oss till att tåga med dig?
Nu vilja vi bränna upp ditt hus jämte dig själv i eld.
Jefta svarade dem: »Jag och mitt folk lågo i svår fejd med Ammons barn; då manade jag eder att komma, men I villen icke frälsa mig ur deras hand.
Och när jag såg att I icke villen frälsa mig, tog jag min själ i min hand och drog åstad mot Ammons barn, och HERREN gav dem i min hand.
Varför haven I då nu dragit upp emot mig till att strida emot mig?»
Och Jefta församlade alla Gileads män och gav sig i strid med Efraim.
Och Gileads män slogo efraimiterna; dessa hade nämligen sagt: »Flyktingar ifrån Efraim ären I; Gilead är ett mellanting, varken Efraim eller Manasse.»
Och gileaditerna besatte vadställena över Jordan för efraimiterna.
Då nu någon av de efraimitiska flyktingarna sade: »Låt mig komma över», frågade Gileads män honom: »Är du en efraimit?»
Om han då svarade nej,
så sade de till honom: »Säg 'schibbolet'.»
Sade han då »sibbolet», därför att han icke nog lade sig vinn om att uttala ordet rätt, så grepo de honom och höggo ned honom där vid vadställena över Jordan.
På detta sätt föllo vid det tillfället fyrtiotvå tusen efraimiter.
Och Jefta var domare i Israel i sex år.
Sedan dog gileaditen Jefta och blev begraven i en av Gileads städer.
Efter honom var Ibsan från Bet-Lehem domare i Israel.
Han hade trettio söner, och trettio döttrar gifte han bort; han fick ock trettio döttrar genom att skaffa hustrur åt sina söner utifrån.
Och han var domare i Israel i sju år.
Sedan dog Ibsan och blev begraven i Bet-Lehem.
Efter honom var sebuloniten Elon domare i Israel; i tio år var han domare i Israel.
Sedan dog sebuloniten Elon och blev begraven i Ajalon, i Sebulons land.
Efter honom var pirgatoniten Abdon, Hillels son, domare i Israel.
Han hade fyrtio söner och trettio sonsöner, vilka plägade rida på sjuttio åsnor.
Och han var domare i Israel i åtta år.
Sedan dog pirgatoniten Abdon, Hillels son, och blev begraven i Pirgaton i Efraims land, i amalekiternas bergsbygd.
Men Israels barn gjorde åter vad ont var i HERRENS ögon; då gav HERREN dem i filistéernas hand, i fyrtio år.
I Sorga levde nu en man av daniternas släkt, vid namn Manoa; hans hustru var ofruktsam och hade icke fött några barn.
Men HERRENS ängel uppenbarade sig för hustrun och sade till henne: »Se, du är ofruktsam och har icke fött några barn, men du skall bliva havande och föda en son.
Tag dig nu till vara, så att du icke dricker vin eller starka drycker ej heller äter något orent.
Ty se, du skall bliva havande och föda en son, på vilkens huvud ingen rakkniv skall komma, ty gossen skall vara en Guds nasir allt ifrån moderlivet; och han skall göra begynnelse till att frälsa Israel ur filistéernas hand.»
Då gick hustrun in och omtalade detta för sin man och sade: »En gudsman kom till mig; han såg ut såsom en Guds ängel, mycket fruktansvärd.
Jag frågade honom icke varifrån han var, och sitt namn lät han mig icke veta.
Och han sade till mig: 'Se, du skall bliva havande och föda en son; drick nu icke vin eller starka drycker och ät icke något orent, ty gossen skall vara en Guds nasir, från moderlivet ända till sin död.'»
Och Manoa bad till HERREN och sade: »Ack Herre, låt gudsmannen som du sände hit åter komma till oss, för att han må lära oss huru vi skola göra med gossen som skall födas.»
Och Gud hörde Manoas röst; Guds ängel kom åter till hans hustru, när hon en gång satt ute på marken och hennes man Manoa icke var hos henne.
Då skyndade hustrun strax åstad och berättade det för sin man; hon sade till honom: »Mannen som kom till mig häromdagen har uppenbarat sig för mig.»
Manoa stod upp och följde sin hustru; och när han kom till mannen, frågade han honom: »Är du den man som förut talade med min hustru?»
Han svarade: »Ja.»
Då sade Manoa: »När det som du har sagt går i fullbordan, vad är då att iakttaga med gossen?
Hur skall man göra med honom?»
HERRENS ängel svarade Manoa »Din hustru skall taga sig till vara för allt varom jag har talat med henne.
Hon skall icke äta något som ha vuxit på vinträd, och vin eller starka drycker får hon icke dricka, ej heller får hon äta något orent.
Allt vad jag har bjudit henne skall hon hålla.»
Och Manoa sade till HERRENS ängel: »Låt oss få hålla dig kvar, så vilja vi tillreda en killing och sätta fram för dig.»
Men HERRENS ängel svarade Manoa: »Om du ock håller mig kvar, skall jag dock icke äta av din mat; men om du vill tillreda ett brännoffer, så offra detta åt HERREN.»
Ty Manoa förstod icke att det var HERRENS ängel.
Och Manoa sade till HERRENS ängel: »Vad är ditt namn?
Säg oss det, för att vi må kunna ära dig, när det som du har sagt går i fullbordan.»
HERRENS ängel sade till honom: »Varför frågar du efter mitt namn?
Det är alltför underbart.»
Och Manoa tog killingen med tillhörande spisoffer och lade upp den på klippan åt HERREN.
Då lät han något underbart ske i Manoas och hans hustrus åsyn.
När lågan steg upp från altaret mot himmelen, for nämligen HERRENS ängel upp, i lågan från altaret.
Då Manoa och hans hustru sågo detta, föllo de ned till jorden på sitt ansikte
Sedan visade sig HERRENS ängel icke mer för Manoa och hans hustru.
Då förstod Manoa att det hade varit HERRENS ängel.
Och Manoa sade till sin hustru: »Nu måste vi dö, eftersom vi hava sett Gud.»
Men hans hustru svarade honom: »Om HERREN hade velat döda oss, så hade han icke tagit emot något brännoffer och spisoffer av vår hand, och icke låtit oss se allt detta, ej heller hade han nu låtit oss höra sådant.»
Därefter födde hans hustru en son och gav honom namnet Simson; och gossen växte upp, och HERREN välsignade honom.
Och HERRENS Ande begynte att verka på honom, medan han var i Dans läger, mellan Sorga och Estaol.
När Simson en gång gick ned till Timna, fick han där i Timna se en kvinna, en av filistéernas döttrar.
Och när han kom upp därifrån, omtalade han det för sin fader och moder och sade: »Jag har i Timna sett en kvinna, en av filistéernas döttrar; henne mån I nu skaffa mig till hustru.»
Hans fader och moder sade till honom: »Finnes då ingen kvinna bland dina bröders döttrar och i hela mitt folk, eftersom du vill gå bort för att skaffa dig en hustru från de oomskurna filistéerna?»
Simson sade till sin fader: »Skaffa mig denna, ty hon behagar mig.»
Men hans fader och moder visste icke att detta kom från HERREN, som sökte sak med filistéerna.
På den tiden rådde nämligen filistéerna över Israel.
Och Simson gick med sin fader och moder ned till Timna; men just som de hade hunnit fram till vingårdarna vid Timna, kom ett ungt lejon rytande emot honom.
Då föll HERRENS Ande över honom, och han slet sönder lejonet, såsom hade han slitit sönder en killing, fastän han icke hade någonting i sin hand; men han talade icke om för sin fader och moder vad han hade gjort.
När han så kom ditned, talade han med kvinnan; och hon behagade Simson.
En tid därefter vände han tillbaka för att hämta henne och vek då av vägen för att se på det döda lejonet; då fick han i lejonets kropp se en bisvärm med honung.
Och han skrapade ut honungen i sina händer och åt därav, medan han gick, han kom så till sin fader och moder och gav dem, och de åto.
Men han talade icke om för dem att det var ur lejonets kropp han hade skrapat honungen.
När nu hans fader kom ned till kvinnan, gjorde Simson där ett gästabud, ty så plägade de unga männen göra.
Och när de fingo se honom, skaffade de trettio bröllopssvenner, som skulle vara hos honom.
Till dem sade Simson: »Jag vill förelägga eder en gåta; om I under de sju gästabudsdagarna sägen mig lösningen på den och gissen rätt, så skall jag giva eder trettio fina linneskjortor och trettio högtidsdräkter.
Men om I icke kunnen säga mig lösningen, så skolen I giva mig trettio fina linneskjortor och trettio högtidsdräkter.»
De sade till honom: »Förelägg oss din gåta, låt oss höra den.»
Då sade han till dem: »Från storätaren utgick ätbart, från den grymme kom sötma.»
Men under tre dagar kunde de icke lösa gåtan.
På sjunde dagen sade de då till Simsons hustru: »Locka din man till att säga oss lösningen på gåtan; eljest skola vi bränna upp dig och din faders hus i eld.
Icke haven I väl bjudit oss hit för att utarma oss?»
Då låg Simsons hustru över honom med gråt och sade: »Du hatar mig allenast och älskar mig alls icke; du har förelagt mina landsmän en gåta, men mig har du icke sagt lösningen på den.»
Han svarade henne: »Icke ens åt min fader eller min moder har jag sagt lösningen; skulle jag då säga den åt dig?»
Men hon låg över honom med gråt under de sju dagar de höllo gästabudet.
Och på sjunde dagen sade han henne lösningen, eftersom hon så hårt ansatte honom; sedan sade hon lösningen på gåtan åt sina landsmän.
Innan solen gick ned på sjunde dagen, gåvo honom alltså männen i staden det svaret: »Vad är sötare än honung, och vad är grymmare än ett lejon?»
Men han sade till dem: »Haden I icke plöjt med min kviga, så haden I icke gissat min gåta.»
Och HERRENS Ande kom över honom, och han gick ned till Askelon och slog där ihjäl trettio män och tog deras kläder och gav högtidsdräkterna åt dem som hade sagt lösningen på gåtan.
Och hans vrede upptändes, och han vände tillbaka upp till sin faders hus.
Då blev Simsons hustru given åt den av hans bröllopssvenner, som han hade haft till sin särskilda följesven.
En tid därefter, medan veteskörden pågick, ville Simson besöka sin hustru, och förde med sig en killing.
Och han sade: »Låt mig gå in till min hustru i kammaren.»
Men hennes fader ville icke tillstädja honom att gå in;
hennes fader sade: »Jag höll för säkert att du hade fattat hat till henne, och därför gav jag henne åt din bröllopssven.
Men hon har ju en yngre syster, som är fagrare än hon; tag denna i stället för den andra.»
Men Simson svarade dem: »Denna gång är jag utan skuld gent emot filistéerna, om jag gör dem något ont.»
Och Simson gick bort och fångade tre hundra rävar; sedan tog han facklor, band så ihop två och två rävar med svansarna och satte in en fackla mitt emellan de två svansarna.
Därefter tände han eld på facklorna och släppte djuren in på filistéernas sädesfält och antände så både sädesskylar och oskuren säd, vingårdar och olivplanteringar.
Då nu filistéerna frågade efter vem som hade gjort detta, fingo de det svaret: »Det har Simson, timnitens måg, därför att denne tog hans hustru och gav henne åt hans bröllopssven.»
Då drogo filistéerna åstad och brände upp både henne och hennes fader i eld.
Men Simson sade till dem: »Om I beten eder så, skall jag sannerligen icke vila, förrän jag har tagit hämnd på eder.»
Och han for våldsamt fram med dem, så att de varken kunde gå eller stå.
Sedan gick han ned därifrån och bodde i bergsklyftan vid Etam.
Då drogo filistéerna upp och lägrade sig i Juda; och de spridde sig i Lehi.
Och Juda män sade: »Varför haven I dragit hitupp mot oss?»
De svarade: »Vi hava dragit hitupp för att binda Simson och för att göra mot honom såsom han har gjort mot oss.»
Då drogo tre tusen män från Juda ned till bergsklyftan vid Etam och sade till Simson: »Du vet ju att filistéerna råda över oss; huru har du då kunnat göra så mot oss?»
Han svarade dem: »Såsom de hava gjort mot mig, så har jag gjort mot dem.»
De sade till honom: »Vi hava kommit hitned för att binda dig och sedan lämna dig i filistéernas hand.»
Simson sade till dem: »Så given mig nu eder ed på att I icke själva viljen stöta ned mig.»
De svarade honom: »Nej, vi vilja allenast binda dig och sedan lämna dig i deras hand, men vi skola icke döda dig.»
Så bundo de honom med två nya tåg och förde honom upp, bort ifrån klippan.
När han nu kom till Lehi, skriade filistéerna och sprungo emot honom.
Då kom HERRENS Ande över honom, och tågen omkring hans armar blevo såsom lintrådar, när de antändas av eld, och banden likasom smälte bort ifrån hans händer.
Och han fick fatt i en åsnekäke som ännu var frisk; och han räckte ut sin hand och tog den, och med den slog han ihjäl tusen män.
Sedan sade Simson: »Med åsnekäken slog jag en skara, ja, två; med åsnekäken slog jag tusen man.»
När han hade sagt detta, kastade han käken ifrån sig.
Och man kallade den platsen Ramat-Lehi .
Men då han därefter blev mycket törstig, ropade han till HERREN och sade: »Du själv har genom din tjänare givit denna stora seger; och nu måste jag dö av törst, och så falla i de oomskurnas hand!»
Då lät Gud fördjupningen i Lehi öppna sig, och därur gick ut vatten, så att han kunde dricka; och hans ande kom tillbaka, och han fick liv igen.
Därav kallades källan Den ropandes källa i Lehi , såsom den heter ännu i dag.
Och han var domare i Israel under filistéernas tid, i tjugu år.
Och Simson gick till Gasa; där fick han se en sköka och gick in till henne.
När då gasiterna fingo höra att Simson hade kommit dit, omringade de platsen och lågo i försåt för honom hela natten vid stadsporten.
Men hela natten höllo de sig stilla; de tänkte: »Vi vilja vänta till i morgon, när det bliver dager; då skola vi dräpa honom.»
Och Simson låg där intill midnatt; men vid midnattstiden stod han upp och grep tag i stadsportens dörrar och i de båda dörrposterna och ryckte loss dem jämte bommen, och lade alltsammans på sina axlar och bar upp det till toppen på det berg som ligger gent emot Hebron.
Därefter fattade han kärlek till en kvinna som hette Delila, vid bäcken Sorek.
Då kommo filistéernas hövdingar upp till henne och sade till henne: »Locka honom till att uppenbara för dig varav det beror att han är så stark, och huru vi skola bliva honom övermäktiga, så att vi kunna binda honom och kuva honom; vi vilja då giva dig ett tusen ett hundra siklar silver var.»
Då sade Delila till Simson: »Säg mig varav det beror att du är så stark, och huru man skulle kunna binda och kuva dig.»
Simson svarade henne: »Om man bunde mig med sju friska sensträngar, som icke hade hunnit torka, så bleve jag svag och vore såsom en vanlig människa.»
Då buro filistéernas hövdingar till henne sju friska sensträngar, som icke hade hunnit torka; och hon band honom med dem.
Men hon hade lagt folk i försåt i den inre kammaren.
Sedan ropade hon till honom: »Filistéerna äro över dig, Simson!»
Då slet han sönder sensträngarna så lätt som en blångarnssnodd slites sönder, när den kommer intill elden.
Alltså hade man ingenting fått veta om hans styrka.
Då sade Delila till Simson: »Du har ju bedragit mig och ljugit för mig.
Men säg mig nu huru man skulle kunna binda dig.»
Han svarade henne: »Om man bunde mig med nya tåg, som ännu icke hade blivit begagnade till något, så bleve jag svag och vore såsom en vanlig människa.»
Då tog Delila nya tåg och band honom med dem och ropade så till honom: »Filistéerna äro över dig, Simson!»; och folk låg i försåt i den inre kammaren.
Men han slet tågen av sina armar, såsom hade det varit trådar.
Då sade Delila till Simson: »Hittills har du bedragit mig och ljugit för mig; säg mig nu huru man skulle kunna binda dig.»
Han svarade henne: »Jo, om du vävde in de sju flätorna på mitt huvud i ränningen till din väv.»
Hon slog alltså fast dem med pluggen och ropade sedan till honom: »Filistéerna äro över dig, Simson!»
När han då vaknade upp ur sömnen, ryckte han loss vävpluggen jämte ränningen till väven.
Då sade hon till honom: »Huru kan du säga att du har mig kär, du som icke är uppriktig mot mig?
Tre gånger har du nu bedragit mig och icke velat säga mig varpå det beror att du är så stark.»
Då hon nu dag efter dag hårt ansatte honom med denna sin begäran och plågade honom därmed, blev han så otålig att han kunde dö,
och yppade så för henne hela sin hemlighet och sade till henne: »Ingen rakkniv har kommit på mitt huvud, ty jag är en Guds nasir allt ifrån min moders liv.
Därför, om man rakar håret av mig, viker min styrka ifrån mig, så att jag bliver svag och är såsom alla andra människor.»
Då nu Delila insåg att han hade yppat för henne hela sin hemlighet, sände hon bud och kallade till sig filistéernas hövdingar; hon lät säga: »Kommen hitupp ännu en gång, ty han har nu yppat för mig hela sin hemlighet.»
Då kommo filistéernas hövdingar ditupp till henne och förde med sig penningarna.
Nu lagade hon så, att han somnade in på hennes knän; och sedan hon hade kallat till sig en man som på hennes befallning skar av de sju flätorna på hans huvud, begynte hon att få makt över honom, och hans styrka vek ifrån honom.
Därefter ropade hon: »Filistéerna äro över dig, Simson!»
När han då vaknade upp ur sömnen, tänkte han: »Jag gör mig väl fri, nu såsom de förra gångerna, och skakar mig lös»; ty han visste icke att HERREN hade vikit ifrån honom.
Men filistéerna grepo honom och stucko ut ögonen på honom.
Därefter förde de honom ned till Gasa och bundo honom med kopparfjättrar, och han måste mala i fängelset.
Men hans huvudhår begynte åter växa ut, sedan det hade blivit avrakat.
Och filistéernas hövdingar församlade sig för att anställa en stor offerfest åt sin gud Dagon och göra sig glada, ty de sade: »Vår gud har givit vår fiende Simson i vår hand.»
Och när folket såg honom, lovade de likaledes sin gud och sade: »Vår gud har givit vår fiende i vår hand honom som förödde vårt land och slog så många av oss ihjäl.»
Då nu deras hjärtan hade blivit glada, sade de: »Låt hämta Simson, för att han må förlusta oss.»
Och Simson blev hämtad ur fängelset och måste vara dem till förlustelse.
Och de hade ställt honom mellan pelarna.
Men Simson sade till den gosse som höll honom vid handen: »Släpp mig och låt mig komma intill pelarna som huset vilar på, så att jag får luta mig mot dem.»
Och huset var fullt med män och kvinnor, och filistéernas alla hövdingar voro där; och på taket voro vid pass tre tusen män och kvinnor, som sågo på, huru Simson förlustade dem.
Men Simson ropade till HERREN och sade: »Herre, HERRE, tänk på mig och styrk mig allenast denna gång, o Gud, så att jag får taga hämnd på filistéerna för ett av mina båda ögon.»
Därefter fattade Simson i de båda mittelpelare som huset vilade på, och tog fast tag mot dem; han fattade i den ena med högra handen och i den andra med vänstra.
Och Simson sade: »Må jag nu själv dö med filistéerna.»
Sedan böjde han sig framåt med sådan kraft, att huset föll omkull över hövdingarna och allt folket som fanns där.
Och de som han så dödade vid sin död voro flera än de som han hade dödat, medan han levde.
Och hans bröder och hela hans familj kommo ditned och togo honom upp med sig och begrovo honom mellan Sorga och Estaol, i hans fader Manoas grav.
Han hade då i tjugu år varit domare i Israel.
I Efraims bergsbygd levde en man som hette Mika.
Denne sade till sin moder: »De ett tusen ett hundra silversiklar som blevo dig fråntagna, och för vilkas skull du uttalade en förbannelse, som jag själv hörde, se, de penningarna finnas hos mig.
Det var jag som tog dem.»
Då sade hans moder: »Välsignad vare du, min son, av HERREN!»
Så gav han de ett tusen ett hundra silversiklarna tillbaka åt sin moder.
Men hans moder sade: »Härmed helgar jag dessa penningar åt HERREN och lämnar dem åt min son, för att han må låta göra en skuren och en gjuten gudabild.
Här lämnar jag dem nu tillbaka åt dig.»
Men han gav penningarna tillbaka åt sin moder.
Då tog hans moder två hundra siklar silver och gav dem åt en guldsmed, och denne gjorde därav en skuren och en gjuten gudabild, vilka sedan ställdes in i Mikas hus.
Mannen Mika hade så ett gudahus; han lät ock göra en efod och husgudar och insatte genom handfyllning en av sina söner till präst åt sig.
På den tiden fanns ingen konung i Israel; var och en gjorde vad honom behagade.
I Bet-Lehem i Juda levde då en ung man av Juda släkt; han var levit och bodde där såsom främling.
Denne man vandrade bort ifrån sin stad, Bet-Lehem i Juda, för att se om han funne någon annan ort där han kunde bo; och under sin färd kom han till Efraims bergsbygd, fram till Mikas hus.
Då frågade Mika honom: »Varifrån kommer du?»
Han svarade honom: »Jag är en levit från Bet-Lehem i Juda, och jag är nu stadd på vandring, för att se om jag finner någon annan ort där jag kan bo.»
Mika sade till honom: »Stanna kvar hos mig, och bliv fader och präst åt mig, så skall jag årligen giva dig tio siklar silver och vad kläder du behöver, och därtill din föda.»
Då följde leviten med honom.
Och leviten gick in på att stanna hos mannen, och denne behandlade den unge mannen såsom sin son.
Och Mika insatte leviten genom handfyllning, så att den unge mannen blev präst åt honom; och han var sedan kvar i Mikas hus.
Och Mika sade: »Nu vet jag att HERREN skall göra mig gott, eftersom jag har fått leviten till präst.»
På den tiden fanns ingen konung i Israel.
Och på den tiden sökte sig daniternas stam en arvedel till att bo i, ty ända dittills hade icke något område tillfallit den såsom arvedel bland Israels övriga stammar.
Så sände då Dans barn ur sin släkt fem män, uttagna bland dem, tappra män, från Sorga och Estaol, till att bespeja landet och undersöka det; och de sade till dem: »Gån åstad och undersöken landet.»
Så kommo de till Efraims bergsbygd, fram till Mikas hus; där stannade de över natten.
När de nu voro vid Mikas hus och kände igen den unge levitens sätt att tala, gingo de fram till honom och frågade honom: »Vem har fört dig hit?
Och vad gör du på detta ställe, och huru har du det här?»
Han omtalade då för dem: »Så och så gjorde Mika med mig; han gav mig lön, och jag blev präst åt honom.»
Då sade de till honom: »Fråga då Gud, så att vi få veta om den resa som vi äro stadda på skall bliva lyckosam.»
Prästen svarade dem: »Gån i frid.
Den resa som I ären stadda på står under HERRENS beskydd.»
Då gingo de fem männen vidare och kommo till Lais; och de sågo huru folket därinne bodde i trygghet, på sidoniernas sätt, stilla och trygga, och att ingen gjorde någon skada i landet genom att tillvälla sig makten; och de bodde långt ifrån sidonierna och hade intet att skaffa med andra människor.
När de sedan kommo åter till sina bröder i Sorga och Estaol, frågade deras bröder dem: »Vad haven I att säga?»
De svarade: »Upp, låt oss draga åstad mot dem!
Ty vi hava besett landet och funnit det mycket gott.
Skolen då I sitta stilla?
Nej, varen ej sena till att tåga åstad, så att I kommen dit och intagen landet.
När I kommen dit, kommen I till ett folk som känner sig tryggt, och landet har utrymme nog.
Ja, Gud har givit det i eder hand -- en ort där ingen brist är på något som jorden kan bära.»
Så bröto sex hundra man av daniternas släkt, omgjordade med vapen, upp därifrån, nämligen från Sorga och Estaol.
De drogo upp och lägrade sig vid Kirjat-Jearim i Juda.
Därför kallar man ännu i dag det stället för Dans läger; det ligger bakom Kirjat-Jearim.
Därifrån drogo de vidare till Efraims bergsbygd och kommo så fram till Mikas hus.
De fem män som hade varit åstad för att bespeja Lais' land togo då till orda och sade till sina bröder: »I mån veta att här i husen finnas en efod och husgudar och en skuren och en gjuten Gudabild.
Så betänken nu vad I bören göra.»
Då drogo de ditfram och kommo till den unge levitens hus, till Mikas hus, och hälsade honom.
Men de sex hundra männen av Dans barn ställde sig vid ingången till porten, omgjordade med sina vapen som de voro.
Och de fem män som hade varit åstad för att bespeja landet gingo upp och kommo ditin och togo den skurna gudabilden och efoden, så ock husgudarna och den gjutna gudabilden, under det att prästen stod vid ingången till porten jämte de sex hundra vapenomgjordade männen.
När nu de fem männen hade gått in i Mikas hus och tagit den skurna gudabilden med efoden och husgudarna och den gjutna gudabilden, sade prästen till dem: »Vad är det I gören!»
De svarade honom: »Tig, lägg handen på din mun, och gå med oss och bliv fader och präst åt oss.
Vilket är bäst för dig: att vara präst för en enskild mans hus eller att vara präst för en hel stam och släkt i Israel?»
Då blev prästens hjärta glatt, och han tog emot efoden och husgudarna och den skurna gudabilden och slöt sig till folket.
Sedan vände de sig åt annat håll och gingo vidare, och läto därvid kvinnor och barn och boskapen och det dyrbaraste godset föras främst i tåget.
Men när Dans barn hade kommit ett långt stycke väg från Mikas hus, upphunnos de av de män som voro bosatta i närheten av Mikas hus, och som under tiden hade samlat sig.
Vid dessas tillrop vände sig nu Dans barn om och frågade Mika: »Vad fattas dig, eftersom du kommer med en sådan hop?»
Han svarade: »I haven tagit de gudar som jag har gjort åt mig, därtill ock prästen, och så gån I eder väg.
Vad har jag nu mer kvar?
Och ändå frågen I mig: 'Vad fattas dig?'!»
Men Dans barn sade till honom: »Låt oss icke höra ett ord mer från dig.
Eljest kan det hända att några män i förbittring hugga ned eder, och då bliver du orsak till att I förloren livet, både du själv och ditt husfolk.»
Därefter fortsatte Dans barn sin väg; och när Mika såg att de voro starkare än han, vände han om och drog tillbaka hem igen.
Sedan de så hade tagit både vad Mika hade låtit förfärdiga och därtill hans präst, föllo de över folket i Lais, som levde stilla och i trygghet, och slogo dem med svärdsegg; men staden brände de upp i eld.
Och ingen kunde komma den till hjälp, ty den låg långt ifrån Sidon, och folket däri hade intet att skaffa med andra människor; den låg i Bet-Rehobs dal.
Sedan byggde de åter upp staden och bosatte sig där.
Och de gåvo staden namnet Dan efter sin fader Dan, som var son till Israel; förut hade staden hetat Lais.
Och Dans barn ställde där upp åt sig den skurna gudabilden; och Jonatan, son till Gersom, Manasses son, och hans söner voro präster åt daniternas stam, ända till dess att landets folk fördes bort i fångenskap.
De ställde upp åt sig den skurna gudabild som Mika hade gjort, och de hade denna kvar under hela den tid Guds hus var i Silo.
På den tiden, då ännu ingen konung fanns i Israel, bodde en levitisk man längst uppe i Efraims bergsbygd.
Denne tog till bihustru åt sig en kvinna från Bet-Lehem i Juda.
Men hans bihustru blev honom otrogen och gick ifrån honom till sin faders hus i Bet-Lehem i Juda; där uppehöll hon sig en tid av fyra månader.
Då stod hennes man upp och begav sig åstad efter henne, för att tala vänligt med henne och så föra henne tillbaka; och han hade med sig sin tjänare och ett par åsnor.
Hon förde honom då in i sin faders hus, och när kvinnans fader fick se honom, gick han glad emot honom.
Och hans svärfader, kvinnans fader, höll honom kvar, så att han stannade hos honom i tre dagar; de åto och drucko och voro där nätterna över.
När de nu på fjärde dagen stodo upp bittida om morgonen och han gjorde sig redo att resa, sade kvinnans fader till sin måg: »Vederkvick dig med ett stycke bröd; sedan mån I resa.»
Då satte de sig ned och åto båda tillsammans och drucko.
Därefter sade kvinnans fader till mannen: »Beslut dig för att stanna här över natten, och låt ditt hjärta vara glatt.»
Och när mannen ändå gjorde sig redo att resa, bad hans svärfader honom så enträget, att han ännu en gång stannade kvar där över natten.
På femte dagen stod han åter upp bittida om morgonen för att resa; då sade kvinnans fader: »Vederkvick dig först, och dröjen så till eftermiddagen.»
Därefter åto de båda tillsammans.
När sedan mannen gjorde sig redo att resa med sin bihustru och sin tjänare, sade hans svärfader, kvinnans fader, till honom: »Se, det lider mot aftonen; stannen kvar över natten, dagen nalkas ju sitt slut; ja, stanna kvar här över natten, och låt ditt hjärta vara glatt.
Sedan kunnen I i morgon bittida företaga eder färd, så att du får komma hem till din hydda.»
Men mannen ville icke stanna över natten, utan gjorde sig redo och reste sin väg, och kom så fram till platsen mitt emot Jebus, det är Jerusalem.
Och han hade med sig ett par sadlade åsnor; och hans bihustru följde honom.
Då de nu voro vid Jebus och dagen var långt framliden, sade tjänaren till sin herre: »Kom, låt oss taga in i denna jebuséstad och stanna där över natten.»
Men hans herre svarade honom: »Vi skola icke taga in i en främmande stad, där inga israeliter bo; låt oss draga vidare, fram till Gibea.»
Och han sade ytterligare till sin tjänare: »Kom, låt oss försöka hinna fram till en av orterna här och stanna över natten i Gibea eller Rama.»
Så drogo de vidare; och när de voro invid Gibea i Benjamin, gick solen ned.
Då togo de in där och kommo för att stanna över natten i Gibea.
Och när mannen kom ditin, satte han sig på den öppna platsen i staden, men ingen ville taga emot dem i sitt hus över natten.
Men då, om aftonen, kom en gammal man från sitt arbete på fältet, och denne man var från Efraims bergsbygd och bodde såsom främling i Gibea; ty folket där på orten voro benjaminiter.
När denne nu lyfte upp sina ögon, fick han se den vägfarande mannen på den öppna platsen i staden.
Då sade den gamle mannen: »Vart skall du resa, och varifrån kommer du?»
Han svarade honom: »Vi äro på genomresa från Bet-Lehem i Juda till den del av Efraims bergsbygd, som ligger längst uppe; därifrån är jag, och jag har gjort en resa till Bet-Lehem i Juda.
Nu är jag på väg till HERRENS hus, men ingen vill här taga emot mig i sitt hus.
Jag har både halm och foder åt våra åsnor, så ock bröd och vin åt mig själv och åt din tjänarinna och åt mannen som åtföljer oss, dina tjänare, så att intet fattas oss.»
Då sade den gamle mannen: »Frid vare med dig!
Men låt mig få sörja för allt som kan fattas dig.
Härute på den öppna platsen må du icke stanna över natten.»
Därefter förde han honom till sitt hus och fodrade åsnorna.
Och sedan de hade tvått sina fötter, åto de och drucko.
Under det att de så gjorde sina hjärtan glada, omringades plötsligt huset av männen i staden, onda män, som bultade på dörren; och de sade till den gamle mannen, som rådde om huset: »För hitut den man som har kommit till ditt hus, så att vi få känna honom.»
Då gick mannen som rådde om huset ut till dem och sade till dem: »Nej, mina bröder, gören icke så illa.
Eftersom nu denne man har kommit in i mitt hus, mån I icke göra en sådan galenskap.
Se, jag har en dotter som är jungfru, och han har själv en bihustru.
Dem vill jag föra hitut, så kunnen I kränka dem och göra med dem vad I finnen för gott.
Men med denne man mån I icke göra någon sådan galenskap.
Men männen ville icke höra på honom; då tog mannen sin bihustru och förde henne ut till dem.
Och de kände henne och hanterade henne skändligt hela natten ända till morgonen; först när morgonrodnaden gick upp, läto de henne gå.
Då kom kvinnan mot morgonen och föll ned vid ingången till mannens hus, där hennes herre var, och låg så, till dess det blev dager.
När nu hennes herre stod upp om morgonen och öppnade dörren till huset och gick ut för att fortsätta sin färd, fick han se sin bihustru ligga vid ingången till huset med händerna på tröskeln.
Han sade till henne: »Stå upp och låt oss gå.»
Men hon gav intet svar.
Då tog han och lade henne på åsnan; sedan gjorde mannen sig redo och reste hem till sitt.
Men när han hade kommit hem, fattade han en kniv och tog sin bi- hustru och styckade henne, efter benen i hennes kropp, i tolv stycken och sände styckena omkring över hela Israels land.
Och var och en som såg detta sade: »Något sådant har icke hänt eller blivit sett allt ifrån den dag då Israels barn drogo upp ur Egyptens land ända till denna dag.
Övervägen detta, rådslån och sägen edert ord.»
Då drogo alla Israels barn ut, och menigheten församlade sig såsom en man, från Dan ända till Beer-Seba, så ock från Gileads land, inför HERREN i Mispa.
Och de förnämsta i hela folket alla Israels stammar, trädde fram i Guds folks församling: fyra hundra tusen svärdbeväpnade mån till fots.
Men Benjamins barn fingo höra att de övriga israeliterna hade dragit upp till Mispa.
Och Israels barn sade: »Omtalen huru denna ogärning har tillgått.»
Då tog den levitiske mannen, den mördade kvinnans man, till orda och sade: »Jag och min bihustru kommo till Gibea i Benjamin för att stanna där över natten.
Då blev jag överfallen av Gibeas borgare; de omringade huset om natten för att våldföra sig på mig.
Mig tänkte de dräpa, och min bihustru kränkte de, så att hon dog.
Då tog jag min bihustru och styckade henne och sände styckena omkring över Israels arvedels hela område, eftersom de hade gjort en sådan skändlighet och galenskap i Israel.
Se, nu ären I allasammans här, I Israels barn.
Läggen nu fram förslag och råd här på stället.»
Då stod allt folket upp såsom en man och sade: »Ingen av oss må gå hem till sin hydda, ingen må begiva sig hem till sitt hus.
Detta är vad vi nu vilja göra med Gibea: vi skola låta lotten gå över det.
På vart hundratal i alla Israels stammar må vi taga ut tio män, och på vart tusental hundra, och på vart tiotusental tusen, för att dessa må skaffa munförråd åt folket, så att folket, när det kommer till Geba i Benjamin, kan göra med staden såsom tillbörligt är för all den galenskap som den har gjort i Israel.»
Så församlade sig vid staden alla män i Israel, endräktigt såsom en man.
Och Israels stammar sände åstad män till alla Benjamins stammar och läto säga; »Vad är det för en ogärning som har blivit begången ibland eder!
Lämnen nu ut de onda män som bo i Gibea, så att vi få döda dem och skaffa bort ifrån Israel vad ont är.»
Men benjaminiterna ville icke lyssna till sina bröders, de övriga israeliternas, ord.
I stället församlade sig Benjamins barn från sina städer till Gibea, för att draga ut till strid mot de övriga israeliterna.
På den dagen mönstrades Benjamins barn, de utgjorde från dessa städer tjugusex tusen svärdbeväpnade män; vid denna mönstring medräknades icke de som bodde i Gibea, vilka utgjorde sju hundra utvalda män.
Bland allt detta folk funnos sju hundra utvalda män som voro vänsterhänta; alla dessa kunde med slungstenen träffa på håret, utan att fela.
Och när Israels män -- Benjamin frånräknad -- mönstrades, utgjorde de fyra hundra tusen svärdbeväpnade män; alla dessa voro krigsmän.
Dessa bröto nu upp och drogo åstad till Betel och frågade Gud.
Israels barn sade: »Vem bland oss skall först draga ut i striden mot Benjamins barn?»
HERREN svarade: »Juda först.»
Då bröto Israels barn upp följande morgon och lägrade sig framför Gibea.
Därefter drogo Israels män ut till strid mot Benjamin; Israels män ställde upp sig till strid mot dem vid Gibea.
Men Benjamins barn drogo ut ur Gibea och nedgjorde på den dagen tjugutvå tusen man av Israel.
Folket, Israels män, tog dock åter mod till sig och ställde upp sig ännu en gång till strid på samma plats där de hade ställt upp sig första dagen.
Israels barn gingo nämligen upp och gräto inför HERRENS ansikte ända till aftonen; och de frågade HERREN: »Skall jag ännu en gång inlåta mig i strid med min broder Benjamins barn?»
Och HERREN svarade: »Dragen ut mot honom.»
När så Israels barn dagen därefter ryckte fram mot Benjamins barn,
drog ock Benjamin på andra dagen ut från Gibea mot Israels barn och nedgjorde av dem ytterligare aderton tusen man, allasammans svärdbeväpnade män.
Då drogo alla Israels barn upp, allt folket, och kommo till Betel och gräto och stannade där inför HERRENS ansikte och fastade på den dagen ända till aftonen; och de offrade brännoffer och tackoffer inför HERRENS ansikte.
Och Israels barn frågade HERREN (ty Guds förbundsark stod på den tiden där,
och Pinehas, son till Eleasar, Arons son, gjorde tjänst inför den på den tiden); de sade: »Skall jag ännu en gång draga ut till strid mot min broder Benjamins barn, eller skall jag avstå därifrån?»
HERREN svarade: »Dragen upp; ty i morgon skall jag giva honom i din hand.»
Då lade Israel manskap i bakhåll mot Gibea, runt omkring det.
Och därefter drogo Israels barn upp mot Benjamins barn, på tredje dagen, och ställde upp sig i slagordning mot Gibea likasom de förra gångerna.
Och Benjamins barn drogo ut mot folket och blevo lockade långt bort ifrån staden; och likasom det hade skett de förra gångerna, fingo de i början slå ihjäl några av folket på vägarna (både på den som går upp till Betel och på den som går till Gibea över fältet), kanhända ett trettiotal av Israels män.
Då tänkte Benjamins barn: »De äro slagna av oss, nu likasom förut.»
Men Israels barn hade träffat det avtalet: »Vi vilja fly och så locka dem långt bort ifrån staden, ut på vägarna.
Och alla Israels män hade brutit upp från platsen där de voro, och hade ställt upp sig i slagordning vid Baal-Tamar, under det att de israeliter som lågo i bakhåll bröto fram ifrån sin plats vid Maare-Geba.
Så kommo då tio tusen man, utvalda ur hela Israel, fram gent emot Gibea, och striden blev hård, utan att någon visste att olyckan var dem så nära.
Och HERREN lät Benjamin bliva slagen av Israel, och Israels barn nedgjorde av Benjamin på den dagen tjugufem tusen ett hundra man, allasammans svärdbeväpnade män.
Nu sågo Benjamins barn att de voro slagna.
Israels män gåvo nämligen plats åt Benjamin, ty de förlitade sig på bakhållet som de hade lagt mot Gibea.
Då skyndade sig de som lågo i bakhåll att falla in i Gibea; de som lågo i bakhåll drogo åstad och slogo alla invånarna i staden med svärdsegg.
Men de övriga israeliterna hade träffat det avtalet med dem som lågo i bakhåll, att dessa skulle låta en tjock rök såsom tecken stiga upp från staden.
Israels män vände alltså ryggen i striden.
Men sedan Benjamin i början hade fått slå ihjäl några av Israels man, kanhända ett trettiotal, och därvid hade tänkt: »Förvisso äro de slagna av oss, nu likasom i den förra striden»,
då kommo de att vända sig om, vid det att rökpelaren, det avtalade tecknet, begynte stiga upp från staden.
Och de fingo nu se hela staden förvandlad i lågor som slogo upp mot himmelen.
När då Israels män åter vände om, blevo Benjamins män förskräckta, ty nu sågo de att olyckan var dem nära.
Och de vände om för Israels män, bort åt öknen till, men fienderna hunno upp dem; och de som bodde i städerna där nedgjorde dem som hade kommit mitt emellan.
De omringade benjaminiterna, de satte efter dem och trampade ned dem på deras viloplats, ända fram emot Gibea, österut.
Så föllo av Benjamin aderton tusen man, allasammans tappert folk.
Då vände de övriga sig mot öknen och flydde dit, till Rimmons klippa; men de andra gjorde en efterskörd bland dem på vägarna, fem tusen man, och satte så efter dem ända till Gideom och slogo av dem två tusen man.
Alltså utgjorde de som på den dagen föllo av Benjamin tillsammans tjugufem tusen svärdbeväpnade män; alla dessa voro tappert folk.
Men av dem som vände sig mot öknen och flydde dit, till Rimmons klippa, hunno sex hundra man ditfram; dessa stannade på Rimmons klippa i fyra månader.
Emellertid vände Israels män tillbaka till Benjamins barn och slogo dem med svärdsegg, både dem av stadens befolkning, som ännu voro oskadda, och jämväl boskapen, korteligen, allt vad de träffade på; därtill satte de eld på alla städer som de träffade på.
Men Israels män hade svurit i Mispa och sagt: »Ingen av oss skall giva sin dotter till hustru åt någon benjaminit.»
Och nu kom folket till Betel och stannade där ända till aftonen inför Guds ansikte; och de brusto ut i bitter gråt
och sade: »Varför, o HERRE, Israels Gud, har sådant fått ske i Israel, att i dag en hel stam fattas i Israel?»
Dagen därefter stod folket bittida upp och byggde där ett altare och offrade brännoffer och tackoffer.
och Israels barn sade: »Finnes någon bland Israels alla stammar, som icke kom upp till HERREN med den övriga församlingen?»
Ty man hade svurit en dyr ed, att den som icke komme upp till HERREN i Mispa skulle straffas med döden.
Och Israels barn ömkade sig över sin broder Benjamin och sade: »Nu har en hel stam blivit borthuggen från Israel.
Vad skola vi göra för dem som äro kvar, så att de kunna få hustrur?
Ty själva hava vi ju svurit vid HERREN att icke åt dem giva hustrur av våra döttrar.»
Och då frågade åter: »Finnes bland Israels stammar någon som icke kom upp till HERREN i Mispa?»
Och se, från Jabes i Gilead hade ingen kommit till lägret, till församlingen där.
Ty när folket mönstrades, befanns det att ingen av invånarna i Jabes i Gilead var där.
Då sände menigheten dit tolv tusen av de tappraste männen och bjöd dessa och sade: »Gån åstad och slån invånarna i Jabes i Gilead med svärdsegg, också kvinnor och barn.
Ja, detta är vad I skolen göra: allt mankön och alla de kvinnor som hava haft med mankön att skaffa skolen I giva till spillo.
Men bland invånarna i Jabes i Gilead funno de fyra hundra unga kvinnor som voro jungfrur och icke hade haft med män, med mankön, att skaffa.
Dessa förde de då till lägret i Silo i Kanaans land.
Sedan sände hela menigheten åstad och underhandlade med de benjaminiter som befunno sig på Rimmons klippa, och tillbjöd dem fred.
Så vände nu Benjamin tillbaka; och man gav dem till hustrur de kvinnor från Jabes i Gilead, som man hade låtit leva.
Men dessa räckte ingalunda till för dem.
Och folket ömkade sig över Benjamin, eftersom HERREN hade gjort en rämna bland Israels stammar.
Och de äldste i menigheten sade: »Vad skola vi göra med dem som äro kvar, så att de kunna få hustrur?
Ty alla kvinnor äro ju utrotade ur Benjamin.»
Och de sade ytterligare: »De undkomna av Benjamin måste få en besittning, så att icke en stam bliver utplånad ur Israel.
Men själva kunna vi icke åt dem giva hustrur av våra döttrar, ty Israels barn hava svurit och sagt: Förbannad vare den som giver en hustru åt Benjamin.»
Och de sade vidare: »En HERREN högtid plägar ju hållas år efter år i Silo, som ligger norr om Betel, öster om den väg som går från Betel upp till Sikem, och söder om Lebona.»
Och de bjödo Benjamins barn och sade: »Gån åstad och läggen eder i försåt i vingårdarna.
När I då fån se Silos döttrar komma ut för att uppföra sina dansar, skolen I komma fram ur vingårdarna, och var och en av eder skall bland Silos döttrar rycka till sig en som kan bliva hans hustru; därefter skolen I begiva eder hem till Benjamins land.
Om sedan deras fäder eller deras bröder komma och beklaga sig för oss, vilja vi säga till dem: 'Förunnen oss dem; ty ingen av oss har tagit sig någon hustru i kriget.
I haven ju då icke själva givit dem åt dessa; ty i sådant fall haden I ådragit eder skuld.'»
Och Benjamins barn gjorde så och skaffade sig hustrur, lika många som de själva voro, bland de dansande kvinnor som de rövade.
Sedan begåvo de sig tillbaka till sin arvedel och byggde åter upp städerna och bosatte sig i dem.
Också de övriga israeliterna begåvo sig bort därifrån, var och en till sin stam och sin släkt, och drogo ut därifrån, var och en till sin arvedel.
På den tiden fanns ingen konung i Israel; var och en gjorde vad honom behagade.
På den tid då domarna regerade uppstod hungersnöd i landet.
Då drog en man från Bet-Lehem i Juda åstad med sin hustru och sina båda söner för att bosätta sig i Moabs land under någon tid.
Mannen hette Elimelek, hans hustru Noomi, och hans båda söner Mahelon och Kiljon; och de voro efratiter, från Bet-Lehem i Juda.
Så kommo de nu till Moabs land och vistades där.
Och Elimelek, Noomis man, dog; men hon levde kvar med sina båda söner.
Dessa skaffade sig moabitiska hustrur; den ena hette Orpa och den andra Rut.
Och sedan de hade bott där vid pass tio år, dogo också de båda, Mahelon och Kiljon; men kvinnan levde kvar efter sina båda söner och sin man.
Då stod hon upp med sina sonhustrur för att vända tillbaka från Moabs land; ty hon hade hört i Moabs land att HERREN hade sett till sitt folk och givit det bröd.
Så begav hon sig, jämte sina båda sonhustrur, från det ställe där hon hade vistats.
Men när de nu gingo sin väg fram, för att komma tillbaka till Juda land,
sade Noomi till sina båda sonhustrur: »Vänden om och gå hem igen, var och en till sin moder.
HERREN bevise godhet mot eder, såsom I haven gjort mot de båda döda och mot mig.
HERREN give eder att I mån finna ro, var i sin mans hus.»
Därefter kysste hon dem.
Men de brusto ut i gråt
och sade till henne: »Nej, vi vilja följa med dig tillbaka till ditt folk.»
Men Noomi svarade: »Vänden om, mina döttrar.
Varför skullen I gå med mig?
Kan väl jag ännu en gång få söner i mitt liv, vilka kunna bliva män åt eder?
Vänden om, mina döttrar, och gån hem, ty jag är nu för gammal att överlämna mig åt en man.
Och om jag än kunde tänka: 'Jag har ännu hopp', ja, om jag ock redan i natt överlämnade mig åt en man och så verkligen födde söner,
icke skullen I därför vänta, till dess att de hade blivit fullvuxna, icke skullen I därför stänga eder inne och förbliva utan män?
Bort det, mina döttrar!
Jag känner redan bedrövelse nog för eder skull, eftersom HERRENS hand så har drabbat mig.»
Då brusto de åter ut i gråt.
Och Orpa kysste sin svärmoder till avsked, men Rut höll sig alltjämt intill henne.
Då sade hon: »Se, din svägerska har vänt tillbaka till sitt folk och till sin gud; vänd ock du tillbaka och följ din svägerska.»
Men Rut svarade: »Sök icke intala mig att övergiva dig och vända tillbaka ifrån dig.
Ty dit du går vill ock jag gå, och där du stannar vill ock jag stanna.
Ditt folk är mitt folk, och din Gud är min Gud.
Där du dör vill ock jag dö, och där vill jag bliva begraven.
HERREN straffe mig nu och framgent, om något annat än döden kommer att skilja mig från dig.»
Då hon nu såg att denna stod fast i sitt beslut att gå med henne, upphörde hon att tala därom med henne.
Så gingo de båda med varandra, till dess att de kommo till Bet-Lehem.
Och när de kommo till Bet-Lehem, kom hela staden i rörelse för deras skull, och kvinnorna sade: »Detta är ju Noomi!»
Men hon sade till dem: »Kallen mig icke Noomi, utan kallen mig Mara, ty den Allsmäktige har låtit mycken bedrövelse komma över mig.
Rik drog jag härifrån, och tomhänt har HERREN låtit mig komma tillbaka.
Varför kallen I mig då Noomi, när HERREN har vittnat emot mig, när den Allsmäktige har låtit det gå mig så illa?»
Så kom då Noomi tillbaka med sin sonhustru, moabitiskan Rut, i det hon vände tillbaka från Moabs land.
Och de kommo till Bet-Lehem, när kornskörden begynte.
Men Noomi hade en frände på sin mans sida, en rik man av Elimeleks släkt, vid namn Boas.
Och moabitiskan Rut sade till Noomi: »Låt mig gå ut på åkern och plocka ax efter någon inför vilkens ögon jag finner nåd.»
Hon svarade henne: »Ja, gå, min dotter.»
Då gick hon åstad och kom till en åker och plockade där ax efter skördemännen; och det hände sig så för henne att åkerstycket tillhörde Boas, som var av Elimeleks släkt.
Och Boas kom just då dit från Bet-Lehem; och han sade till skördemännen: »HERREN vare med eder.»
De svarade honom: »HERREN välsigne dig.»
Och Boas frågade den bland tjänarna, som hade uppsikt över skördemännen: »Vem tillhör den unga kvinnan där?»
Tjänaren som hade uppsikt över skördemännen svarade och sade: »Det är en moabitisk kvinna, den kvinna som med Noomi har kommit hit från Moabs land.
Hon bad att hon skulle få plocka och hopsamla ax bland kärvarna, efter skördemännen; och så kom hon, och hon har hållit på allt sedan i morse ända till denna stund, utom att hon nyss har vilat något litet därinne.»
Då sade Boas till Rut: »Hör, min dotter: du skall icke gå bort och plocka ax på någon annan åker, ej heller gå härifrån, utan du skall hålla dig till mina tjänarinnor här.
Se efter, var skördemännen arbeta på åkern, och gå efter dem; jag har förbjudit mina tjänare att göra dig något för när.
Och om du bliver törstig, så gå till kärlen och drick av det som mina tjänare hämta.»
Då föll hon ned på sitt ansikte och bugade sig mot jorden och sade till honom: »Varför har jag funnit sådan nåd för dina ögon, att du tager dig an mig, fastän jag är en främling?»
Boas svarade och sade till henne: »För mig har blivit berättat allt vad du har gjort mot din svärmoder efter din mans död, huru du har övergivit din fader och din moder och ditt fädernesland, och vandrat åstad till ett folk som du förut icke kände.
HERREN vedergälle dig för vad du har gjort; ja, må full lön tillfalla dig från HERREN, Israels Gud, till vilken du har kommit, för att finna tillflykt under hans vingar.»
Hon sade: »Så må jag då finna nåd för dina ögon, min herre; ty du har tröstat mig och talat vänligt med din tjänarinna, fastän jag icke är såsom någon av dina tjänarinnor.»
Och när måltidsstunden var inne, sade Boas till henne: »Kom hitfram och ät av brödet och doppa ditt brödstycke i vinet.»
Då satte hon sig vid sidan av skördemännen; och han lade för henne rostade ax, och hon åt och blev mätt och fick därtill över.
Och när hon därefter stod upp för att plocka ax, bjöd Boas sina tjänare och sade: »Låten henne ock få plocka ax mellan kärvarna, och förfördelen henne icke.
Ja, I mån till och med draga ut strån ur knipporna åt henne och låta dem ligga, så att hon får plocka upp dem, och ingen må banna henne därför.»
Så plockade hon ax på åkern ända till aftonen; och när hon klappade ut det som hon hade plockat, var det vid pass en efa korn.
Och hon tog sin börda och gick in i staden, och hennes svärmoder fick se vad hon hade plockat.
Därefter tog hon fram och gav henne vad hon hade fått över, sedan hon hade ätit sig mätt.
Då sade hennes svärmoder till henne: »Var har du i dag plockat ax, och var har du arbetat?
Välsignad vare han som har tagit sig an dig!»
Då berättade hon för sin svärmoder hos vem hon hade arbetat; hon sade: »Den man som jag i dag har arbetat hos heter Boas.»
Då sade Noomi till sin sonhustru: »Välsignad vare han av HERREN, därför att han icke har undandragit sig att bevisa godhet både mot de levande och mot de döda!»
Och Noomi sade ytterligare till henne: »Den mannen är vår nära frände, en av våra bördemän.»
Moabitiskan Rut sade: »Han sade ock till mig: 'Håll dig till mina tjänare, ända till dess att de hava inbärgat hela min skörd.'»
Då sade Noomi till sin sonhustru Rut: »Ja, det är bäst, min dotter, att du går med hans tjänarinnor, så att man icke behandlar dig illa, såsom det kunde ske på en annan åker.»
Så höll hon sig då till Boas' tjänarinnor och plockade ax där, till dess både korn- och veteskörden voro avslutade.
Men hon bodde hos sin svärmoder.
Och hennes svärmoder Noomi sade till henne: »Min dotter, jag vill söka skaffa dig ro, för att det må gå dig väl.
Så hör då: Boas, med vilkens tjänarinnor du har varit tillsammans, är ju vår frände.
Och just i natt kastar han korn på sin tröskplats.
Så två dig nu och smörj dig och kläd dig, och gå ned till tröskplatsen.
Men laga så, att mannen icke får se dig, förrän han har ätit och druckit.
När han då lägger sig, så se efter, var han lägger sig, och gå dit och lyft upp täcket vid hans fötter och lägg dig där; han skall då själv säga dig vad du bör göra.»
Hon svarade: »Allt vad du säger vill jag göra.»
Och hon gick ned till tröskplatsen och gjorde alldeles såsom hennes svärmoder hade bjudit henne.
Ty när Boas hade ätit och druckit, så att hans hjärta blev glatt, och sedan han hade gått åstad och lagt sig invid sädeshögen, kom hon oförmärkt och lyfte upp täcket vid hans fötter och lade sig där.
Vid midnattstiden blev mannen uppskrämd och böjde sig framåt och fick då se en kvinna ligga vid hans fötter.
Och han sade: »Vem är du?»
Hon svarade: »Jag är Rut, din tjänarinna.
Bred ut din mantelflik över din tjänarinna, ty du är min bördeman.»
Då sade han: »Välsignad vare du av HERREN, min dotter!
Du har nu givit ett större bevis på din kärlek än förut, därigenom att du icke har lupit efter unga män, vare sig fattiga eller rika.
Så frukta nu icke, min dotter; allt vad du säger vill jag göra dig.
Ty allt folket i min stad vet att du är en rättskaffens kvinna.
Nu är det visserligen sant att jag är din bördeman; men en annan bördeman finnes, som är närmare än jag.
Stanna nu kvar i natt; om han i morgon vill taga dig efter bördesrätt, gott, må han då göra det, så sant HERREN lever.
Ligg nu kvar ända till morgonen.»
Så låg hon vid hans fötter ända till morgonen, men hon fick stå upp, innan ännu någon kunde känna igen den andre; ty han tänkte: »Det får icke bliva känt att kvinnan har kommit hit till tröskplatsen.»
Och han sade: »Räck hit manteln som du har på dig, och håll fram den.»
Och hon höll fram den.
Då mätte han upp sex mått korn och gav henne att bära; därefter gick hon in i staden.
Och när hon kom till sin svärmoder, sade denna: »Huru har det gått för dig, min dotter?»
Då berättade hon för henne allt vad mannen hade gjort mot henne;
och hon sade: »Dessa sex mått korn gav han mig, i det han sade: 'Du skall icke komma tomhänt hem till din svärmoder.'»
Då svarade hon: »Bida, min dotter, till dess du får se huru saken avlöper; ty mannen skall icke giva sig till ro, med mindre han i dag för saken till sitt slut.»
Och Boas hade gått upp till stadsporten och satt sig där.
Då hände sig att den bördeman som Boas hade talat om gick där fram; då nämnde han honom vid namn och sade: »Kom hit och sätt dig här.»
Och han kom och satte sig.
Därefter tog Boas till sig tio män av de äldste i staden och sade: »Sätten eder här.»
Och de satte sig.
Sedan sade han till bördemannen: »Det åkerstycke som tillhörde vår broder Elimelek har Noomi sålt, hon som kom tillbaka från Moabs land.
Därefter tänkte jag att jag skulle underrätta dig därom och säga: Köp det inför dem som här sitta och inför mitt folks äldste.
Om du vill taga det efter bördesrätt, så säg mig det, så att jag får veta det, ty ingen annan äger bördesrätt än du och, näst dig, jag själv.»
Han sade: »Jag vill taga det efter bördesrätt.»
Då sade Boas: »När du köper åkern av Noomis hand, då köper du den ock av moabitiskan Rut, den dödes hustru, med skyldighet att uppväcka den dödes namn och fästa det vid hans arvedel.»
Bördemannen svarade: »Då kan jag icke begagna mig av min bördesrätt, ty jag skulle därmed fördärva min egen arvedel.
Börda du åt dig vad jag skulle hava bördat, ty jag kan icke göra det.»
Men när någon bördade något eller avtalade ett byte, var det fordom sed i Israel att han, till stadfästelse av ett sådant avtal, drog av sig sin sko och gav den åt den andre; och detta gällde såsom ett vittnesbörd i Israel.
Så sade nu bördemannen till Boas: »Köp du det»; och han drog därvid av sig sin sko.
Då sade Boas till de äldste och till allt folket: »I ären i dag vittnen till att jag nu har köpt av Noomis hand allt vad som har tillhört Kiljon och Mahelon.
Därjämte har jag ock köpt moabitiskan Rut, Mahelons hustru, till hustru åt mig, för att uppväcka den dödes namn och fästa det vid hans arvedel, på det att den dödes namn icke må bliva utrotat bland hans bröder eller ur porten till hans stad.
I ären i dag vittnen härtill.»
Och allt folket i stadsporten, så ock de äldste, svarade: »Ja, och HERREN låte den kvinna som nu går in i ditt hus bliva lik Rakel och Lea, de båda som hava byggt upp Israels hus.
Och må du förkovra dig storligen i Efrata och göra dig ett namn i Bet-Lehem.
Och blive ditt hus såsom Peres' hus, hans som Tamar födde åt Juda, genom de avkomlingar som HERREN skall giva dig med denna unga kvinna.»
Så tog då Boas Rut till sig, och hon blev hans hustru, och han gick in till henne; och HERREN gav henne livsfrukt, och hon födde en son.
Då sade kvinnorna till Noomi: »Lovad vare HERREN, som i dag har så gjort, att det icke fattas dig en bördeman som skall få ett namn i Israel!
Han skall bliva dig en tröstare och en försörjare på din ålderdom; ty din sonhustru, som har dig kär, har fött honom, hon som är mer för dig än sju söner.»
Och Noomi tog barnet och lade det i sin famn och blev dess sköterska.
Och grannkvinnorna sade: »Noomi har fått en son»; och de gåvo honom namn, de kallade honom Obed.
Han blev fader till Isai, Davids fader.
Och detta är Peres' släktregister: Peres födde Hesron;
Hesron födde Ram; Ram födde Amminadab;
Amminadab födde Naheson; Naheson födde Salma;
Salmon födde Boas; Boas födde Obed;
Obed födde Isai, och Isai födde David.
I Ramataim-Sofim, i Efraims bergsbygd, levde en man som hette Elkana, son till Jeroham, son till Elihu, son till Tohu, son till Suf, en efraimit.
Han hade två hustrur; den ena hette Hanna, den andra Peninna.
Och Peninna hade barn, men Hanna var barnlös.
Den mannen begav sig år efter år upp från sin stad för att tillbedja och offra åt HERREN Sebaot i Silo, där Elis båda söner, Hofni och Pinehas, då voro HERRENS präster.
En dag offrade nu Elkana.
Och han plägade giva sin hustru Peninna och alla hennes söner och döttrar var sin andel av offret;
men åt Hanna gav han då en dubbelt så stor andel, ty han hade Hanna kär, fastän HERREN hade gjort henne ofruktsam.
Men hennes medtävlerska plägade, för att väcka hennes vrede, mycket retas med henne, därför att HERREN hade gjort henne ofruktsam.
För vart år, så ofta hon hade kommit upp till HERRENS hus, gjorde han på samma sätt, och den andra retades då med henne på samma sätt.
Och nu grät hon och åt intet.
Då sade hennes man Elkana till henne: »Hanna, varför gråter du?
Varför äter du icke?
Varför är du så sorgsen?
Är jag icke mer för dig än tio söner?
En gång när de hade ätit och druckit i Silo hände sig, medan prästen Eli satt på sin stol vid dörren till HERRENS tempel, att Hanna stod upp
och i sin djupa bedrövelse begynte bedja till HERREN under bitter gråt.
Och hon gjorde ett löfte och sade: HERRE Sebaot, om du vill se till din tjänarinnas lidande och tänka på mig och icke förgäta din tjänarinna, utan giva din tjänarinna en manlig avkomling, så vill jag giva denne åt HERREN för hela hans liv, och ingen rakkniv skall komma på hans huvud.»
När hon nu länge så bad inför HERREN och Eli därvid gav akt på hennes mun
-- Hanna talade nämligen i sitt hjärta; allenast hennes läppar rörde sig, men hennes röst hördes icke -- då trodde Eli att hon var drucken.
Därför sade Eli till henne: »Huru länge skall du bete dig såsom en drucken?
Laga så, att ruset går av dig.»
Men Hanna svarade och sade: »Nej, min herre, jag är en hårt prövad kvinna; vin och starka drycker har jag icke druckit, men jag utgöt nu min själ för HERREN.
Anse icke din tjänarinna för en ond kvinna, ty det är mitt myckna bekymmer och min myckna sorg som har drivit mig att tala ända till denna stund.»
Då svarade Eli och sade: »Gå i frid.
Israels Gud skall giva dig vad du har utbett dig av honom.»
Hon sade: »Låt din tjänarinna finna nåd för dina ögon.»
Så gick kvinnan sin väg och fick sig mat, och hon såg sedan icke mer så sorgsen ut.
Bittida följande morgon, sedan de hade tillbett inför HERREN, vände de tillbaka och kommo hem igen till Rama.
Och Elkana kände sin hustru Hanna, och HERREN tänkte på henne,
Och Hanna blev havande och födde en son, när tiden hade gått om; denne gav hon namnet Samuel, »ty», sade hon, »av HERREN har jag utbett mig honom.»
När sedan mannen Elkana med hela sitt hus begav sig upp för att offra åt HERREN sitt årliga slaktoffer och sitt löftesoffer,
gick Hanna icke med ditupp, utan sade till sin man: »Jag vill vänta, till dess att gossen har blivit avvand, då skall jag föra honom med mig, för att han må ställas fram inför HERRENS ansikte och sedan stanna där för alltid.»
Hennes man Elkana sade till henne: »Gör vad du finner för gott; stanna, till dess du har avvant honom; må HERREN allenast uppfylla sitt ord.»
Så stannade då hustrun hemma och gav sin son di, till dess hon skulle avvänja honom.
Men sedan hon hade avvant honom, tog hon honom med sig ditupp, jämte tre tjurar, en efa mjöl och en vinlägel; så förde hon honom in i HERRENS hus i Silo.
Men gossen var ännu helt ung.
Och de slaktade tjuren och förde så gossen fram till Eli.
Och hon sade: »Hör mig, min herre; så sant du lever, min herre, jag är den kvinna som stod här bredvid dig och bad till HERREN.
Om denne gosse bad jag; nu har HERREN givit mig vad jag utbad mig av honom.
Därför vill ock jag nu giva honom tillbaka åt HERREN; så länge han lever, skall han vara given åt HERREN.»
Och de tillbådo där HERREN.
Och Hanna bad och sade: »Mitt hjärta fröjdar sig i HERREN; mitt horn är upphöjt genom HERREN.
Min mun är vitt upplåten mot mina fiender; ty jag gläder mig över din frälsning.
Ingen är helig såsom HERREN ty ingen finnes förutom dig; ingen klippa är såsom vår Gud.
Fören icke beständigt så mycket högmodigt tal; vad fräckt är gånge icke ut ur eder mun.
Ty HERREN är en Gud som vet allt, och hos honom vägas gärningarna.
Hjältarnas bågar äro sönderbrutna, men de stapplande omgjorda sig med kraft.
De som voro mätta måste taga lega för bröd, men de som ledo hunger hungra icke mer.
Ja, den ofruktsamma föder sju barn, men den moder som fick många barn vissnar bort.
HERREN dödar och gör levande, han för ned i dödsriket och upp därifrån.
HERREN gör fattig, han gör ock rik; han ödmjukar, men han upphöjer ock.
Han upprättar den ringe ur stoftet, ur dyn lyfter han den fattige upp, ty han vill låta dem sitta bredvid furstar, och en härlig tron giver han dem till arvedel.
Ty jordens grundfästen äro HERRENS, och jordkretsen har han ställt på dem.
Sina frommas fötter bevarar han, men de ogudaktiga förgöras i mörkret, ty ingen förmår något genom egen kraft.
De som strida mot HERREN bliva krossade, ovan dem dundrar han i himmelen; ja, HERREN dömer jordens ändar.
Men han giver makt åt sin konung, han upphöjer sin smordes horn.
Och Elkana gick hem igen till Rama; gossen däremot gjorde tjänst inför HERREN under prästen Eli.
Men Elis söner voro onda män, de ville icke veta av HERREN.
På följande sätt plägade nämligen prästerna gå till väga med folket: så ofta någon offrade ett slaktoffer, kom prästens tjänare, medan köttet koktes, och hade en treuddig gaffel i sin hand;
den stack han ned i kitteln eller pannan eller krukan eller grytan, och allt vad han så fick upp med gaffeln, det tog prästen.
Så gjorde de mot alla israeliter som kommo dit till Silo.
Ja, till och med innan man hade förbränt det feta, kom prästens tjänare och sade till den som offrade: »Giv hit kött, så att jag kan steka det åt prästen, ty han vill icke hava kokt kött av dig, utan rått.»
Om då mannen svarade honom: »Först skall man nu förbränna det feta; tag sedan vad dig lyster», så sade han: »Nej, nu strax skall du lämna det, eljest tager jag det med våld.»
Och de unga männens synd var så mycket större inför HERREN som folket därigenom lärde sig att förakta HERRENS offer.
Men Samuel gjorde tjänst inför HERRENS ansikte, och var redan såsom gosse iklädd linne-efod.
Därtill plägade hans moder vart år göra åt honom en liten kåpa, som hon hade med sig till honom, när hon jämte sin man begav sig upp för att offra det årliga slaktoffret.
Då plägade Eli välsigna Elkana jämte hans hustru och säga: »HERREN skänke dig ytterligare avkomma med denna kvinna, i stället för den som hon utbad sig genom sin bön till HERREN.»
Och så gingo de hem igen.
Och HERREN såg till Hanna, och hon blev havande och födde tre söner och två döttrar.
Men gossen Samuel växte upp i HERRENS hus.
Då nu Eli, som var mycket gammal, fick höra allt vad hans söner gjorde mot hela Israel, och att de lågo hos de kvinnor som hade tjänstgöring vid ingången till uppenbarelsetältet,
sade han till dem: »Varför gören sådant, allt detta onda som jag hör allt folket här tala om eder?
Icke så, mina söner!
Det rykte jag hör vara gängse bland HERRENS folk är icke gott.
Om en människa försyndar sig mot en annan, så kan Gud medla för henne; men om en människa försyndar sig mot HERREN, vem kan då göra sig till medlare för henne?»
Men de lyssnade icke till sin faders ord, ty HERREN ville döda dem.
Gossen Samuel däremot växte till i ålder och välbehag både för HERREN och för människor.
Och en gudsman kom till Eli och sade till honom: »Så säger HERREN: Har jag icke uppenbarat mig för din faders hus, när de ännu voro i Egypten och tjänade Faraos hus?
Och har jag icke utvalt honom bland alla Israels stammar till präst åt mig, till att offra på mitt altare och antända rökelse och bära efod inför mitt ansikte?
Och gav jag icke åt din faders hus Israels barns alla eldsoffer?
Varför förtrampen I då de slaktoffer och spisoffer som jag har påbjudit i min boning?
Och huru kan du ära dina söner mer än mig, så att I göden eder med det bästa av var offergåva som mitt folk Israel bär fram?
Därför säger HERREN, Israels Gud: Väl har jag sagt att ditt och din faders hus skulle få göra tjänst inför mig evärdligen.
Men nu säger HERREN: Bort det!
Ty dem som ära mig vill jag ock ära, men de som förakta mig skola komma på skam.
Se, dagar skola komma, då jag skall avhugga din arm och din faders hus' arm, så att ingen skall bliva gammal i ditt hus.
Och du skall få se min boning lida nöd, trots allt det goda som vederfares Israel.
Och ingen skall någonsin bliva gammal i ditt eget hus.
Dock vill jag icke från mitt altare utrota var man av din slakt, så att jag kommer dina ögon att förtvina och din själ att försmäkta; men alla som växa upp i ditt hus skola dö, när de hava hunnit till manlig ålder.
Och tecknet härtill skall för dig vara det som skall övergå dina båda söner Hofni och Pinehas: på en och samma dag skola de båda dö.
Men jag skall låta en präst uppstå åt mig, som bliver beståndande, en som gör efter vad i mitt hjärta och min själ är; åt honom skall jag bygga ett hus som bliver beståndande, och han skall göra tjänst inför min smorde beständigt.
Och var och en som bliver kvar: av ditt hus skall komma och falla ned för honom, för att få en silverpenning eller en kaka bröd; han skall säga: 'Anställ mig vid någon prästsyssla, så att jag får en bit bröd att äta.'»
Så gjorde nu den unge Samuel tjänst inför HERREN under Eli.
Och HERRENS ord var sällsynt på den tiden, profetsyner voro icke vanliga.
Då nu en gång Eli, vilkens ögon hade begynt att bliva skumma, så att han icke kunde se, låg och sov på sin plats,
innan ännu Guds lampa hade slocknat, och medan också Samuel låg och sov, då hände sig i HERRENS tempel, där Guds ark stod,
att HERREN ropade på Samuel Denne svarade: »Här är jag.»
Därefter skyndade han till Eli och sade: »Här är jag; du ropade ju på mig.»
Men han svarade: »Jag har icke ropat; gå tillbaka och lägg dig.»
Och han gick och lade sig.
Men HERREN ropade ännu en gång på Samuel; och Samuel stod upp och gick till Eli och sade: »Här är jag; du ropade ju på mig.»
Men han svarade: »Jag har icke ropat, min son; gå tillbaka och lägg dig.»
Samuel hade nämligen ännu icke lärt att känna igen HERREN, och ännu hade icke något HERRENS ord blivit uppenbarat för honom.
Men HERREN ropade åter på Samuel, för tredje gången; och han stod upp och gick till Eli och sade: »Här är jag; du ropade ju på mig.
Då förstod Eli att det var HERREN som ropade på ynglingen.
Därför sade Eli till Samuel: »Gå och lägg dig; och om han vidare ropar på dig, så säg: 'Tala, HERRE; din tjänare hör.»
Och Samuel gick och lade sig på sin plats.
Då kom HERREN och ställde sig där och ropade såsom de förra gångerna: »Samuel!
Samuel!»
Samuel svarade: »Tala, din tjänare hör.»
Då sade HERREN till Samuel: »Se, jag skall i Israel göra något som kommer att genljuda i båda öronen på var och en som får höra det.
På den dagen skall jag låta komma över Eli allt vad jag har uttalat över hans hus, det första till det sista.
Ty jag har förkunnat för honom att jag skall vara domare över hans hus till evig tid, därför att han har syndat, i det han visste huru hans söner drogo förbannelse över sig och dock icke höll dem tillbaka.
Därför har jag ock med ed betygat om Elis hus: Sannerligen, Elis hus' missgärning skall icke någonsin kunna försonas, vare sig med slaktoffer eller med någon annat offergåva.»
Och Samuel låg kvar ända tills morgonen, då han öppnade dörrarna till HERRENS hus.
Och Samuel fruktade för att omtala synen for Eli.
Men Eli ropade på Samuel och sade: »Samuel, min son!
Denne svarade: »Här är jag.»
Han sade: »Vad var det han ta lade till dig?
Dölj det icke för mig.
Gud straffe dig nu och framgent, om du döljer for mig något enda ord av det han talade till dig.»
Då omtalade Samuel för honom alltsammans och dolde intet för honom.
Och han sade: »Han är HERREN; han göre vad honom täckes.
Men Samuel växte upp, och HERREN var med honom och lät intet av allt vad han hade talat falla till jorden.
Och hela Israel, från Dan ända till Beer-Seba, förstod att Samuel var betrodd att vara HERRENS profet.
Och HERREN fortfor att låta se sig i Silo; ty HERREN uppenbarade sig för Samuel i Silo genom HERRENS ord.
Och Samuels ord kom till hela Israel.
Och Israel drog ut till strid mot filistéerna och lägrade sig vid Eben-Haeser, under det filistéerna hade lägrat sig vid Afek.
Filistéerna ställde då upp sig i slagordning mot Israel, och striden utbredde sig, och israeliterna blevo slagna av filistéerna; dessa nedgjorde på slagfältet vid pass fyra tusen man.
När folket kom tillbaka till lägret sade de äldste i Israel: »Varför har HERREN i dag låtit oss bliva slagna av filistéerna?
Låt oss hämta hit till oss från Silo HERRENS förbundsark, för att den må komma och vara ibland oss och frälsa oss från våra fienders hand.»
Så sände då folket till Silo, och de buro därifrån HERREN Sebaots förbundsark, hans som tronar på keruberna; och Elis båda söner, Hofni och Pinehas, följde därvid med Guds förbundsark.
Då nu HERRENS förbundsark kom in i lägret, hov hela Israel upp ett stort jubelrop, så att det dånade i marken.
När då filistéerna hörde jubelropet, sade de: »Vad betyder detta stora jubelrop i hebréernas läger?»
Och de fingo veta att HERRENS ark hade kommit in i lägret.
Då blevo filistéerna förskräckta, ty de tänkte: »Gud har kommit in i lägret.»
Och de sade: »Ve oss!
Något sådant har förut icke hänt.
Ve oss!
Vem kan rädda oss från denne väldige Guds hand?
Det var denne Gud som slog egyptierna med alla slags plågor i öknen.
Men fatten dock mod och varen män, I filistéer, så att I icke bliven trälar åt hebréerna, såsom de hava varit trälar åt eder.
Ja, varen män och striden.»
Så stridde nu filistéerna, och israeliterna blevo slagna och flydde var och en till sin hydda, och nederlaget blev mycket stort: av Israel föllo trettio tusen man fotfolk.
Därtill blev Guds ark tagen, och Elis båda söner, Hofni och Pinehas, blevo dödade.
Och en benjaminit sprang från slagfältet och kom till Silo samma dag, med sönderrivna kläder och med jord på sitt huvud.
Och när han kom dit, satt Eli på sin stol vid sidan av vägen och såg utåt, ty hans hjärta bävade av oro för Guds ark.
Då nu mannen kom in i staden med budskapet, höjde hela staden upp klagorop.
Och när Eli hörde klagoropet, sade han: »Vad betyder detta larm?»
Då kom mannen skyndsamt dit och berättade det för Eli.
Men Eli var nittioåtta år gammal och hans ögon voro starrblinda, så att han icke kunde se.
Och mannen sade till Eli: »Jag är den som har kommit från slagfältet; jag har i dag flytt ifrån slagfältet.»
Då sade han: »Huru har det gått, min son?»
Budbäraren svarade och sade: »Israel har flytt för filistéerna, mycket folk har också stupat; dina båda söner, Hofni och Pinehas, äro ock döda, och därtill har Guds ark blivit tagen.»
När han nämnde om Guds ark, föll Eli baklänges av stolen vid sidan av porten och bröt nacken av sig och dog; ty mannen var gammal och tung.
Han hade då varit domare i Israel i fyrtio år.
Och när hans sonhustru, Pinehas' hustru, som var havande och nära att föda, fick höra ryktet om att Guds ark var tagen, och att hennes svärfader och hennes man voro döda, sjönk hon ned och födde sitt barn, ty födslovåndorna kommo över henne.
Och när hon då höll på att dö, sade kvinnorna som stodo omkring henne: »Frukta icke; du har fött en son.»
Men hon svarade intet och aktade icke därpå.
Och hon kallade gossen I-Kabod, och sade: »Härligheten är borta från Israel.»
Därmed syftade hon på att Guds ark var tagen, så ock på sin svärfader och sin man.
Hon sade: »Härligheten är borta från Israel», eftersom Guds ark var tagen.
När filistéerna hade tagit Guds ark, förde de den från Eben-Haeser till Asdod.
Där togo filistéerna Guds ark och förde in den i Dagons tempel och ställde den bredvid Dagon.
Men när asdoditerna bittida dagen därefter kommo dit, fingo de se Dagon ligga framstupa på jorden framför HERRENS ark.
Då togo de Dagon och satte honom upp igen på hans plats.
Men när de dagen därefter åter kommo dit bittida om morgonen, fingo de ånyo se Dagon ligga framstupa på jorden framför HERRENS ark; och Dagons huvud och hans båda händer lågo avslagna på tröskeln, allenast fiskdelen satt kvar på honom.
I Asdod trampar därför ännu i dag ingen på Dagons tröskel, varken någon av Dagons präster, ej heller någon annan som går in i Dagons tempel.
Och HERRENS hand var tung över asdoditerna; han anställde förödelse bland dem, i det han slog dem med bölder, såväl i Asdod som inom tillhörande områden.
Då nu invånarna i Asdod sågo att så skedde, sade de: »Israels Guds ark får icke stanna hos oss, ty hans hand vilar hårt på oss och på vår gud Dagon.»
Och de sände bud och läto församla till sig alla filistéernas hövdingar och sade: »Vad skola vi göra med Israels Guds ark?»
De svarade: »Israels Guds ark må flyttas till Gat.»
Då flyttade de Israels Guds ark dit.
Men sedan de hade flyttat den dit, kom genom HERRENS hand en mycket stor förvirring i staden; han slog invånarna i staden, både små och stora, så att bölder slogo upp på dem.
Då sände de Guds ark till Ekron.
Men när Guds ark kom till Ekron, ropade ekroniterna: »De hava flyttat Israels Guds ark till oss för att döda oss och vårt folk.»
Och de sände bud och läto för samla alla filistéernas hövdingar och sade: »Sänden bort Israels Guds ark, så att den får komma tillbaka till sin plats igen och icke dödar oss och vårt folk.»
Ty en dödlig förvirring hade uppstått i hela staden; Guds hand låg mycket tung på den.
De av invånarna som icke dogo blevo slagna med bölder; och ropet från staden steg upp mot himmelen.
Sedan nu HERRENS ark hade varit i filistéernas land i sju månader,
tillkallade filistéerna sina präster och spåmän och sade: »Vad skola vi göra med HERRENS ark?
Låten oss veta på vilket sätt vi skola sända den till dess plats igen.»
De svarade: »Om I viljen sända bort Israels Guds ark, skolen I icke sända bort den utan skänker; I måsten giva åt honom ett skuldoffer.
Då skolen I bliva botade, och det skall då också bliva eder kunnigt varför hans hand icke drager sig tillbaka från eder.»
Då frågade de: »Vad för ett skuldoffer skola vi giva åt honom?»
De svarade: »Fem bölder av guld och fem jordråttor av guld, lika många som filistéernas hövdingar; ty en och samma hemsökelse har träffat alla, också edra hövdingar.
I skolen göra avbildningar av edra bölder och avbildningar av jordråttorna som fördärva edert land; given så ära åt Israels Gud.
Kanhända tager han då bort sin tunga hand från eder, så ock från eder gud och från edert land.
Varför tillsluten I edra hjärtan, såsom egyptierna och Farao tillslöto sina hjärtan?
Måste icke dessa, sedan han hade utfört stora gärningar bland dem, släppa israeliterna, så att de fingo gå?
Så gören eder nu en ny vagn, och tagen två kor som giva di, och som icke hava burit något ok, och spännen korna för vagnen, men skiljen deras kalvar ifrån dem och låten dem stanna hemma.
Tagen så HERRENS ark och sätten den på vagnen, och läggen de gyllene klenoder I given honom såsom skuldoffer ned i ett skrin vid sidan av den, och låten den så gå åstad.
Sedan skolen I se efter: om den tager vägen till sitt land, upp mot Bet-Semes, så var det han som gjorde oss allt detta stora onda; men om så icke sker, då veta vi att det icke var hans hand som hemsökte oss.
Detta har då träffat oss allenast av en händelse.»
Männen gjorde så; de togo två kor som gåvo di och spände dem för vagnen; men deras kalvar behöllo de hemma.
Och de satte HERRENS ark på vagnen, därtill ock skrinet med jordråttorna av guld och med avbildningarna av svulsterna.
Och korna gingo raka vägen fram åt Bet-Semes till; de höllo alltjämt samma stråt och gingo där råmande, utan att vika av vare sig till höger eller till vänster.
Och filistéernas hövdingar gingo efter dem ända till Bet-Semes' område.
Men betsemesiterna höllo på med veteskörd i dalen.
När de nu lyfte upp sina ögon, fingo de se arken; och de blevo glada, då de sågo den.
Men när vagnen kom till betsemesiten Josuas åker, stannade den där; och där låg en stor sten.
Då höggo de sönder trävirket på vagnen och offrade korna till brännoffer åt HERREN.
Leviterna hade nämligen lyft ned HERRENS ark jämte skrinet som stod därbredvid, det vari de gyllene klenoderna funnos, och hade satt detta på den stora stenen.
Sedan offrade invånarna i Bet-Semes på den dagen brännoffer och slaktoffer åt HERREN.
Och när filistéernas fem hövdingar hade sett detta, vände de samma dag tillbaka till Ekron.
De svulster av guld som filistéerna gåvo såsom skuldoffer åt HERREN utgjorde: för Asdod en, för Gasa en, för Askelon en, för Gat en, för Ekron en.
Men jordråttorna av guld voro lika många som filistéernas alla städer under de fem hövdingarna, varvid medräknas både befästa städer och landsbygdens byar, intill den stora Sorgestenen, på vilken de satte ned HERRENS ark, och som finnes kvar ännu i dag, på betsemesiten Josuas åker.
Av invånarna i Bet-Semes blevo ock många slagna, därför att de hade sett på HERRENS ark; han slog sjuttio man bland folket, femtio tusen man.
Och folket sörjde däröver att HERREN hade slagit så många bland folket.
Och invånarna i Bet-Semes sade: »Vem kan bestå inför HERREN, denne helige Gud?
Och till vem skall han draga bort ifrån oss?»
Och de skickade sändebud till dem som bodde i Kirjat-Jearim och läto säga: »Filistéerna hava sänt tillbaka HERRENS ark; kommen hitned och hämten den upp till eder.
Då kommo Kirjat-Jearims män och hämtade HERRENS ark ditupp och förde den in i Abinadabs hus på höjden.
Och hans son Eleasar helgade de till att hava vården om HERRENS ark.
Och från den dag då arken fick sin plats i Kirjat-Jearim förflöt en lång tid: tjugu år förgingo; och hela Israels hus suckade nu efter HERREN.
Men Samuel sade till hela Israels hus: »Om I av allt edert hjärta viljen vända om till HERREN, så skaffen bort ifrån eder de främmande gudarna och Astarterna, och rikten edra hjärtan till HERREN och tjänen honom allena, så skall han rädda eder ifrån filistéernas hand.»
Då skaffade Israels barn bort Baalerna och Astarterna och tjänade HERREN allena.
Och Samuel sade: »Församlen hela Israel i Mispa, så vill jag där bedja till HERREN för eder.»
Då församlade de sig i Mispa och öste upp vatten och göto ut det in. för HERREN och fastade den dagen; och de sade där: »Vi hava syndat mot HERREN.»
Och Samuel dömde Israels barn i Mispa.
Men när filistéerna hörde att Israels barn hade församlat sig i Mispa, drogo filistéernas hövdingar ditupp mot Israel.
Då Israels barn hörde detta, blevo de förskräckta för filistéerna.
Och Israels barn sade till Samuel: »Hör icke upp att ropa för oss till HERREN, vår Gud, att han må frälsa oss ifrån filistéernas hand.»
Då tog Samuel ett dilamm och offrade det såsom ett heloffer, till brännoffer åt HERREN; och Samuel ropade till HERREN för Israel, och HERREN bönhörde honom.
Under det att Samuel offrade brännoffret, ryckte nämligen filistéerna fram till strid mot Israel; men HERREN lät ett starkt tordön dundra över filistéerna på den dagen och förvirrade dem, så att de blevo slagna av Israel.
Och Israels män drogo ut från Mispa och förföljde filistéerna och nedgjorde dem, under det att de förföljde dem ända till trakten nedanför Bet-Kar.
Då tog Samuel en sten och reste den mellan Mispa och Sen och gav den namnet Eben-Haeser, i det han sade: »Allt härintill har HERREN hjälpt oss.»
Så blevo filistéerna kuvade och kommo icke mer in i Israels land Och HERRENS hand var emot filistéerna, så länge Samuel levde.
Och de städer som filistéerna hade tagit från Israel kommo tillbaka till Israel, allasammans, från Ekron ända till Gat; och det tillhörande området tog Israel också igen ifrån filistéerna.
Och mellan Israel och amoréerna blev fred.
Och Samuel var domare i Israel, så länge han levde.
Vart år färdades han omkring till Betel, Gilgal och Mispa; och han dömde Israel på alla dessa platser.
Sedan plägade han vända tillbaka till Rama, ty där var hans hem, och där dömde han eljest Israel där byggde han ock ett altare åt HERREN.
Men när Samuel blev gammal, satte han sina söner till domare över Israel
Hans förstfödde son hette Joel, och hans andre son Abia; de hade sitt domarsäte i Beer-Seba.
Men hans söner vandrade icke på hans väg, utan veko av därifrån och sökte orätt vinning; de togo mutor och vrängde rätten.
Då församlade sig alla de äldste i Israel och kommo till Samuel i Rama.
Och de sade till honom: »Du är ju nu gammal, och dina söner vandra icke på dina vägar.
Så sätt nu en konung över oss till att döma oss, såsom alla andra folk hava.»
Men det misshagade Samuel, detta att de sade då: »Giv oss en konung, for att han må döma oss.»
Och Samuel bad till HERREN.
Då sade HERREN till Samuel »Lyssna till folkets ord, och gör allt vad de begära av dig; ty det är icke dig de hava förkastat, nej, mig hava de förkastat, i det de icke vilja att jag skall vara konung över dem.
Såsom de alltid hava gjort, från den dag då jag förde dem upp ur Egypten ända till denna dag, i det att de hava övergivit mig och tjänat andra gudar, så göra de nu ock mot dig.
Så lyssna nu till deras ord.
Dock må du högtidligt varna dem och förkunna för dem den konungs rätt, som kommer att regera över dem.»
Och Samuel sade till folket, som hade begärt en konung av honom, allt vad HERREN hade talat.
Han sade: »Detta bliver den konungs rätt, som kommer att regera över eder: Edra söner skall han taga och skall sätta dem på sina vagnar och hästar, till sin tjänst, eller ock skola de nödgas löpa framför hans vagnar.
Andra av dem skall han taga och sätta till sina över- och underhövitsmän, och andra skola nödgas plöja hans åkerjord och inbärga hans skörd och förfärdiga hans krigsredskap och hans vagnsredskap.
Edra döttrar skall han taga till salvoberederskor, kokerskor och bagerskor.
Edra bästa åkrar, vingårdar och olivplanteringar skall han taga och skall giva dem åt sina tjänare;
och han skall taga tionde av edra sädesfält och edra vingårdar och giva åt sina hovmän och tjänare.
Därtill skall han taga edra tjänare och edra tjänarinnor och edra bästa ynglingar, så ock edra åsnor, och bruka dem för sitt behov.
Av eder småboskap skall han taga tionde, och I skolen vara hans trälar.
När I då ropen om hjälp för dem konungs skull som I själva haven utvalt åt eder, då skall HERREN icke svara eder.
Men folket ville icke lyssna till Samuels ord, utan sade: »Nej, en konung måste vi hava över oss.»
Vi vilja bliva lika alla andra folk; vi vilja hava en konung som dömer oss, och som drager ut i spetsen för oss till att föra våra krig.»
Då nu Samuel hörde allt detta som folket sade, framförde han det till HERREN.
Men HERREN sade till Samuel: »Lyssna till deras ord, och sätt en konung över dem.»
Då sade Samuel till Israels män: »Gån hem, var och en till sin stad.»
I Benjamin levde en man som hette Kis, son till Abiel, son till Seror, son till Bekorat, son till Afia, son till en benjaminit; och han var en rik man.
Han hade en son som hette Saul, en ståtlig och fager man; bland Israels barn fanns ingen man som var fagrare än han; han var huvudet högre än allt folket.
Nu hade Kis', Sauls faders, åsninnor kommit bort för honom; därför sade Kis till sin son Saul: »Tag med dig en av tjänarna och stå upp och gå åstad och sök efter åsninnorna.»
Då gick han genom Efraims bergsbygd och därefter genom Salisalandet; men de funno dem icke.
Så gingo de genom Saalimslandet, men där voro de icke; sedan gick han genom Benjamins land, men de funno dem icke heller där.
När de så hade kommit in i Sufs land, sade Saul till tjänaren som han hade med sig: »Kom, låt oss gå hem igen; min fader kunde eljest, stället för att tänka på åsninnorna, bliva orolig för vår skull.»
Men han svarade honom: »Se, i denna stad finnes en gudsman; han är en ansedd man; allt vad han säger, det sker.
Låt oss nu gå dit; måhända kan han säga oss något om den färd vi hava företagit oss.»
Då sade Saul till sin tjänare: »Men om vi gå dit, vad skola vi då taga med oss åt mannen?
Brödet är ju slut i våra ränslar, och vi hava icke heller någon annan gåva att taga med oss åt gudsmannen.
Eller vad hava vi väl?»
Tjänaren svarade Saul ännu en gång och sade: »Se, här har jag i min ägo en fjärdedels sikel silver; den vill jag giva åt gudsmannen, för att han må säga oss vilken väg vi böra gå.»
(Fordom sade man så i Israel, när man gick för att fråga Gud: »Kom, låt oss gå till siaren.»
Ty den som man nu kallar profet kallade man fordom siare.)
Saul sade till sin tjänare: »Ditt förslag är gott; kom, låt oss gå.»
Så gingo de till staden där gudsmannen fanns.
När de nu gingo uppför höjden där staden låg, träffade de några flickor som hade gått ut för att hämta vatten; dem frågade de: »Är siaren här?»
De svarade dem och sade: »Ja, helt nära.
Skynda dig nu, ty han har i dag kommit till staden; folket firar nämligen i dag en offerfest på offerhöjden.
Om I nu gån in i staden, träffen I honom, innan han går upp på höjden till måltiden, ty folket äter icke, förrän han kommer.
Han skall välsigna offret; först sedan begynna de inbjudna att äta.
Gån därför nu ditupp, ty just nu kunnen I träffa honom.»
Så gingo de upp till staden.
Och just när de kommo in i staden, mötte de Samuel, som var stadd på väg upp till offerhöjden.
Men dagen innan Saul kom hade HERREN uppenbarat för Samuel och sagt:
»I morgon vid denna tid skall jag sända till dig en man från Benjamins land, och honom skall du smörja till furste över mitt folk Israel; han skall frälsa mitt folk ifrån filistéernas hand.
Ty jag har sett till mitt folk, eftersom deras rop har kommit till mig.»
När nu Samuel fick se Saul, gav HERREN honom den uppenbarelsen: »Se där är den man om vilken jag sade till dig: Denne skall styra mitt folk.»
Men Saul gick fram till Samuel i porten och sade: »Säg mig var siaren bor.»
Samuel svarade Saul och sade: »Jag är siaren.
Gå före mig upp på offerhöjden, ty I skolen äta där med mig i dag.
Men i morgon vill jag låta dig gå; och om allt vad du har på hjärtat vill jag giva dig besked.
Och vad angår åsninnorna, som nu i tre dagar hava varit borta för dig, skall du icke bekymra dig för dem, ty de äro återfunna.
Vem tillhör för övrigt allt vad härligt är i Israel, om icke dig och hela din faders hus?»
Saul svarade och sade: »Jag är ju en benjaminit, från en av de minsta stammarna i Israel, och min släkt är ju den ringaste bland alla släkter i Benjamins stammar.
Varför talar du då till mig på det sättet?»
Men Samuel tog Saul och hans tjänare och förde dem upp i salen och gav dem plats överst bland de inbjudna, vilka voro vid pass trettio män.
Och Samuel sade till kocken: »Giv hit det stycke som jag gav dig, och som jag sade att du skulle förvara hos dig.»
Då tog kocken fram lårstycket med vad därtill hörde, och satte det fram för Saul; och Samuel sade: »Se, här sättes nu fram för dig det som har blivit sparat; ät därav.
Ty just för denna stund blev det undanlagt åt dig, då när jag sade att jag hade inbjudit folket.»
Så åt Saul den dagen med Samuel.
Därefter gingo de ned från offerhöjden och in i staden.
Sedan samtalade han med Saul uppe på taket.
Men bittida följande dag, när morgonrodnaden gick upp, ropade Samuel uppåt taket till Saul och sade: »Stå upp, så vill jag ledsaga dig till vägs.»
Då stod Saul upp, och de gingo båda åstad, han och Samuel.
När de så voro på väg ned mot ändan av staden, sade Samuel till Saul: »Säg till tjänaren att han skall gå före oss» -- och han fick gå -- »men du själv må nu stanna här, så vill jag låta dig höra vad Gud har talat.»
Och Samuel tog sin oljeflaska och göt olja på hans huvud och kysste honom och sade: »Se, HERREN har smort dig till furste över sin arvedel.
När du nu går ifrån mig, skall du invid Rakels grav, vid Benjamins gräns, vid Selsa, träffa två män; dessa skola säga till dig: 'Åsninnorna som du gick åstad att söka äro återfunna; din fader tänker därför icke mer på åsninnorna, men han är orolig för eder skull och säger: Vad skall jag göra för att finna min son?'
Och när du har gått därifrån ett stycke fram och kommit till Tabors terebint skall du där möta tre män som äro på väg upp till Gud i Betel.
En bär tre killingar, en bar tre brödkakor, och en bär en vinlägel.
Dessa skola hälsa dig och giv dig två bröd, och du skall taga emot vad de giva.
Sedan kommer du till Guds Gibea, där filistéernas fogdar äro.
Och när du kommer dit in i staden, skall du träffa på en skara profeter, som komma ned från offerhöjden där, med psaltare, puka, flöjt och harpa före sig, under det att de själva äro i profetisk hänryckning.
Och HERRENS Ande skall komma över dig, så att också du fattas av hänryckning likasom de; och du skall då bliva förvandlad till en annan människa.
När du nu ser att dessa tecken inträffa, då må du göra vad tillfället giver vid handen, ty Gud är med dig.
Sedan må du gå ned före mig till Gilgal, så skall jag komma ditned till dig, för att offra brännoffer och tackoffer; sju dagar skall du vänta till dess jag kommer till dig och förkunnar för dig vad du skall göra.
I det han nu vände sig om för att gå ifrån Samuel, förvandlade Gud hans sinne och gav honom ett annat hjärta; och alla dessa tecken inträffade samma dag.
När de kommo till Gibea, mötte honom där en skara profeter; då kom Guds Ande över honom, så att han, mitt ibland dem, själv fattades av profetisk hänryckning.
Då nu alla som förut kände honom fingo se honom vara i hänryckning likasom profeterna, sade folket sinsemellan: »Vad har skett med Kis' son?
Är ock Saul bland profeterna?»
Men en av männen därifrån svarade och sade: »Vem är då dessas fader?» -- Härav uppkom ordspråket: »Är ock Saul bland profeterna?»
Men när hans profetiska hänryckning hade upphört, gick han upp på offerhöjden.
Då frågade Sauls farbroder honom och hans tjänare: »Var haven I varit?»
Han svarade: »Borta för att söka åsninnorna.
Men när vi sågo att de ingenstädes voro att finna, gingo vi till Samuel.»
Då sade Sauls farbroder: »Tala om for mig vad Samuel sade till eder.»
Saul svarade sin farbroder: »Han omtalade för oss att åsninnorna voro återfunna.»
Men vad Samuel hade sagt om konungadömet omtalade han icke för honom.
Därefter kallade Samuel folket tillsammans till HERREN, i Mispa.
Och han sade till Israels barn: »Så säger HERREN, Israels Gud: Jag har fört Israel upp ur Egypten, och jag räddade eder icke allenast undan Egypten, utan ock undan alla andra konungadömen som förtryckte eder.
Men nu haven I förkastat eder Gud, som själv frälste eder ur alla edra olyckor och trångmål, och haven sagt till honom: 'Sätt en konung över oss.'
Så träden nu fram inför HERREN efter edra stammar och edra ätter.»
Därpå lät Samuel alla Israels stammar gå fram; då träffades Benjamin stam av lotten.
När han sedan lät Benjamins stam gå fram efter dess släkter, träffade Matris släkt av lotten; därpå träffades Saul, Kis' son, av lotten, men när de då sökte efter honom, stod han icke att finna.
Då frågade de HERREN ännu en gång: »Har någon mer kommit hit?
HERREN svarade: »Han har gömt sig bland trossen.»
Då skyndade de dit och hämtad honom därifrån, och när han nu trädde fram bland folket, var han huvudet högre än allt folket.
Och Samuel sade till allt folket: »Här sen I nu den som HERREN har utvalt; ingen är honom lik bland allt folket.»
Då jublade allt folket och ropade: »Leve konungen!»
Och Samuel kungjorde för folket konungadömets rätt och tecknade upp den i en bok och lade ned den inför HERREN.
Sedan lät Samuel allt folket gå hem, var och en till sitt.
Också Saul gick hem till Gibea; och honom följde en härskara av män vilkas hjärtan Gud hade rört.
Men några onda män sade: »Vad hjälp skulle denne kunna giva oss?»
Och de föraktade honom och buro icke fram skänker till honom.
Men han låtsade som om han icke märkte det.
Och ammoniten Nahas drog upp och belägrade Jabes i Gilead.
Då sade alla män i Jabes till Nahas: »Slut fördrag med oss, så vilja vi bliva dig underdåniga.»
Men ammoniten Nahas svarade dem: »På det villkoret vill jag sluta fördrag med eder, att jag får sticka ut högra ögat på eder alla och därmed tillfoga hela Israel smälek.»
De äldste i Jabes sade till honom: »Giv oss sju dagars uppskov, så att vi kunna skicka sändebud över hela Israels land; om då ingen vill hjälpa oss, så skola vi giva oss åt dig.»
Så kommo nu sändebuden till Sauls Gibea och omtalade detta för folket.
Då brast allt folket ut i gråt.
Men just då kom Saul gående bakom sina oxar från åkern.
Och Saul frågade: »Vad fattas folket, eftersom de gråta?»
Och de förtäljde för honom vad mannen från Jabes hade sagt.
Då kom Guds Ande över Saul, när han hörde detta, och hans vrede upptändes högeligen.
Och han tog ett par oxar och styckade dem och sände styckena omkring över hela Israels land med sändebuden och lät säga: »Den som icke drager ut efter Saul och Samuel, med hans oxar skall så göras.»
Då föll en förskräckelse ifrån HERREN över folket, så att de drogo ut såsom en man.
Och han mönstrade dem i Besek, och Israels barn utgjorde då tre hundra tusen, och Juda män trettio tusen.
Och de sade till sändebuden som hade kommit: »Så skolen I säga till männen i Jabes i Gilead: I morgon skolen I få hjälp, när solen bränner som hetast.»
Och sändebuden kommo och förkunnade detta för männen i Jabes; och dessa blevo glada däröver.
Nu läto männen i Jabes säga: »I morgon vilja vi giva oss åt eder, och I mån då göra med oss vadhelst I finnen för gott.»
Dagen därefter fördelade Saul folket i tre hopar; och de trängde in i lägret vid morgonväkten och nedgjorde ammoniterna, och upphörde först när det var som hetast på dagen.
Och de som kommo undan blevo så kringspridda, att icke två av dem kommo undan tillsammans.
Då sade folket till Samuel: »Vilka voro de som sade: 'Skulle Saul bliva konung över oss!'
Given hit dessa män, så att vi få döda dem.»
Men Saul sade: »På denna dag skall ingen dödas, ty i dag har HERREN givit seger åt Israel.»
Och Samuel sade till folket: »Kom, låt oss gå till Gilgal och där förnya konungadömet.»
Då gick allt folket till Gilgal och gjorde Saul till konung där, inför HERRENS ansikte, i Gilgal; och de offrade där tackoffer inför HERRENS ansikte.
Och Saul och alla Israels män voro där uppfyllda av glädje.
Och Samuel sade till hela Israel: »Se, jag har lyssnat till edra ord och gjort allt vad I haven begärt av mig; jag har satt en konung över eder.
Nu är det eder konung som skall vara eder ledare, nu då jag är gammal och grå; I haven ju redan mina söner ibland eder.
Hittills är det jag som har varit eder ledare, från min ungdom ända till denna dag.
Se har står jag, vittnen nu mot mig inför HERREN och inför hans smorde.
Har jag tagit någons oxe, eller har jag tagit någons åsna?
Har jag förtryckt någon eller övat våld mot någon?
Har jag tagit mutor av någon, för att jag skulle se genom fingrarna med honom?
Jag vill då giva eder ersättning därför.»
De svarade: »Du har icke förtryckt oss, du har icke övat våld mot oss; och från ingen människa har du tagit något.»
Då sade han till dem: »HERREN vare vittne mot -- eder, och hans smorde vare ock vittne denna dag, att I icke haven funnit något i min hand.»
De svarade: »Ja, vare det så.»
Samuel sade till folket: »Ja, HERREN vare vittne, han som lät Mose och Aron uppstå och förde edra fäder upp ur Egyptens land.
Så träden nu fram, för att jag må gå till rätta med eder inför HERREN angående allt gott som HERREN i sin rättfärdighet har gjort mot eder och mot edra fäder.
När Jakob hade kommit fram till Egypten, ropade edra fäder till HERREN, och HERREN sände Mose och Aron, som förde edra fäder ut ur Egypten och läto dem bosätta sig här i landet.
Men när de glömde HERREN, sin Gud, sålde han dem i Siseras hand, härhövitsmannens i Hasor, och i filistéernas hand och i Moabs konungs hand, och dessa stridde mot dem.
Men då ropade till HERREN och sade: 'Vi hava syndat, ty vi hava övergivit HERREN och tjänat Baalerna och Astarterna; men rädda oss nu från våra fienders hand, så vilja vi tjäna dig.'
Då sände HERREN Jerubbaal och Bedan och Jefta och Samuel och räddade eder från edra fienders hand runt omkring, så att I fingen bo i trygghet.
Men när I sågen att Nahas, Ammons barns konung, kom emot eder, saden I till mig: 'Nej, en konung måste regera över oss', fastän det är HERREN, eder Gud, som är eder konung.
Och se, här är nu den konung I haven utvalt, den som I haven begärt; se, HERREN har satt en konung över eder.
Allenast man I nu frukta HERREN och tjäna honom och höra hans röst och icke vara gensträviga mot HERRENS befallning.
Ja, både I och den konung som regerar över eder mån följa HERREN, eder Gud.
Men om I icke hören HERRENS röst, utan ären gensträviga mot HERRENS befallning, då skall HERRENS hand drabba eder likasom edra fäder.
Träden nu ock fram och sen det stora under som HERREN skall göra inför edra ögon.
Nu är ju tiden för veteskörden; men jag vill ropa till HERREN att han må låta det dundra och regna.
Så skolen I märka och se huru mycket ont I haven gjort i HERRENS ögon genom eder begäran att få en konung.»
Och Samuel ropade till HERREN, och HERREN lät det dundra och regna på den dagen.
Då betogs allt folket av stor fruktan för HERREN och för Samuel.
Och allt folket sade till Samuel: »Bed för dina tjänare till HERREN, din Gud, att vi icke må dö, eftersom vi till alla våra andra synder ock hava lagt det onda att vi hava begärt att få en konung.»
Samuel sade till folket: »Frukten icke.
Väl haven I gjort allt detta onda; men viken nu blott icke av ifrån HERREN, utan tjänen HERREN av allt edert hjärta.
Viken icke av; ty då följen I tomma avgudar, som varken kunna hjälpa eller rädda, eftersom de äro allenast tomhet.
Ty HERREN skall icke förskjuta sitt folk, för sitt stora namns skull, eftersom HERREN har behagat att göra eder till sitt folk.
Vare det ock fjärran ifrån mig att jag skulle så synda mot HERREN, att jag upphörde att bedja för eder!
Jag vill fastmer lära eder den goda och rätta vägen.
Allenast frukten HERREN och tjänen honom troget av allt edert hjärta.
Ty sen vilka stora ting han har gjort med eder!
Men om I gören vad ont är, så skolen både I och eder konung förgås.»
Saul hade varit konung ett år, och när han nu regerade över Israel på andra året,
utvalde han åt sig tre tusen män ur Israel.
Av dessa hade Saul själv hos sig två tusen i Mikmas och i Betels bergsbygd, och ett tusen hade Jonatan hos sig i Gibea i Benjamin.
Men det övriga folket hade han låtit gå hem, var och en till sin hydda.
Och Jonatan dräpte filistéernas fogde i Geba; och filistéerna fingo höra det.
Men Saul lät stöta i basun över hela landet och säga: »Detta må hebréerna höra.»
Så fick hela Israel höra omtalas att Saul hade dräpt filistéernas fogde, och att Israel därigenom hade blivit förhatligt för filistéerna.
Och folket bådades upp att följa Saul till Gilgal.
Under tiden hade filistéerna församlat sig för att strida mot Israel: trettio tusen vagnar och sex tusen ryttare, och fotfolk så talrikt som sanden på havets strand; och de drogo upp och lägrade sig vid Mikmas, öster om Bet-Aven.
Då nu israeliterna sågo sig vara i nöd, i det att folket svårt ansattes, gömde sig folket i grottor, i skogssnår och bland klippor, i fasta valv och i gropar.
Och somliga av hebréerna gingo över Jordan in i Gads och Gileads land.
Men Saul var ännu kvar i Gilgal; och allt folket följde honom med bävan.
När han nu hade väntat sju dagar, intill den tid Samuel hade bestämt men Samuel likväl icke kom till Gilgal, begynte folket skingra sig och gå ifrån honom.
Då sade Saul: »Fören fram till mig brännoffers- och tackoffersdjuren.»
Därpå frambar han brännoffret.
Men just när han hade slutat att frambära brännoffret, kom Samuel.
Då gick Saul honom till mötes för att hälsa honom.
Men Samuel sade: »Vad har du gjort!»
Saul svarade: »När jag såg att folket skingrade sig och gick ifrån mig, under det att du icke kom inom den bestämda tiden, fastän filistéerna voro församlade vid Mikmas,
då tänkte jag: Nu komma filistéerna hitned mot mig i Gilgal, och jag har ännu icke bönfallit inför HERREN.
Då tog jag mod till mig och offrade brännoffret.»
Samuel sade till Saul: »Du har handlat dåraktigt.
Du har icke hållit det bud HERREN, din Gud, har givit dig; eljest skulle HERREN hava befäst ditt konungadöme över Israel för evig tid.
Men nu skall ditt konungadöme icke bliva beståndande.
HERREN har sökt sig en man efter sitt hjärta, och honom har HERREN förordnat till furste över sitt folk, eftersom du icke har hållit vad HERREN bjöd dig.»
Därefter stod Samuel upp och gick från Gilgal till Gibea i Benjamin.
Men Saul mönstrade det folk som fanns hos honom: vid pass sex hundra man.
Och Saul och hans son Jonatan stannade i Geba i Benjamin med det folk som fanns hos dem, under det att filistéerna hade lägrat sig vid Mikmas.
Och en härskara, delad i tre hopar, drog ut ur filistéernas läger för att härja: en hop tog vägen till Ofra i Sualslandet,
en hop tog vägen till Bet-Horon, och en hop tog vägen till det område som vetter åt Seboimsdalen, åt öknen till.
Ingen smed fanns då i hela Israels land, ty filistéerna fruktade att hebréerna skulle låta göra sig svärd eller spjut.
Och så måste en israelit alltid begiva sig ned till filistéerna, om han ville låta vässa sin lie eller sin plogbill eller sin yxa eller sin skära,
när det hade blivit något fel med eggen på skärorna eller plogbillarna, eller med gafflarna eller yxorna, eller när oxpikarnas uddar behövde rätas.
Härav kom sig, att när striden skulle stå, ingen enda av Sauls och Jonatans folk hade ett svärd eller ett spjut; allenast Saul själv och hans son Jonatan hade sådana.
Men filistéerna läto en utpost rycka fram till passet vid Mikmas.
Så hände sig nu en dag att Jonatan, Sauls son, sade till sin vapendragare: »Kom, låt oss gå över till filistéernas utpost där på andra sidan.»
Men han omtalade det icke för sin fader.
Saul vistades då vid Gibeas gräns, under granatträdet i Migron, och folket som han hade hos sig utgjorde vid pass sex hundra man;
och Ahia, son till Ahitub, som var broder till I-Kabod, son till Pinehas, son till Eli, HERRENS präst i Silo, har då efoden.
Och folket visste icke om, att Jonatan hade gått bort.
Men i passet, där Jonatan sökte gå över för att komma till filistéernas utpost, låg på vardera sidan en brant klippa; den ena hette Boses och den andra Sene.
Den ena klippan reste sig i norr, mitt emot Mikmas, den andra i söder, mitt emot Geba.
Och Jonatan sade till sin vapendragare: »Kom, låt oss gå över till dessa oomskurnas utpost, kanhända skall HERREN göra något för oss.
Ty intet hindrar HERREN att giva seger genom få likasåväl som genom många.»
Hans vapendragare svarade honom: »Gör allt vad du har i sinnet.
Gå du åstad; jag följer dig vart du vill.»
Då sade Jonatan: »Välan, vi skola gå över till männen där och laga så, att de få se oss.
Om de då säga till oss så: 'Stån stilla, till dess vi komma fram till eder', då skola vi stanna där vi äro och icke stiga upp till dem.
Om de däremot säga så: 'Kommen hitupp till oss', då skola vi stiga ditupp, ty då har HERREN givit dem i vår hand; detta skall för oss vara tecknet härtill.»
När nu de två hade blivit synliga för filistéernas utpost, sade filistéerna: »Se, hebréerna krypa ut ur hålen där de hava gömt sig.»
Därpå ropade utpostens manskap till Jonatan och hans vapendragare och sade: »Kommen hitupp till oss, så skola vi väl lära eder!»
Då sade Jonatan till sin vapendragare: »Följ mig ditupp, ty HERREN har givit dem i Israels hand.»
Och Jonatan klättrade på händer och fötter uppför, och hans vapendragare följde honom.
Och de föllo för Jonatan; och hans vapendragare gick efter honom och gav dem dödsstöten.
I det första anfallet nedgjorde så Jonatan och hans vapendragare vid pass tjugu män, på en sträcka av vid pass ett halvt plogland.
Då uppstod förskräckelse i lägret på fältet och bland allt folket; utposterna och de som hade gått ut för att härja grepos ock av förskräckelse.
Och marken darrade, så att en förskräckelse ifrån Gud uppstod.
Och Sauls väktare i Gibea i Benjamin fingo se att hopen var i upplösning, och att man sprang hit och dit.
Då sade Saul till folket som han hade hos sig: »Hållen mönstring och sen efter, vem som har gått ifrån oss.»
När de då höllo mönstring, funno de att Jonatan och hans vapendragare icke voro där.
Då sade Saul till Ahia: »För hit Guds ark.»
Ty Guds ark fanns på den tiden bland Israels barn.
Medan Saul ännu talade med prästen, tilltog larmet i filistéernas läger allt mer och mer.
Då sade Saul till prästen: »Låt det vara.»
Och Saul och allt det folk som han hade hos sig församlade sig och drogo till stridsplatsen; där fingo de se att den ene hade lyft sitt svärd mot den andre, så att en mycket stor förvirring hade uppstått.
Och de hebréer som sedan gammalt lydde under filistéerna, och som hade dragit hitupp med dem och voro här och där i lägret, dessa slöto sig nu ock till de israeliter som anfördes av Saul och Jonatan.
Och när de israeliter som hade gömt sig i Efraims bergsbygd hörde att filistéerna flydde, satte alla dessa också efter dem och deltogo i striden.
Så gav HERREN Israel seger på den dagen, och striden fortsattes ända bortom Bet-Aven.
När nu Israels män på den dagen voro hårt ansträngda, band Saul folket med följande ed: »Förbannad vare den man som förtär någon föda före aftonen, och innan jag har tagit hämnd på mina fiender.»
Så smakade då ingen av folket någon föda.
Och när de allasammans kommo in i skogsbygden, låg honung på marken.
Men när folket hade kommit in i skogsbygden och fått se den utflutna honungen, vågade dock ingen föra handen upp till munnen, ty folket fruktade för eden.
Jonatan däremot hade icke hört, när hans fader band folket med eden; därför räckte han ut staven som han hade i sin hand och doppade dess ända i honungskakan, och förde så handen till munnen; då kunde hans ögon åter se klart.
Men en man bland folket tog till orda och sade: »Din fader har bundit folket med en dyr ed och sagt: 'Förbannad vare den man som dag förtär någon föda.'»
Och folket var uttröttat.
Jonatan svarade: »Min fader har därmed dragit olycka över landet.
Sen huru klara mina ögon hava blivit, därför att jag smakade något litet av honungen här.
Huru mycket mer, om folket i dag hade fått äta sig mätta av bytet som de hade tagit från sina fiender -- huru mycket större skulle icke då filistéernas nederlag hava blivit!»
Emellertid slogo de filistéerna på den dagen och förföljde dem från Mikmas till Ajalon.
Och folket var mycket uttröttat.
Därför kastade sig folket över bytet och tog får, oxar och kalvar och slaktade dem på marken; och folket åt sedan köttet med blodet i.
När man berättade detta för Saul och sade: »Se, folket syndar mot HERREN genom att äta kött med blodet i», utropade han: »I haven handlat brottsligt.
Vältren nu fram till mig en stor sten.»
Och Saul sade vidare: »Gån ut bland folket och sägen till dem 'Var och en före fram till mig sin oxe och sitt får, och slakten dem här och äten; synden icke mot HERREN genom att äta köttet med blodet i.'»
Då förde allt folket, var och en med egen hand, om natten fram sina oxar och slaktade dem där.
Och Saul byggde ett altare åt HERREN; detta var det första altare som han byggde åt HERREN.
Och Saul sade: »Låt oss i natt draga ned och förfölja filistéerna och anställa plundring bland dem, ända till dess det bliver dager i morgon, och låt oss laga så, att ingen av dem bliver kvar.»
De svarade: »Gör allt vad dig täckes.»
Men prästen sade: »Låt oss träda fram hit till Gud.»
Då frågade Saul Gud: »Skall jag draga ned och förfölja filistéerna?
Vill du då giva dem i Israels hand?»
Men han gav honom intet svar den dagen.
Då sade Saul: »Kommen hitfram, alla I folkets förnämsta män, för att I mån få veta och se vari den synd består, som i dag har blivit begången.
Ty så sant HERREN lever, han som har givit Israel seger: om den ock vore begången av min son Jonatan, skall han döden dö.»
Men ingen bland allt folket svarade honom.
Då sade han till hela Israel: »Ställen I eder på ena sidan, så vill jag med min son Jonatan ställa mig på andra sidan.»
Folket svarade Saul: »Gör vad dig täckes.»
Och Saul sade till HERREN, »Israels Gud: »Låt sanningen komma i dagen.»
Då träffades Jonatan och Saul av lotten, och folket gick fritt.
Saul sade: »Kasten lott mellan mig och min son Jonatan.»
Då träffades Jonatan av lotten.
Saul sade till Jonatan: »Omtala för mig vad du har gjort.»
Då omtalade Jonatan det för honom och sade: »Med ändan av staven som jag hade i min hand tog jag litet honung och smakade därpå -- och så skall jag nu dö!»
Saul svarade: »Ja, Gud straffe mig nu och framgent: du måste döden dö, Jonatan.»
Men folket sade till Saul: »Skulle Jonatan dö, han som har förskaffat Israel denna stora seger?
Bort det!
Så sant HERREN lever, icke ett hår från hans huvud skall falla till jorden; ty med Guds hjälp har han i dag utfört detta.»
Och folket köpte Jonatan fri ifrån döden.
Och Saul drog hem, utan att vidare förfölja filistéerna; filistéerna begåvo sig ock hem till sitt.
När Saul nu hade tagit konungadömet över Israel i besittning, förde han krig mot alla sina fiender runt omkring: mot Moab, mot Ammons barn, mot Edom, mot konungarna i Soba och mot filistéerna; och vart han vände sig tuktade han dem.
Han gjorde mäktiga ting och slog Amalek och räddade så Israel från dess plundrares hand.
Sauls söner voro Jonatan, Jisvi och Malki-Sua; och av hans båda döttrar hette den äldre Merab och den yngre Mikal.
Sauls hustru hette Ahinoam, Ahimaas' dotter.
Hans härhövitsman hette Abiner, son till Ner, som var Sauls farbroder.
Ty Kis, Sauls fader, och Ner, Abners fader, voro söner till Abiel.
Men kriget mot filistéerna pågick häftigt, så länge Saul levde.
Och varhelst Saul såg någon rask och krigsduglig man tog han honom i sin tjänst.
Men Samuel sade till Saul: »Det var mig HERREN sände att smörja dig till konung över sitt folk Israel.
Så hör nu HERRENS ord.
Så säger HERREN Sebaot: Jag vill hemsöka Amalek för det som han gjorde mot Israel, att han lade sig i vägen för honom, när han drog upp ur Egypten.
Så drag nu åstad och slå amalekiterna och giv dem till spillo, med allt vad de hava, och skona dem icke, utan döda både män och kvinnor, både barn och spenabarn, både fäkreatur och får, både kameler och åsnor.»
Då bådade Saul upp folket och mönstrade dem i Telaim: två hundra tusen man fotfolk, och dessutom tio tusen man från Juda.
När Saul sedan kom till Amaleks stad, lade han ett bakhåll i dalen.
Men till kainéerna lät Saul säga: »Skiljen eder från amalekiterna och dragen ned, för att jag icke må utrota eder tillsammans med dem.
I bevisaden ju barmhärtighet mot alla Israels barn, när de drogo ut ur Egypten.»
Då skilde sig kainéerna från amalekiterna.
Och Saul slog amalekiterna och förföljde dem från Havila fram emot Sur, som ligger öster om Egypten.
Och han tog Agag, Amaleks konung, levande till fånga, och allt folket gav han till spillo, och han slog dem med svärdsegg.
Men Saul och folket skonade Agag, så ock det bästa och det näst bästa av får och fäkreatur jämte lammen, korteligen, allt som var av värde; sådant ville de icke giva till spillo.
All boskap däremot, som var dålig och mager, gåvo de till spillo.
Då kom HERRENS ord till Samuel; han sade:
»Jag ångrar att jag har gjort Saul till konung, ty han har vänt sig bort ifrån mig och icke fullgjort mina befallningar.»
Detta gick Samuel hårt till sinnes, och han ropade till HERREN hela den natten.
Och bittida om morgonen stod Samuel upp och gick för att möta Saul.
Då blev det berättat för Samuel att Saul hade kommit till Karmel och där rest åt sig en minnesstod, och att han sedan hade vänt om och dragit därifrån ned till Gilgal.
När nu Samuel kom till Saul, sade Saul till honom: »Välsignad vare du av HERREN.
Jag har nu fullgjort HERRENS befallning.»
Men Samuel sade: »Vad är det då för ett läte av får som ljuder i mina öron, och vad är det för ett läte av fäkreatur som jag hör?»
Saul svarade: »Från amalekiterna hava de fört dem med sig, ty folket skonade det bästa av fåren och fäkreaturen för att offra det åt HERREN, din Gud; men det övriga hava vi givit till spillo.»
Då sade Samuel till Saul: »Håll nu upp, så vill jag förkunna för dig vad HERREN i natt har talat till mig.
Han sade till honom: »Tala.»
Samuel sade: »Se, fastän du var ringa i dina egna ögon, har du blivit ett huvud för Israels stammar, ty HERREN smorde dig till konung över Israel.
Och HERREN sände dig åstad och sade: 'Gå och giv till spillo amalekiterna, de syndarna, och strid mot dem, till dess att du har förgjort dem.'
Varför har du då icke hört HERRENS röst, utan kastat dig över bytet och gjort vad ont är i HERRENS ögon?»
Saul svarade Samuel: »Jag har ju hört HERRENS röst och gått den väg på vilken HERREN har sänt mig.
Jag har fört hit Agag, Amaleks konung, och givit Amalek till spillo.
Men folket tog av bytet far och fäkreatur, det bästa av det tillspillogivna, för att offra det åt HERREN din Gud, i Gilgal.»
Då sade Samuel: »Menar du att HERREN har samma behag till brännoffer och slaktoffer som därtill att man hör HERRENS röst?
Nej, lydnad är bättre än offer, och hörsamhet bättre än det feta av vädurar.
Ty gensträvighet är trolldomssynd, och motspänstighet är avguderi och husgudsdyrkan.
Eftersom du har förkastat HERRENS ord, har han ock förkastat dig, och du skall icke längre vara konung.»
Saul sade till Samuel: »Jag har syndat därmed att jag har överträtt HERRENS befallning och handlat emot dina ord; ty jag fruktade för folket och lyssnade till deras ord.
Men förlåt mig nu min synd, och vänd tillbaka med mig, så att jag får tillbedja HERREN.»
Samuel sade till Saul: »Jag vänder icke tillbaka med dig; ty då du har förkastat HERRENS ord, har HERREN ock förkastat dig, så att du icke längre får vara konung över Israel.»
När nu Samuel vände sig om för att gå, fattade han i hörnet på hans mantel, och den rycktes sönder.
Och Samuel sade till honom: »HERREN har i dag ryckt Israels konungarike från dig och givit det åt en annan, som är bättre än du.
Och den Härlige i Israel ljuger icke och ångrar sig icke; ty han är icke en människa, så att han skulle kunna ångra sig.»
Han svarade: »Jag har syndat; men bevisa mig dock nu den äran inför de äldste i mitt folk och inför Israel, att du vänder tillbaka med mig, så att jag får tillbedja HERREN, din Gud.»
Då vände Samuel tillbaka och följde med Saul; och Saul tillbad HERREN.
Och Samuel sade: »Fören fram till mig Agag, Amaleks konung.»
Då gick Agag med glatt mod fram till honom.
Och Agag sade: »Välan, snart är dödens bitterhet överstånden.»
Men Samuel sade: »Såsom ditt svärd har gjort kvinnor barnlösa så skall ock din moder bliva barnlös framför andra kvinnor.»
Därpå högg Samuel Agag i stycken inför HERREN, i Gilgal.
Sedan begav sig Samuel till Rama; men Saul drog upp till sitt hem i Sauls Gibea.
Och Samuel ville icke mer se Saul så länge han levde, ty Samuel sörjde över Saul, eftersom HERREN ångrade att han hade gjort Saul till konung över Israel.
Och HERREN sade till Samuel: »Huru länge tänker du sörja över Saul?
Jag har ju förkastat honom, ty jag vill icke längre att han skall vara konung över Israel.
Fyll ditt horn med olja och gå åstad jag vill sända dig till betlehemiten Isai, ty en av hans söner har jag utsett åt mig till konung.»
Men Samuel sade: »Huru skall jag kunna gå dit?
Om Saul får höra det, så dräper han mig.»
HERREN svarade: »Tag en kviga med dig och säg: 'Jag har kommit för att offra åt HERREN.'
Sedan skall du inbjuda Isai till offret, och jag skall då själv låta dig veta vad du bör göra, och du skall smörja åt mig den jag säger dig.»
Samuel gjorde vad HERREN hade sagt, och kom så till Bet-Lehem Men när de äldste i staden fingo se honom, blevo de förskräckta och frågade: »Allt står väl rätt till?»
Han svarade: »Ja.
Jag har kommit för att offra åt HERREN.
Helgen eder och kommen med mig tid offret.»
Och han helgade Isai och hans söner och inbjöd dem till offret.
När de nu kommo dit och han fick se Eliab, tänkte han: »Förvisso står HERRENS smorde här inför honom.»
Men HERREN sade till Samuel »Skåda icke på hans utseende och på hans högväxta gestalt, ty jag har förkastat honom.
Ty det är icke såsom en människa ser; en människa ser på det som är för ögonen men HERREN ser till hjärtat.»
Då kallade Isai på Abinadab och lät honom gå fram för Samuel.
Men han sade: »Icke heller denne har HERREN utvalt.»
Då lät Isai Samma gå fram.
Men han sade: »Icke heller denne har HERREN utvalt.»
På detta sätt lät Isai sju av sina söner gå fram för Samuel; men Samuel sade till Isai: »HERREN har icke utvalt någon av dessa.»
Och Samuel frågade Isai: »Är detta alla ynglingarna?»
Han svarade: »Ännu återstår den yngste, men han går nu i vall med fåren.»
Då sade Samuel till Isai: »Sänd åstad och hämta hit honom, ty vi skola icke sätta oss till bords, förrän han kommer hit.»
Då sände han åstad och lät hämta honom, och han var ljuslätt och hade sköna ögon och ett fagert utseende.
Och HERREN sade: »Stå upp och smörj honom, ty denne är det.»
Då tog Samuel sitt oljehorn och smorde honom mitt ibland hans bröder; och HERRENS Ande kom över David, från den dagen och allt framgent.
Sedan stod Samuel upp och gick till Rama.
Men sedan HERRENS Ande hade vikit ifrån Saul, kvaldes han av en ond ande från HERREN.
Då sade Sauls tjänare till honom: »Eftersom en ond ande från Gud kväljer dig,
må du, vår herre, tillsäga dina tjänare, som stå inför dig, att de söka upp en man som är kunnig i harpospel, på det att han må spela på harpan, när den onde anden från Gud kommer över dig; så skall det bliva bättre med dig.»
Då sade Saul till sina tjänare: »Sen eder för min räkning om efter en man som är skicklig i strängaspel, och fören honom till mig.»
En av männen svarade då och sade: »Betlehemiten Isai har en son som jag har funnit vara kunnig i strängaspel, en käck stridsman och en förståndig man, därtill en fager man; och HERREN är med honom.»
Så sände då Saul bud till Isai och lät säga: »Sänd till mig din son David, som vaktar fåren.»
Då tog Isai en åsna, som han lastade med bröd, vidare en vinlägel och en killing, och sände detta med sin son David till Saul.
Så kom David till Saul och trädde i hans tjänst och blev honom mycket kär, så att han fick bliva hans vapendragare.
Och Saul sände till Isai och lät säga: »Låt David stanna kvar i min tjänst, ty han har funnit nåd för mina ögon.»
När nu anden från Gud kom över Saul, tog David harpan och spelade; då kände Saul lindring, och det blev bättre med honom, och den onde anden vek ifrån honom.
Men filistéerna församlade sina härar till strid; de församlade sig vid det Soko som hör till Juda.
Och de lägrade sig mellan Soko och Aseka, vid Efes-Dammim.
Saul och Israels män hade ock församlat sig och lägrat sig i Terebintdalen; och de ställde upp sig till strid mot filistéerna.
Filistéerna stodo vid berget på ena sidan, och israeliterna stodo vid berget på andra sidan, så att de hade dalen emellan sig.
Då framträdde ur filistéernas skaror en envigeskämpe vid namn Goljat, från Gat; han var sex alnar och ett kvarter lång.
Han hade en kopparhjälm på sitt huvud och var klädd i ett fjällpansar, och hans pansar hade en vikt av fem tusen siklar koppar.
Och han hade benskenor av koppar och bar en lans av koppar på sin rygg.
Skaftet på hans spjut liknade en vävbom, och spetsen på spjutet höll sex hundra siklar järn.
Och hans sköldbärare gick framför honom.
Han trädde nu fram och ropade till Israels här och sade till dem: »Varför dragen I ut och ställen upp eder till strid?
Jag står här på filistéernas vägnar, och I ären Sauls tjänare; väljen nu ut åt eder en man som må komma hitned till mig.
Om han förmår strida mot mig och slår ned mig, så skola vi vara eder underdåniga; men om jag bliver hans överman och slår ned honom, så skolen I vara oss underdåniga och tjäna oss.»
Och filistéen sade ytterligare: »Jag har i dag smädat Israels här.
Skaffen nu hit någon, så att vi få strida med varandra!
Då Saul och hela Israel hörde dessa filistéens ord, blevo de gripna av förfäran och stor fruktan.
Men David var son till den omtalade efratiten från Bet-Lehem i Juda, som hette Isai och hade åtta söner; denne var på Sauls tid en gammal man vid framskriden ålder.
Nu hade Isais tre äldsta söner dragit åstad och följt med Saul ut i kriget.
Av dessa hans tre söner, som hade dragit ut i kriget, hette den förstfödde Eliab, hans andre son Abinadab och den tredje Samma.
David var den yngste.
De tre äldsta hade nu följt med Saul.
Men David lämnade understundom Saul och gick hem för att vakta sin faders får i Bet-Lehem.
Och filistéen kom fram både bittida och sent; i fyrtio dagar kom han och ställde sig där.
Nu sade Isai en gång till sin son David: »Tag för dina bröders räkning en efa av dessa rostade ax jämte dessa tio bröd, och skaffa detta skyndsamt till dina bröder i lägret.
Och dessa tio ostar skall du föra till deras överhövitsman.
Du skall se efter, om det står väl till med dina bröder, och begära av dem en mottagningspant.
Saul och de och alla Israels män äro nämligen i Terebintdalen och strida mot filistéerna.»
Bittida följande morgon överlämnade David fåren åt en vaktare, tog med sig vad han skulle och begav sig åstad, såsom Isai hade bjudit honom.
När han kom fram till vagnborgen, hov hären, som då skulle draga ut i slagordning, upp sitt härskri.
Och Israel och filistéerna ställde upp sig i slagordning mot varandra.
Då lämnade David ifrån sig sakerna åt trossvaktaren och skyndade bort till hären; och när han kom dit, hälsade han sina bröder.
Under det att han talade med dem, trädde nu envigeskämpen, han som hette Goljat, filistéen ifrån Gat, fram ur filistéernas här och talade såsom förut; och David hörde det.
Och alla Israels män flydde för mannen, när de fingo se honom och fruktade storligen.
Och Israels män sade: »Sen I mannen där, som nu träder upp?
Han träder upp för att smäda Israel.
Men den man som slår ned honom vill konungen begåva med stor rikedom, och åt honom vill han giva sin dotter, och hans faders hus vill han göra skattefritt i Israel.»
Och David sade till de man som stodo bredvid honom: »Vad får den man som slår ned denne filisté och därmed tager bort sådan smälek från Israel?
Ty vem är denne oomskurne filisté, som vågar smäda den levande Gudens här?»
Folket upprepade då för honom det som nyss hade blivit sagt; de sade: »Detta får den man som slår ned honom.»
Men Eliab, hans äldste broder, hörde huru han talade med männen; då upptändes Eliabs vrede mot David, och han sade: »Varför har du kommit hitned, och åt vem har du överlämnat den lilla fårhjorden där i öknen?
Jag känner ditt övermod och ditt hjärtas ondska; för att se på striden är det som du har kommit hitned.»
David svarade: »Vad har jag då gjort?
Det var ju allenast en fråga.»
Sedan vände han sig ifrån honom till en annan och upprepade sin fråga, och folket gav honom samma svar som förut.
Men vad David hade talat blev bekant; och man berättade det för Saul, och denne lät hämta honom.
Och David sade till Saul: »Må ingen låta sitt mod falla.
Din tjänare vill gå åstad och strida mot denne filisté.»
Saul sade till David: »Icke kan du gå åstad mot denne filisté och strida mot honom; du är du ju allenast en yngling, och han är en stridsman allt ifrån ungdomen.»
Men David svarade Saul: »Din tjänare har gått i vall med sin faders får; om då ett lejon eller en björn kom och tog bort ett får av hjorden,
så följde jag efter vilddjuret och slog ned det och ryckte rovet ur munnen på det; och om det då reste sig upp mot mig, så fattade jag det i skägget och slog ned det och dödade det.
Har nu din tjänare slagit ned både lejon och björn, så skall det gå denne oomskurne filisté såsom det gick vart och ett av dessa djur, ty han har smädat den levande Gudens här.»
Och David sade ytterligare: »HERREN, som räddade mig undan lejon och björn, han skall ock rädda mig undan denne filisté.»
Då sade Saul till David: »Gå då åstad; HERREN skall vara med dig.»
Och Saul klädde på David sina egna kläder och satte en kopparhjälm på hans huvud och klädde på honom ett pansar.
Och David omgjordade sig med hans svärd utanpå kläderna och prövade på att gå därmed, ty han hade aldrig försökt något sådant.
Och David sade till Saul: »Jag kan icke gå så klädd, ty jag har aldrig försökt sådant.»
Därpå lade David det av sig.
Och han tog sin stav i handen och valde ut åt sig fem släta stenar ur bäcken och lade dem i sin herdeväska och i barmen, och tog sin slunga i handen; därefter gick han fram mot filistéen.
Och filistéen gick framåt och kom David allt närmare, och hans sköld bärare gick framför honom.
Då nu filistéen såg upp och fick se David, föraktade han honom; ty denne var ännu en yngling, ljuslätt och skön.
Och filistéen sade till David: »Menar du att jag är en hund, eftersom du kommer emot mig med käppar?»
Och filistéen förbannade David, i det han svor vid sina gudar.
Sedan sade filistéen till David: »Kom hit till mig, så skall jag giva ditt kött åt himmelens fåglar och åt markens djur.»
David svarade filistéen: »Du kommer mot mig med svärd och spjut och lans, men jag kommer mot dig i HERREN Sebaots namn, hans som är Israels härs Gud, den härs som du har smädat.
HERREN skall denna dag överlämna dig i min hand, så att jag skall slå ned dig och taga ditt huvud av dig, och jag skall denna dag giva de filisteiska krigarnas döda kroppar åt himmelens fåglar och åt jordens vilda djur; så skola alla länder förnimma att Israel har en Gud.
Och hela denna hop skall förnimma att det icke är genom svärd och spjut som HERREN giver seger; ty striden är HERRENS, och han skall giva eder i vår hand.»
När då filistéen gjorde sig redo och gick framåt och närmade sig David, sprang David med hast fram mot hären, filistéen till mötes.
Och David stack sin hand i väskan och tog därur en sten och slungade och träffade filistéen i pannan; och stenen trängde in i pannan, så att han föll omkull med ansiktet mot jorden.
Så övervann David filistéen med slunga och sten och slog filistéen till döds,
utan att David därvid hade något svärd i sin hand.
Sedan sprang David fram och ställde sig invid filistéen och fattade i hans svärd; och när han hade dragit det ut ur skidan, gav han honom dödsstöten och högg av hans huvud därmed.
När filistéerna nu sågo att deras kämpe var död, flydde de.
Men Israels och Juda man stodo upp och höjde ett härskri och förföljde filistéerna ända dit där vägen går till Gai, och ända intill Ekrons portar; och filistéer föllo och lågo slagna på vägen till Saaraim, och sedan ända till Gat och ända till Ekron.
Sedan Israels barn sålunda häftigt hade förföljt filistéerna, vände de tillbaka och plundrade deras läger.
Och David tog filistéens huvud och förde det till Jerusalem, men hans vapen lade han i sitt tält.
När Saul såg David gå ut mot filistéen, frågade han härhövitsmannen Abner: »Vems son är denne yngling, Abner?»
Abner svarade: »Så sant du lever, konung, jag vet det icke.»
Då sade konungen: »Hör då efter, vems son den unge mannen är.»
När sedan David vände tillbaka, efter att hava slagit ihjäl filistéen, tog Abner honom med sig och förde honom inför Saul, medan han ännu hade filistéens huvud i sin hand.
Då sade Saul till honom: »Vems son är du, yngling» David svarade: »Din tjänare Isais, betlehemitens, son.»
Sedan, efter det att David hade talat ut med Saul, fäste sig Jonatans hjärta så vid Davids hjärta, att Jonatan hade honom lika kär som sitt eget liv.
Och Saul tog honom till sig på den dagen och lät honom icke mer vända tillbaka till sin faders hus.
Och Jonatan slöt ett förbund med David, då han nu hade honom lika kär som sitt eget liv.
Och Jonatan tog av sig manteln som han hade på sig och gav den åt David, så ock sina övriga kläder, ända till sitt svärd, sin båge och sitt bälte
Och när David drog ut, hade han framgång överallt dit Saul sände honom; Saul satte honom därför över krigsfolket.
Och allt folket fann behag i honom, också de som voro Sauls tjänare.
Och när de kommo hem, då David vände tillbaka, efter att hava slagit ned filistéen, gingo kvinnorna ut från alla Israels städer, under sång och dans, för att möta konung Saul med jubel, med pukor och trianglar.
Och kvinnorna sjöngo med fröjd sålunda: »Saul har slagit sina tusen, men David sina tio tusen.»
Då blev Saul mycket vred, ty det talet misshagade honom, och han sade: »Åt David hava de givit tio tusen, och åt mig hava de givit tusen; nu fattas honom allenast konungadömet.»
Och Saul såg med ont öga på David från den dagen och allt framgent.
Dagen därefter kom en ond ande från Gud över Saul, så att han rasade i sitt hus; men David spelade på harpan, såsom han dagligen plägade.
Och Saul hade sitt spjut i handen.
Och Saul svängde spjutet och tänkte: »Jag skall spetsa David fast vid väggen.»
Men David böjde sig undan för honom, två gånger.
Och Saul fruktade för David, eftersom HERREN var med honom, sedan han hade vikit ifrån Saul.
Därför avlägsnade Saul honom ifrån sig, i det att han gjorde honom till överhövitsman i sin här; han blev så folkets ledare och anförare.
Och David hade framgång på alla sina vägar, och HERREN var med honom.
Då nu Saul såg att han hade så stor framgång, fruktade han honom än mer.
Men hela Israel och Juda hade David kär, eftersom han var deras ledare och anförare.
Och Saul sade till David: »Se, min äldsta dotter, Merab, vill jag giva dig till hustru; skicka dig allenast såsom en tapper man i min tjänst, och för HERRENS krig.»
Ty Saul tänkte: »Min hand må icke drabba honom, filistéernas hand må drabba honom.»
Men David svarade Saul: »Vem är jag, vilka hava mina levnadsförhållanden varit, och vad är min faders släkt i Israel, eftersom jag skulle bliva konungens måg?»
När tiden kom att Sauls dotter Merab skulle hava givits åt David, blev hon emellertid given till hustru åt meholatiten Adriel. --
Men Sauls dotter Mikal hade David kär.
Och när man omtalade detta för Saul, behagade det honom.
Saul tänkte nämligen: »Jag skall giva henne åt honom, för att hon må bliva honom en snara, så att filistéernas hand drabbar honom.»
Och Saul sade till David: »För andra gången kan du nu bliva min måg.»
Och Saul bjöd sina tjänare att de hemligen skulle tala så med David: »Se, konungen har behag till dig, och alla hans tjänare hava dig kär; du hör nu bliva konungens måg.»
Och Sauls tjänare talade dessa ord i Davids öron.
Men David sade: »Tyckes det eder vara en så ringa sak att bliva konungens måg?
Jag är ju en fattig och ringa man.»
Detta omtalade Sauls tjänare för honom och sade: »Så har David sagt.»
Då tillsade Saul dem att de skulle säga så till David: »Konungen begär ingen annan brudgåva än förhudarna av ett hundra filistéer, för att hämnd så må tagas på konungens fiender.»
Saul hoppades nämligen att han skulle få David fälld genom filistéernas hand.
När så hans tjänare omtalade för David vad han hade sagt, ville David gärna på det villkoret bliva konungens måg; och innan tiden ännu var förlupen,
stod David upp och drog åstad med sina män och slog av filistéerna två hundra man.
Och David tog deras förhudar med sig, och fulla antalet blev överlämnat åt konungen, för att han skulle bliva konungens måg.
Och Saul gav honom så sin dotter Mikal till hustru.
Men Saul såg och förstod att HERREN var med David; Och Sauls dotter Mikal hade honom kär.
Då fruktade Saul ännu mer för David, och så blev Saul Davids fiende för hela livet.
Men filistéernas furstar drogo i fält; och så ofta de drogo ut, hade David större framgång än någon annan av Sauls tjänare, så att hans namn blev mycket berömt.
Och Saul talade med sin son Jonatan och med alla sina tjänare om att döda David; men Sauls son Jonatan var David mycket tillgiven.
Därför omtalade Jonatan detta för David och sade: »Min fader Saul söker att döda dig.
Tag dig alltså till vara i morgon och håll dig gömd på någon plats där du kan vara dold.
Men själv vill jag gå ut och ställa mig bredvid min fader på marken, där du är, och jag vill tala om dig med min fader; om jag då märker något, skall jag sedan omtala det för dig.
Och Jonatan talade till Davids bästa med sin fader Saul och sade till honom: »Konungen må icke försynda sig på sin tjänare David ty han har icke försyndat sig mot dig, utan vad han har gjort har varit till stort gagn för dig.
Han tog ju sin själ i sin hand och slog ned filistéen, och HERREN gav så hela Israel en stor seger; du har själv sett det och glatt dig däråt.
Varför skulle du då försynda dig på oskyldigt blod genom att döda David utan sak?»
Och Saul lyssnade till Jonatans ord; och Saul svor: »Så sant HERREN lever, han skall icke dödas.»
Sedan kallade Jonatan David till sig; och Jonatan omtalade för honom allt som hade blivit sagt.
Därefter förde Jonatan David till Saul, och han var i hans tjänst såsom förut.
När så kriget åter begynte, drog David ut och stridde mot filistéerna och tillfogade dem ett stort nederlag, så att de flydde för honom.
Men en ond ande från HERREN kom över Saul, där han satt i sitt hus med spjutet i handen, under det att David spelade på harpan.
Då sökte Saul att med spjutet spetsa David fast vid väggen; men denne vek undan för Saul, så att han allenast stötte spjutet in i väggen.
Och David flydde och kom undan samma natt.
Emellertid sände Saul till Davids hus några män med uppdrag att vakta på honom och att sedan om morgonen döda honom.
Men Mikal, Davids hustru, omtalade detta för honom och sade: »Om du icke i natt räddar ditt liv, så är du i morgon dödens man.»
Därefter släppte Mikal ned David genom fönstret; och han begav sig på flykten och kom så undan.
Sedan tog Mikal husguden och lade honom i sängen och satte myggnätet av gethår över huvudgärden och höljde täcket över honom.
När sedan Saul sände sina män med uppdrag att hämta David, sade hon: »Han är sjuk.»
Då sände Saul dit männen med uppdrag att skaffa sig tillträde till David själv och sade: »Bären honom i sängen hitupp till mig, så att jag får döda honom.»
Men när männen kommo in, fingo de se att det var husguden som låg i sängen, med myggnätet över huvudgärden.
Då sade Saul till Mikal: »Varför har du så bedragit mig och släppt min fiende, så att han har kommit undan?»
Mikal svarade Saul: »Han sade till mig: 'Släpp mig; eljest dödar jag dig.'»
När David nu hade flytt och kommit undan, begav han sig till Samuel i Rama och omtalade för denne allt vad Saul hade gjort honom.
Och han och Samuel gingo till Najot och stannade där.
Och det blev berättat för Saul att David var i Najot vid Rama.
Då sände Saul dit några män med uppdrag att hämta David.
Men när Sauls utskickade fingo se skaran av profeterna i profetisk hänryckning, och fingo se Samuel stå där såsom deras anförare, kom Guds Ande över dem, så att också de fattades av hänryckning.
När man omtalade detta för Saul, sände han dit andra män; men också de fattades av hänryckning.
Och när han då ytterligare, för tredje gången, sände dit män med samma uppdrag, fattades också dessa av hänryckning.
Då begav han sig själv till Rama; och när han kom till den stora brunnen i Seku, frågade han: »Var äro Samuel och David?»
Man svarade: »De äro i Najot vid Rama.»
Då begav han sig dit, till Najot vid Rama.
Men Guds Ande kom också över honom, så att han hela vägen gick i profetisk hänryckning, ända till dess att han kom fram till Najot vid Rama.
Då kastade också han av sig sina kläder, i det att också han blev fattad av hänryckning inför Samuel; och han föll ned och låg där naken hela den dagen och hela natten.
Därför plägar man säga: »Är ock Saul bland profeterna?»
Men David flydde från Najot vid Rama och kom till Jonatan och sade: »Vad har jag gjort?
Vilken missgärning, vilken synd har jag begått mot dig fader, eftersom han står efter mitt liv?»
Han svarade honom: »Bort det!
Du skall icke dö.
Min fader gör ju intet, varken något viktigt eller något oviktigt, utan att uppenbara det för mig.
Varför skulle då min fader dölja detta för mig?
Nej, så skall icke ske.»
Men David betygade ytterligare med ed och sade: »Din fader vet väl att jag har funnit nåd för dina ögon; därför tänker han: 'Jonatan skall icke få veta detta, på det att han icke må bliva bedrövad.'
Men så sant HERREN lever, och så sant du själv lever: det är icke mer än ett steg mellan mig och döden.»
Då sade Jonatan till David: »Vadhelst du önskar skall jag göra för dig.»
David sade till Jonatan: »I morgon är ju nymånad, och jag skulle då rätteligen sitta till bords med konungen; men låt mig nu gå och gömma mig ute på marken till i övermorgon afton.
Om då din fader saknar mig, så säg: 'David utbad sig tillstånd av mig att få göra ett hastigt besök i sin stad, Bet-Lehem, där hela släkten nu firar sin årliga offerfest.'
Om han då säger: 'Gott!', så kan din tjänare vara trygg.
Men om han bliver vred, så märker du därav att han har beslutit min ofärd.
Visa så din nåd mot din tjänare, eftersom du har låtit din tjänare ingå ett HERRENS förbund med dig.
Men om det finnes någon missgärning hos mig, så döda mig du, ty varför skulle du föra mig till din fader?»
Då sade Jonatan: »Bort det!
Om jag märker att min fader har beslutit att låta ofärd komma över dig, skall jag förvisso omtala det för dig.»
Men David sade till Jonatan: »Vem skall omtala för mig detta, eller säga mig om din fader giver dig ett hårt svar?»
Jonatan sade till David: »Kom, låt oss gå ut på marken.»
Och de gingo båda ut på marken.
Och Jonatan sade till David: »Vid HERREN» Israels Gud: om jag finner att det låter gott för David, när jag i morgon eller i övermorgon vid denna tid utforskar min fader, så skall jag förvisso sända bud till dig och uppenbara det för dig.
HERREN straffe Jonatan nu och framgent, om jag, såframt min fader åstundar din ofärd, icke uppenbarar det för dig och låter dig komma undan, så att du får gå dina färde i trygghet.
Och HERREN vare då med dig, såsom han har varit med min fader.
Och nog skall du väl, om jag då ännu är i livet, ja, nog skall du väl bevisa barmhärtighet mot mig, såsom HERREN är barmhärtig, så att jag slipper att dö?
Icke skall du väl någonsin taga bort din barmhärtighet från mitt hus, icke ens då när HERREN har tagit bort alla Davids fiender ifrån jorden?»
Jonatan slöt då ett förbund med Davids hus; och HERREN utkrävde sedan av Davids fiender vad de hade förskyllt.
Och Jonatan besvor David ytterligare vid sin kärlek till honom, ty han hade honom lika kär som han hade sitt eget liv;
Jonatan sade till honom: »I morgon är nymånad, och du skall då saknas, ty din plats kommer ju att stå tom.
Men gå i övermorgon skyndsamt ned till den plats där du gömde dig den dag då ogärningen skulle hava skett, och uppehåll dig bredvid Eselstenen.
Jag vill då själv i dess närhet avskjuta mina tre pilar, såsom sköte jag till måls.
Sedan skall jag skicka min tjänare att gå och söka upp pilarna.
Om jag då säger till tjänaren: »Se, pilarna ligga bakom dig, närmare hitåt', så tag du upp dem och kom fram, ty då kan du vara trygg och ingenting är på färde, så sant HERREN lever.
Men om jag säger så till den unge mannen: 'Se, pilarna ligga framför dig, längre bort', så gå dina färde, ty då sänder HERREN dig bort.
Och i fråga om det som jag och du nu hava talat, är HERREN vittne mellan mig och dig till evig tid.»
Och David gömde sig ute på marken.
Och när nymånaden var inne, satte konungen sig till bords för att äta.
Konungen satte sig på sin vanliga sittplats, platsen vid väggen; och Jonatan stod upp, och Abner satte sig vid Sauls sida.
Men Davids plats stod tom.
Saul sade dock intet den dagen, ty han tänkte: »Något har hänt honom; han är nog icke ren, säkerligen är han icke ren.»
Men när Davids plats stod tom också dagen efter nymånadsdagen, dagen därefter, sade Saul till sin son Jonatan: »Varför har Isais son varken i går eller i dag kommit till måltiden?»
Jonatan svarade Saul: »David utbad sig tillstånd av mig att få gå till Bet-Lehem;
han sade: 'Låt mig gå, ty vi fira en släktofferfest i staden, och min broder har själv bjudit mig att komma; om jag har funnit nåd för dina ögon, så låt mig nu slippa härifrån för att besöka mina bröder.'
Därför har han icke kommit till konungens bord.»
Då upptändes Sauls vrede mot Jonatan, och han sade till honom: »Du son till en otuktig kvinna!
Visste jag då icke att du hade funnit behag i Isais son, till skam för dig själv och till skam för din moders blygd!
Ty så länge Isais son lever på jorden, är varken du eller din konungamakt säker.
Sänd därför nu åstad och låt hämta honom hit till mig, ty han är dödens barn.»
Jonatan svarade sin fader Saul och sade till honom: »Varför skall han dödas?
Vad har han gjort?»
Då svängde Saul spjutet mot honom för att genomborra honom; och nu märkte Jonatan att hans fader hade beslutit att döda David.
Och Jonatan stod upp från bordet i vredesmod och åt intet på den andra nymånadsdagen, ty han var bedrövad för Davids skull, därför att hans fader hade gjort sådan orätt mot denne.
Följande morgon gick Jonatan ut på marken, vid den tid han hade utsatt för David; och han hade en liten gosse med sig.
Och han sade till gossen: »Spring och sök reda på pilarna som jag skjuter av.»
Medan nu gossen sprang, sköt han pilen över honom.
Och när gossen kom till det ställe dit Jonatan hade avskjutit pilen, ropade Jonatan efter gossen och sade: »Pilen ligger ju framför dig, längre bort.»
Och Jonatan ropade ytterligare efter gossen: »Fort, skynda dig, stanna icke!»
Och gossen som Jonatan hade med sig tog upp pilen och kom till sin herre.
Men gossen visste icke varom fråga var; allenast Jonatan och David visste det.
Och Jonatan lämnade sina vapen åt gossen som han hade med sig och sade till honom: »Gå och bär dem in i staden.»
Men sedan gossen hade gått, reste David sig upp på södra sidan; och han föll ned till jorden på sitt ansikte och bugade sig tre gånger; och de kysste varandra och gräto med varandra, och David grät överljutt.
Och Jonatan sade till David: »Gå i frid.
Blive det såsom vi båda svuro vid HERRENS namn, när vi sade: 'HERREN vare vittne mellan mig och dig, mellan mina efterkommande och dina, till evig tid.'»
Sedan stod han upp och gick sina färde, men Jonatan gick in i staden igen.
Och David kom till prästen Ahimelek i Nob.
Men Ahimelek blev förskräckt, när han fick se David, och frågade honom: »Varför kommer du ensam och har ingen med dig?»
David svarade prästen Ahimelek: »Konungen har givit mig ett uppdrag, men han sade till mig: 'Ingen får veta något om det uppdrag vari jag sänder dig, och som jag har givit dig.'
Och mina män har jag visat till det och det stället.
Giv mig nu vad du har till hands, fem bröd eller vad som kan finnas.»
Prästen svarade David och sade »Vanligt bröd har jag icke till hands; allenast heligt bröd finnes -- om eljest dina män hava avhållit sig från kvinnor.»
David svarade prästen och sade till honom: »Ja, sannerligen, kvinnor hava på sista tiden varit skilda från oss; när jag drog åstad, voro ock mina mäns tillhörigheter heliga.
Därför, om också vårt förehavande är av helt vanligt slag, är det dock i dag heligt, vad våra tillhörigheter angår.»
Då gav prästen honom av det heliga; ty där fanns icke något annat bröd än skådebröden, som hade legat inför HERRENS ansikte, men som man hade burit undan, för att lägga fram nybakat bröd samma dag det gamla togs bort.
Men där befann sig den dagen en av Sauls tjänare, som var satt i förvar inför HERREN, en edomé vid namn Doeg, den förnämste av Sauls herdar.
Och David frågade Ahimelek ytterligare: »Har du icke här till hands något spjut eller något svärd?
Ty varken mitt svärd eller mina andra vapen tog jag med mig, eftersom konungens uppdrag krävde så stor skyndsamhet.»
Prästen svarade: »Jo, det svärd som har tillhört filistéen Goljat, honom som du slog ned i Terebintdalen; det finnes, inhöljt i ett kläde, där bakom efoden.
Vill du taga det med dig, så tag det; ty något annat än det har jag icke.»
David sade: »Dess like finnes icke; giv mig det.»
Och David stod upp och flydde samma dag för Saul och kom till Akis, konungen i Gat.
Men Akis' tjänare sade till honom: »Detta är ju David, landets konung!
Det är ju till dennes ära man sjunger så under dansen: 'Saul har slagit sina tusen, men David sina tio tusen.'
David lade märke till dessa ord, och han begynte storligen frukta för Akis, konungen i Gat.
Därför ställde han sig vansinnig inför deras ögon och betedde sig såsom en ursinnig, när de ville fasthålla honom, och ritade på dörrarna i porten och lät spotten rinna ned i sitt skägg.
Då sade Akis till sina tjänare: »I sen ju huru vanvettigt mannen beter sig.
Varför fören I honom till mig?
Har jag då sådan brist på vanvettiga människor, att I behövden föra denne hit, för att han skulle bete sig vanvettigt inför mig?
Skulle en sådan få komma in i mitt hus?»
Då begav sig David därifrån och flydde undan till Adullams grotta.
Och när hans bröder och hela hans faders hus fingo höra detta, kommo de ditned till honom.
Och till honom församlade sig alla slags män som voro i något trångmål, alla som ansattes av fordringsägare och alla missnöjda, och han blev deras hövding; vid pass fyra hundra man slöto sig så till honom.
Därifrån begav sig David till Mispe i Moab.
Och han sade till konungen i Moab: »Låt min fader och min moder få komma hitöver och vara hos eder till dess jag får veta vad Gud vill göra med mig.»
Och han förde dem fram inför konungen i Moab; och de fingo stanna hos denne, så länge David var på borgen.
Men profeten Gad sade till David: »Du skall icke stanna här på borgen; drag bort härifrån och begiv dig in i Juda land.»
Då drog David bort därifrån och kom till Heretskogen.
Och Saul fick höra att man hade fått spaning på David och de män som voro med honom.
Då nu Saul en dag satt i Gibea under tamarisken på höjden, med sitt spjut i handen, under det att alla hans tjänare stodo omkring honom,
sade han till sina tjänare, där de stodo omkring honom: »Hören, I benjaminiter.
Skall då också Isais son åt eder alla giva åkrar och vingårdar och göra eder alla till över- och underhövitsmän?
Ty I haven ju alla sammansvurit eder mot mig, och ingen har uppenbarat för mig att min son har slutit förbund med Isais son.
Ingen av eder bekymrar sig så mycket om mig, att han har uppenbarat det för mig.
Min son har ju uppeggat min tjänare till att stämpla mot mig, såsom nu sker.»
Edoméen Doeg, som ock stod där bland Sauls tjänare, svarade då och sade: »Jag har sett Isais son komma till Ahimelek, Ahitubs son, i Nob.
Denne frågade då HERREN för honom och gav honom reskost; han gav honom ock filistéen Goljats svärd.»
Då sände konungen och lät kalla till sig prästen Ahimelek, Ahitubs son, och hela hans faders hus, prästerna i Nob.
Och de kommo alla till konungen.
Då sade Saul: »Hör mig, du Ahitubs son.»
Han svarade: »Jag hör dig, min herre.»
Saul sade till honom: »Varför haven I sammansvurit eder mot mig, du och Isais son, i det att du har givit honom bröd och svärd och frågat Gud för honom, så att han skulle kunna sätta sig upp mot mig och stämpla mot mig, såsom nu sker?»
Ahimelek svarade konungen och sade: »Vem bland alla dina tjänare är väl så betrodd som David, han som därtill är konungens måg och hövding för din livvakt och högt ärad i ditt hus?
Är det då nu för första gången som jag har frågat Gud för honom?
Bort det!
Icke må konungen lägga mig, sin tjänare, och hela min faders hus något till last, ty din tjänare visste alls intet om allt detta.»
Men konungen sade: »Du måste döden dö, Ahimelek, du själv och hela din faders hus.»
Och konungen sade till drabanterna som stodo där omkring honom: »Träden fram och döden HERRENS präster; ty också de hålla med David; och fastän de visste att han flydde, uppenbarade de det icke för mig.»
Men konungens tjänare ville icke uträcka sina händer till att stöta ned HERRENS präster.
Då sade konungen till Doeg: »Träd du fram och stöt ned prästerna.»
Edoméen Doeg trädde då fram och stötte ned prästerna och dödade på den dagen åttiofem män som buro linne-efod.
Och invånarna i präststaden Nob blevo slagna med svärdsegg, både män och kvinnor, både barn och spenabarn; också fäkreatur, åsnor och får blevo slagna med svärdsegg.
Allenast en son till Ahimelek, Ahitubs son, vid namn Ebjatar, kom undan, och denne flydde bort till David.
Och Ebjatar omtalade för David att Saul hade dräpt HERRENS präster.
Då sade David till Ebjatar: »Jag förstod redan då att edoméen Doeg, eftersom han var där, skulle omtala allt för Saul.
Det är jag som är orsaken till att hela din faders hus har förgåtts.
Bliv kvar hos mig, frukta intet; ty den som står efter mitt liv, han står ock efter ditt liv.
Hos mig är du i gott förvar.»
Och man berättade för David: »Filistéerna hålla nu på att belägra Kegila, och de plundra logarna.»
Då frågade David HERREN: »Skall jag draga åstad och slå dessa filistéer?»
HERREN svarade David: »Drag åstad och slå filistéerna och fräls Kegila.»
Men Davids män sade till honom: »Vi leva ju i fruktan redan här i Juda.
Och nu skulla vi därtill draga åstad till Kegila, mot filistéernas här!»
Då frågade David HERREN ännu en gång, och HERREN svarade honom och sade: »Stå upp och drag ned till Kegila; ty jag vill giva filistéerna i din hand.»
Då drog David med sina män till Kegila och stridde mot filistéerna och förde bort deras boskap och tillfogade dem ett stort nederlag.
Så frälste David invånarna i Kegila.
När Ebjatar, Ahimeleks son, flydde till David i Kegila, förde han efoden med sig ditned.
Och det blev berättat för Saul att David hade dragit in i Kegila.
Då sade Saul: »Gud har förkastat honom och givit honom i min hand, ty han har själv stängt in sig genom att gå in i en stad med portar och bommar.»
Därefter bådade Saul upp allt folket till strid, för att draga ned till Kegila och där innesluta David och hans man.
Men när David fick veta att Saul stämplade ont mot honom, sade han till prästen Ebjatar: »Bär hit efoden.»
Och David sade: »HERRE, Israels Gud, din tjänare har hört att Saul har i sinnet att komma mot Kegila och fördärva staden för min skull.
Skola Kegilas borgare då utlämna mig åt honom?
Skall Saul komma hitned, såsom din tjänare har hört?
HERRE, Israels Gud, förkunna det för din tjänare.»
HERREN svarade: »Han skall komma hitned.»
David frågade ytterligare: »Skola Kegilas borgare då utlämna mig och mina man åt Saul?»
HERREN svarade: »De skola utlämna eder.»
Då bröt David upp med sitt folk, som utgjorde vid pass sex hundra man, och de drogo ut från Kegila och vandrade vart de kunde.
När det då blev berättat för Saul att David hade flytt undan från Kegila avstod han från att draga ut.
Så uppehöll sig nu David i öknen på bergfästena; han uppehöll sig bland bergen i öknen Sif.
Och Saul sökte alltjämt efter honom, men Gud gav honom icke i hans hand.
Och medan David var i Hores i öknen Sif, förnam han att Saul hade dragit ut för att söka döda honom.
Men Jonatan, Sauls son, stod upp och gick till David i Hores och styrkte hans mod i Gud.
Han sade till honom: »Frukta icke; ty min fader Sauls hand skall icke träffa dig, utan du skall bliva konung över Israel, och jag skall då hava andra platsen, näst efter dig.
Detta vet ock min fader Saul.»
Sedan slöto de båda ett förbund inför HERREN.
Och David stannade kvar i Hores, men Jonatan gick hem igen.
Men några sifiter drogo upp till Saul i Gibea och sade: »David håller sig nu gömd hos oss på bergfästena i Hores, på Hakilahöjden, som ligger söder om ödemarken.
Så drag nu ditned, o konung, så snart det lyster dig att göra det. står sak bliver det då att utlämna honom åt konungen.»
Då sade Saul: »Varen välsignade av HERREN, därför att I haven velat spara mig bekymmer.
Men gån nu och skaffen eder ytterligare visshet, och tagen reda på och sen efter, på vilket ställe han nu vistas, och vem som har sett honom där; ty man har sagt mig att han är mycket listig.
Och sen efter och tagen reda på alla gömställen där han kan gömma sig; och kommen så igen till mig, när I haven fått visshet, så vill jag sedan gå med eder.
Ty finnes han i landet, skall jag veta att söka upp honom, om jag än måste söka bland alla Juda ätter.»
Då stodo de upp och gingo till Sif före Saul.
Men David och hans män voro i öknen Maon, på hedmarken, söder om ödemarken.
När nu Saul drog åstad med sina män för att söka efter David, om talade man det för denne, och han drog då ned till klippan och stannade så i öknen Maon.
När Saul hörde detta, satte han efter David in i öknen Maon.
Och Saul gick på ena sidan om berget, och David med sina män på andra sidan.
Men just som David var stadd på flykt för att komma undan Saul, under det att Saul och hans män sökte kringränna David och hans män för att taga dem till fånga
kom en budbärare till Saul och sade: »Skynda dig och kom, ty filistéerna hava fallit in i landet.»
Då upphörde Saul att förfölja David och drog mot filistéerna.
Därav fick det stället namnet Sela-Hammalekot.
Men David drog upp därifrån och uppehöll sig sedan på En-Gedis bergfästen.
Och när Saul kom tillbaka från tåget mot filistéerna, omtalade man för honom att David var i En-Gedis öken.
Då tog Saul tre tusen män, utvalda ur hela Israel, och drog åstad för att söka efter David och hans män på Stenbocksklipporna.
Och när han kom till boskapsgårdarna vid vägen, fanns där en grotta; då gick han ditin för något avsides bestyr.
Men David och hans män sutto längst inne i grottan.
Då sade Davids män till honom: »Se, detta är den dag om vilken HERREN har sagt till dig: Jag vill nu giva din fiende i din hand, så att du far göra med honom vad du finner för gott.»
Då stod David upp och skar oförmärkt av en flik på Sauls mantel.
Men därefter slog Davids samvete honom, därför att han hade skurit av fliken på Sauls mantel.
Och han sade till sina män: »HERREN låte det vara fjärran ifrån mig att jag skulle göra detta mot min herre, mot HERRENS smorde, att jag skulle uträcka min hand mot honom; han är ju HERRENS Smorde.»
Och David höll sina män tillbaka med stränga ord och tillstadde dem icke att överfalla Saul.
Men när Saul hade stått upp och gått ut ur grottan och fortsatt sin färd,
då stod ock David upp och gick ut ur grottan och ropade efter Saul: »Min herre konung!»
När då Saul såg sig tillbaka, böjde David sig ned, med ansiktet mot jorden, och bugade sig.
Och David sade till Saul: »Varför hör du på sådana människors ord, som säga att David söker din ofärd?
Du har ju i dag med egna ögon sett hurusom jag skonade dig, när HERREN i dag hade givit dig i min hand i grottan Och man uppmanade mig att dräpa dig; jag tänkte: 'Jag vill icke uträcka min hand mot min herre; han är ju HERRENS Smorde.
Se själv, min fader, ja, se här fliken av din mantel i min hand.
Ty därav att jag skar av fliken på din mantel, men icke dräpte dig, må du märka och se att jag icke har velat göra något ont eller begå någon förbrytelse, och att jag icke har försyndat mig mot dig, fastän du traktar efter att taga mitt liv.
HERREN skall döma mellan mig och dig, och HERREN skall hämnas mig på dig, men min hand skall icke röra dig.
Det är såsom det gamla ordspråket säger: 'Från de ogudaktiga kommer vad ogudaktigt är'; därför skall hand icke röra dig.»
Efter vem har Israels konung dragit ut?
Efter vem är det du jagar?
Efter en död hund, efter en enda liten loppa!
Så vare då HERREN domare och döme mellan mig och dig; må han se härtill och utföra min sak, ja, må han döma mig fri ifrån din hand.»
När David hade talat dessa ord till Saul, sade Saul: »De är ju din röst, min son David.»
Och Saul brast ut i gråt.
Och han sade till David: »Du är rättfärdigare än jag, ty du har bevisat mig gott, under det jag har bevisat dig ont.
Du har i dag låtit mig se din godhet mot mig, därigenom att du icke har dräpt mig, fastän HERREN hade överlämnat mig i din hand.
Ty när någon träffar på sin fiende, plägar han då låta honom gå sin väg i ro?
HERREN vedergälle dig med sitt goda för vad du denna dag har gjort mig.
Och nu vet jag väl att du skall bliva konung, och att Israels konungadöme skall förbliva i din hand.
Men lova mig nu med ed vid HERREN att du icke utrotar mina avkomlingar efter mig och icke utplånar mitt namn ur min faders hus.»
Då svor David Saul denna ed.
Därefter drog Saul hem; men David och hans män drogo upp till borgen.
Och Samuel dog, och hela Israel församlade sig och höll dödsklagan efter honom; och de begrovo honom där han bodde i Rama.
Och David stod upp och drog ned till öknen Paran.
I Maon fanns då en man som hade sin boskapsskötsel i Karmel, och den mannen var mycket rik; han ägde tre tusen får och ett tusen getter.
Och han höll just då på att klippa sina får i Karmel.
Mannen hette Nabal, och hans hustru hette Abigail.
Hustrun hade ett gott förstånd och ett skönt utseende; men mannen var hård och ondskefull; och han var en avkomling av Kaleb.
När nu David i öknen fick höra att Nabal klippte sina får,
sände han dit tio unga män; och David sade till männen: »Gån upp till Karmel och begiven eder till Nabal och hälsen honom från mig.
Och I skolen säga till mina bröder där: »Frid vare med dig själv frid vare med ditt hus, och frid vare med allt vad du har.
Jag har nu hört att du håller på med fårklippning.
Nu är det så att dina herdar hava vistats i vårt grannskap, utan att vi hava gjort dem något förfång, och utan att något har kommit bort för dem under hela den tid de hava varit i Karmel.
Fråga dina tjänare därom, så skola de själva säga dig det.
Låt nu våra män finna nåd för dina ögon.
Vi hava ju kommit hit på en glad dag.
Giv därför åt dina tjänare och åt din son David vad du kan hava till hands.»
När nu Davids män kommo dit, talade de på Davids vägnar till Nabal alldeles såsom det var dem befallt, och sedan väntade de stilla.
Men Nabal svarade Davids tjänare och sade: »Vem är David, vem är Isais son?
I denna tid är det många tjänare som rymma från sina herrar.
Skulle jag taga min mat och min dryck och slaktdjuren, som jag har slaktat åt mina fårklippare, och giva detta åt män om vilka jag icke ens vet varifrån de äro?»
Då vände Davids män om och gingo sin väg; och när de hade kommit tillbaka, berättade de for honom allt, såsom det hade tillgått.
Då sade David till sina män: »Var och en omgjorde sig med sitt svärd.»
Och var och en omgjordade sig med sitt svärd; jämväl David själv omgjordade sig med sitt svärd.
Och vid pass fyra hundra man följde med David ditupp, men två hundra stannade vid trossen.
Men en av tjänarna berättade för Abigail, Nabals hustru, och sade: »David har skickat sändebud hit från öknen och låtit hälsa vår herre, men han visade av dem.
Dessa män hava likväl varit oss mycket nyttiga; vi hava aldrig lidit något förfång, och aldrig har något kommit bort för oss under hela den tid vi drogo omkring i deras närhet, medan vi voro därute på marken.
De voro en mur för oss både dag och natt under hela den tid vi vistades i deras grannskap, medan vi vaktade hjorden.
Så betänk nu och se till, vad du bör göra, ty något ont är nog beslutet mot vår herre och över hela hans hus; och han är ju en ond man, så att ingen vågar säga något åt honom.»
Då gick Abigail strax och tog två hundra bröd, två vinläglar, fem tillredda får, fem sea-mått rostade ax, ett hundra russinkakor och två hundra fikonkakor, och lastade detta på åsnor.
Och hon sade till sina tjänare: »Gån framför mig, jag vill komma efter eder.»
Men för sin man Nabal sade hon intet härom.
När hon nu red på sin åsna och kom ned i en hålväg i berget, fick hon se David och hans män komma ned från motsatta sidan, så att hon måste möta dem.
Men David hade sagt: »Förgäves har jag skyddat allt vad den mannen hade i öknen, så att intet av allt vad han ägde har kommit bort; men har har vedergällt mig med ont för gott.
Så sant Gud må straffa Davids fiender nu och framgent, jag skall av allt som tillhör honom icke låta någon av mankön leva kvar till i morgon.»
Då nu Abigail fick se David, steg hon strax ned från åsnan och föll ned inför David på sitt ansikte och bugade sig mot jorden.
Hon föll till hans fötter och sade: »På mig vilar denna missgärning, herre.
Men låt din tjänarinna få tala inför dig, och hör på din tjänarinnas ord.
Icke må min herre fästa något avseende vid Nabal, den onde mannen, ty vad hans namn betyder, det är han; Nabal heter han, och dårskap bor i honom.
Men jag, din tjänarinna, har icke sett de män som du, min herre, sände.
Och nu, min herre, så sant HERREN lever, och så sant du själv lever, du som av HERREN har avhållits från att ådraga dig blodskuld och skaffa dig rätt med egen hand: må det nu gå dina fiender och dem som söka bereda min herre ofärd såsom det må gå Nabal.
Och låt nu dessa hälsningsskänker, som din trälinna har medfört till min herre, givas åt de män som följa min herre.
Förlåt din tjänarinna vad hon har brutit.
Ty HERREN skall förvisso åt min herre uppbygga ett hus som bliver beståndande, eftersom min herre för HERRENS krig; och du skall icke bliva skyldig till något ont, så länge du lever.
Och om någon står upp för att förfölja dig och söka döda dig, så må min herres liv vara inknutet i de levandes pung hos HERREN, din Gud; men dina fienders liv må han lägga i sin slunga och slunga det bort.
När nu HERREN gör med min herre allt det goda varom han har talat till dig, och förordnar dig till furste över Israel,
skall alltså detta icke bliva dig en stötesten eller vara till hjärteångest för min herre, att du har utgjutit blod utan sak, och att min herre själv har skaffat sig rätt.
Men när HERREN gör min herre gott, så tänk på din tjänarinna.»
Då sade David till Abigal: »Välsignad vare HERREN, Israels Gud som i dag har sänt dig mig till mötes!
Och välsignat vare ditt förstånd, och välsignad vare du själv, som i dag har hindrat mig från att ådraga mig blodskuld och skaffa mig rätt med egen hand!
Men så sant HERREN, Israels Gud, lever, han som har avhållit mig från att göra dig något ont: om du icke strax hade kommit mig till mötes, så skulle i morgon, när det hade blivit dager, ingen av mankön hava funnits kvar av Nabals hus.»
Därefter tog David emot av henne vad hon hade medfört åt honom; och han sade till henne: »Far i frid hem igen.
Se, jag har lyssnat till dina ord och gjort dig till viljes.»
När sedan Abigail kom hem till Nabal, höll denne just i sitt hus ett gästabud, som var såsom en konungs gästabud; och Nabals hjärta var glatt i honom, och han var mycket drucken.
Därför omtalade hon alls intet för honom förrän om morgonen, när det blev dager.
Men om morgonen, när ruset hade gått av Nabal, omtalade hans hustru för honom vad som hade hänt.
Då blev hans hjärta såsom dött i hans bröst, och han blev såsom en sten.
Och vid pass tio dagar därefter slog HERREN Nabal, så att han dog.
När David hörde att Nabal var död, sade han: »Lovad vare HERREN, som på Nabal har hämnats den smälek han tillfogade mig, och som har bevarat sin tjänare från att göra vad ont var, under det att HERREN lät Nabals ondska komma tillbaka över hans eget huvud!»
Och David sände åstad och lät säga Abigail att han önskade få henne till sin hustru.
När så Davids tjänare kommo till Abigail i Karmel, talade de till henne och sade: »David har sänt oss till dig för att få dig till hustru åt sig.»
Då stod hon upp och föll ned till jorden på sitt ansikte och sade: »Må din tjänarinna bliva en trälinna, som tvår min herres tjänares fötter.»
Därefter stod Abigail upp med hast och satte sig på sin åsna, likaledes de fem tärnor som utgjorde hennes följe.
Och hon följde med dem som David hade sänt till henne och blev hans hustru.
David hade ock tagit till hustru Ahinoam från Jisreel, så att dessa båda blevo hans hustrur.
Men Saul hade givit sin dotter Mikal, Davids hustru, åt Palti, Lais' son, från Gallim.
Och sifiterna kommo till Saul i Gibea och sade: »David håller sig nu gömd på Hakilahöjden, gent emot ödemarken.»
Då bröt Saul upp och drog ned till öknen Sif med tre tusen män utvalda ur Israel, för att söka efter David i öknen Sif.
Och Saul lägrade sig på Hakilahöjden, som ligger gent emot ödemarken, vid vägen.
Men David uppehöll sig då i öknen.
Och när David förnam att Saul hade kommit efter honom in i öknen,
sände han ut spejare och fick så full visshet om att Saul hade kommit.
Då bröt David upp och begav sig till det ställe där Saul hade lägrat sig; och David såg platsen där Saul låg med sin härhövitsman Abner, Ners son.
Saul låg nämligen i vagnborgen, och folket var lägrat runt
Och David tog till orda och sade I till hetiten Ahimelek och till Abisai, Serujas son, Joabs broder: »Vem vill gå med mig ned till Saul i lägret?»
Då svarade Abisai: »Jag vill gå med dig ditned.»
Så kommo då David och Abisai om natten till folket där, och sågo Saul ligga och sova i vagnborgen, med spjutet nedstött i jorden invid huvudgärden; och Abner och folket lågo runt omkring honom.
Då sade Abisai till David: »Gud har i dag överlämnat din fiende i din hand; så låt mig nu få spetsa honom fast i jorden med spjutet; det skall ske genom en enda stöt, jag skall icke behöva giva honom mer än den.»
Men David svarade Abisai: »Du får icke förgöra honom; ty vem har uträckt sin hand mot HERRENS smorde och förblivit ostraffad?»
Och David sade ytterligare: »Så sant HERREN lever, HERREN må själv slå honom, eller ock må hans dödsdag komma i vanlig ordning, eller må han draga ut i strid och så få sin bane;
men HERREN låte det vara fjärran ifrån mig att jag skulle uträcka min hand mot HERRENS smorde.
Tag nu likväl spjutet som står vid hans huvudgärd och vattenkruset; och låt oss sedan gå vår väg.
Och David tog spjutet och vattenkruset från Sauls huvudgärd, och sedan gingo de sin väg.
Men ingen såg eller märkte det eller ens vaknade, utan allasammans sovo; ty HERREN hade låtit en tung sömn falla över dem.
Sedan, när David hade kommit över på andra sidan, ställde han sig på toppen av berget, långt ifrån så att avståndet var stort mellan dem.
Och David ropade till folket och till Abner, Ners son, och sade: »Vill du icke svara, Abner?»
Abner svarade och sade: »Vem är du som så ropar till konungen?»
David sade till Abner: »Du är ju en man som icke har sin like i Israel.
Varför har du då icke vakat över din herre, konungen?
En av folket har ju kommit in för att förgöra konungen, din herre.
Vad du har gjort är icke väl gjort.
Så sant HERREN lever, I haden förtjänat att dö, därför att I icke haven vakat över eder herre, HERRENS smorde.
Se nu efter: var äro konungens spjut och vattenkruset som stodo vid hans huvudgärd?»
Då kände Saul igen Davids röst och sade: »Det är ju din röst, min son David.»
David svarade: »Ja, min herre konung.»
Och han sade ytterligare: »Varför jagar min herre så efter sin tjänare?
Vad har jag då gjort, och vad för ont är i min hand?
Må nu min herre konungen höra sin tjänares ord: Om det är HERREN som har uppeggat dig emot mig, så låt honom få känna lukten av en offergåva; men om det är människor, så vare de förbannade inför HERREN, därför att de nu hava drivit mig bort, så att jag icke får uppehålla mig i HERRENS arvedel.
De säga ju: 'Gå bort och tjäna andra gudar.'
Och må nu icke mitt blod falla på jorden fjärran ifrån HERRENS ansikte, då Israels konung har dragit ut för att söka efter en enda liten loppa, såsom man jagar rapphöns på bergen.»
Då sade Saul: »Jag har syndat.
Kom tillbaka, min son David; ty jag vill icke mer göra dig något ont, eftersom mitt liv i dag har varit dyrt aktat i dina ögon.
Se, ja har handlat i mycket stor dårskap och förvillelse.»
David svarade och sade: »Se här är spjutet, o konung; låt nu en av dina män komma hitöver och hämta det.
Och HERREN skall vedergälla var och en för hans rättfärdighet och trofasthet.
HERREN gav dig ju dag i min hand, men jag ville icke uträcka min hand mot HERRENS smorde.
Och likasom ditt liv i dag har varit högt aktat i mina ögon, så så ock mitt liv vara högt aktat i HERRENS ögon, så att han räddar mig ur all nöd.»
Saul sade till David: »Välsignad vare du, min son David!
Vad du företager dig, det skall du ock förmå utföra.»
Därefter gick David sin väg, och Saul vände tillbaka hem igen.
Men David sade till sig själv: »En dag skall jag nu i alla fall omkomma genom Sauls hand.
Ingen annan räddning finnes för mig än att fly undan till filistéernas land; då måste Saul avstå ifrån att vidare söka efter mig över hela Israels område, och så undkommer jag hans hand.»
Och David bröt upp och drog med sina sex hundra man över till Akis, Maoks son, konungen i Gat.
Och David stannade hos Akis i Gat med sina män, var och en med sitt husfolk, David med sina båda hustrur, Ahinoam från Jisreel och Abigail, karmeliten Nabals hustru.
Och när det blev berättat för Saul att David hade flytt till Gat, sökte han icke vidare efter honom.
Men David sade till Akis: »Om jag har funnit nåd för dina ögon, så låt mig få min bostad i någon av landsortsstäderna, så att jag får vistas där.
Varför skulle din tjänare bo i huvudstaden hos dig?»
Då gav Akis honom samma dag Siklag.
Därför hör Siklag ännu i dag under Juda konungar.
Den tid David bodde i filistéernas land var sammanräknat ett år och fyra månader.
Men David drog upp med sina män, och de företogo plundringståg i gesuréernas, girsiternas och amalekiternas land.
Ty dessa stammar bodde sedan gammalt där i landet, fram emot Sur och ända intill Egyptens land.
Och så ofta David härjade i landet, lät han varken män eller kvinnor bliva vid liv; men får och fäkreatur och åsnor och kameler och kläder tog han med sig och vände så tillbaka och kom till Akis.
När då Akis sade: »Haven I väl i dag företagit något plundringståg?», svarade David: »Ja, i den del av Sydlandet, som tillhör Juda», eller: »I den del av Sydlandet, som tillhör jerameeliterna», eller: »I den del av Sydlandet, som tillhör kainéerna.»
Men att David lät varken män eller kvinnor bliva vid liv och komma till Gat, det skedde därför att han tänkte: »De kunde eljest förråda oss och säga: 'Så och så har David gjort, så har han betett sig under hela den tid han har bott i filistéernas land.'»
Därför trodde Akis David och tänkte: »Han har nu gjort sig förhatlig för sitt folk Israel och kommer att bliva min tjänare för alltid.
Vid den tiden församlade filistéerna sina krigshärar för att strida mot Israel.
Och Akis sade till David: »Du må veta att du med dina män nu måste draga ut med mig i härnad.»
David svarade Akis: »Välan, då skall du ock få märka vad din tjänare kan uträtta.»
Akis sade till David »Välan, jag sätter dig alltså till väktare över mitt huvud för beständigt.»
Samuel var nu död, och hela Israel hade hållit dödsklagan efter honom; och de hade begravit honom i hans stad, i Rama.
Och Saul hade utdrivit andebesvärjare och spåmän ur landet.
Så församlade sig nu filistéerna och kommo och lägrade sig vid Sunem.
Då församlade ock Saul hela Israel, och de lägrade sig vid Gilboa.
Men när Saul såg filistéernas läger, fruktade han och förskräcktes högeligen i sitt hjärta.
Och Saul frågade HERREN, men HERREN svarade honom icke, varken genom drömmar eller genom urim eller genom profeter.
Då sade Saul till sina tjänare: »Söken upp åt mig någon andebesvärjerska, så vill jag gå till henne och fråga henne.»
Hans tjänare svarade honom: »I En-Dor finnes en andebesvärjerska.»
Då gjorde Saul sig oigenkännlig och tog på sig andra kläder och gick åstad med två män; och de kommo till kvinnan om natten.
Och han sade: »Spå åt mig genom anden, och mana upp åt mig den jag säger dig.»
Men kvinnan svarade honom: »Du vet ju själv vad Saul har gjort, huru han har utrotat andebesvärjare och spåmän ur landet.
Varför lägger du då ut en snara för mitt liv och vill döda mig?»
Då svor Saul henne en ed vid HERREN och sade: »Så sant HERREN lever, i denna sak skall intet tillräknas dig såsom missgärning.»
Kvinnan frågade: »Vem skall jag då mana upp åt dig?»
Han svarade: »Mana upp Samuel åt mig.»
Men när kvinnan fick se Samuel, gav hon till ett högt rop.
Och kvinnan sade till Saul: »Varför har du bedragit mig?
Du är ju Saul.»
Konungen sade till henne: »Frukta icke.
Vad är det då du ser?»
Kvinnan svarade Saul: »Jag ser ett gudaväsen komma upp ur jorden.»
Han frågade henne: »Huru ser han ut?»
Hon svarade: »Det är en gammal man som kommer upp, höljd i en kåpa.»
Då förstod Saul att det var Samuel, och böjde sig ned med ansiktet mot jorden och bugade sig.
Och Samuel sade till Saul: »Varför har du stört min ro och manat mig upp?»
Saul svarade: »Jag är i stor nöd: filistéerna hava begynt krig mot mig, och Gud har vikit ifrån mig och svarar mig icke mer, varken genom profeter eller genom drömmar.
Därför har jag kallat dig upp, på det att du må låta mig veta vad jag skall göra.»
Men Samuel svarade: »Varför frågar du mig, då nu HERREN har vikit ifrån dig och blivit din fiende?
HERREN har efter sitt behag gjort vad han hade sagt genom mig: HERREN har ryckt riket ur din hand och givit det åt en annan, åt David.
Eftersom du icke hörde HERRENS röst och icke lät Amalek känna hans vredes glöd, därför har HERREN nu gjort dig detta.
HERREN skall giva både dig och Israel i filistéernas hand, och i morgon skall du med dina söner vara hos mig; ja, också Israels läger skall HERREN giva i filistéernas hand.»
Då föll Saul strax raklång till jorden; så förfärad blev han över Samuels ord.
Också voro hans krafter uttömda, ty på ett helt dygn hade han ingenting ätit.
Men kvinnan gick fram till Saul, och när hon såg huru högeligen förskräckt han var, sade hon till honom: »Se, din tjänarinna lyssnade till din begäran; Jag tog min själ i min hand och hörsammade den önskan du uttalade till mig.
Så lyssna nu också du till dina tjänarinnas ord och låt mig sätta fram litet mat för dig, och ät, så att du hämtar krafter, innan du går dina färde.»
Men han vägrade och sade: »Jag vill icke äta.»
Då bådo honom hans tjänare jämte kvinnan så enträget, att han lyssnade till deras ord; han stod upp från jorden och satte sig på vilobädden.
Och kvinnan hade en gödd kalv i huset; den slaktade hon nu i hast.
Därpå tog hon mjöl och knådade det och bakade därav osyrat bröd.
Sedan satte hon fram det för Saul: och hans tjänare, och de åto.
Därefter stodo de upp och gingo samma natt sina färde.
Filistéerna församlade nu alla sina härar i Afek, medan israeliterna voro lägrade vid källan i Jisreel.
Då nu filistéernas hövdingar tågade fram med avdelningar på hundra och tusen, och David och hans män därvid tågade sist fram, tillika med Akis,
sade filistéernas furstar: »Vad hava dessa hebréer här att göra?»
Men Akis svarade filistéernas furstar: »Denne David är ju Sauls, Israels konungs, tjänare, som nu har varit hos mig över år och dag, och jag har icke funnit något ont hos honom, från den dag han gick över till mig ända till denna dag.
Då blevo filistéernas furstar förtörnade på honom; och filistéernas furstar sade till honom: »Låt mannen vända om och gå tillbaka till den ort du har anvisat honom; han får icke draga med med oss till strid, för att han icke under striden må bliva vår motståndare.
Ty varigenom skulle han väl bättre kunna göra sig behaglig för sin herre än genom dessa mäns huvuden?
Han är ju den David till vilkens ära man sjunger så under dansen: 'Saul har slagit sina tusen, men David sina tio tusen.'»
Då kallade Akis David till sig och sade till honom: »Så sant HERREN lever, du är en redlig man, och att du går ut och in här hos mig i lägret är mig välbehagligt, ty jag har icke funnit något ont hos dig, från den dag du kom till mig ända till denna dag; men för hövdingarna är du icke välbehaglig.
Så vänd nu tillbaka och gå i frid, för att du icke må göra något som misshagar filistéernas hövdingar.»
David sade till Akis: »Vad har jag då gjort, och vad har du funnit hos din tjänare, från den dag jag kom i din tjänst ända till denna dag, eftersom jag icke får gå åstad och strida mot min herre konungens fiender?»
Akis svarade och sade till David: »Jag vet bäst att du är mig välbehaglig såsom en Guds ängel; men filistéernas furstar säga: 'Han får icke draga upp med oss i striden.'
Så stå nu upp bittida i morgon, jämte din herres tjänare som hava kommit hit med dig; och när morgon haven stått bittida upp, mån I draga edra färde, så snart det har blivit dager.»
Då stod David bittida upp med sina män för att om morgonen drag tillbaka till filistéernas land.
Men filistéerna drogo upp till Jisreel.
När David med sina män på tredje dagen kom till Siklag, hade amalekiterna infallit i Sydlandet och i Siklag; och de hade intagit Siklag och bränt upp det i eld.
Och kvinnorna som voro därinne, både små och stora, hade de fört bort såsom fångar, utan att döda någon; de hade allenast fört bort dem och gått sin väg.
När nu David med sina män kom till staden och fick se att den var uppbränd i eld, och att deras hustrur jämte deras söner och döttrar voro bortförda såsom fångar,
brast han ut i gråt, så ock hans folk; och de gräto, till dess att de icke förmådde gråta mer.
Davids båda hustrur, Ahinoam från Jisreel och Abigail, karmeliten Nabals hustru, voro också fångna.
Och David kom i stor nöd, ty folket tänkte stena honom; så förbittrat var allt folket, var och en för sina söners och döttrars skull.
Men David hämtade styrka hos HERREN, sin Gud.
Och David sade till prästen Ebjatar, Ahimeleks son: »Bär hit till mig efoden.»
Då bar Ebjatar fram efoden till David.
David frågade nu HERREN: »Skall jag sätta efter denna rövarskara?
Kan jag då hinna upp den?»
Han svarade honom: »Sätt efter dem; ty du skall förvisso hinna upp dem och skaffa räddning.»
Då begav sig David åstad med sina sex hundra man, och de kommo till bäcken Besor; där stannade de som nödgades bliva efter.
Men David fortsatte förföljelsen med fyra hundra man; ty de som sade blivit för trötta, och som därför stannade, utan att gå över bäcken Besor, utgjorde två hundra man.