Ty jag säger eder: Härefter skolen I icke få se mig, intill den tid då I sägen: 'Välsignad vare han som kommer, i Herrens namn.'»
Och Jesus gick därifrån, ut ur helgedomen.
Hans lärjungar trädde då fram och bådo honom giva akt på helgedomens byggnader.
Då svarade han och sade till dem: »Ja, I sen nu allt detta; men sannerligen säger jag eder: Här skall icke lämnas sten på sten; allt skall bliva nedbrutet.»
När han sedan satt på Oljeberget, trädde hans lärjungar fram till honom, medan de voro allena, och sade: »Säg oss när detta skall ske, och vad som bliver tecknet till din tillkommelse och tidens ände.»
Då svarade Jesus och sade till dem: »Sen till, att ingen förvillar eder.
Ty många skola komma under mitt namn och säga: 'Jag är Messias' och skola förvilla många.
Och I skolen få höra krigslarm och rykten om krig; sen då till, att I icke förloren besinningen, ty sådant måste komma, men därmed är ännu icke änden inne.
Ja, folk skall resa sig upp mot folk och rike mot rike, och det skall bliva hungersnöd och jordbävningar på den ena orten efter den andra;
men allt detta är allenast begynnelsen till 'födslovåndorna'.
Då skall man prisgiva eder till misshandling, och man skall dräpa eder, och I skolen bliva hatade av alla folk, för mitt namns skull.
Och då skola många komma på fall, och den ene skall förråda den andre, och den ene skall hata den andre.
Och många falska profeter skola uppstå och skola förvilla många.
Och därigenom att laglösheten förökas, skall kärleken hos de flesta kallna.
Men den som är ståndaktig intill änden, han skall bliva frälst.
Och detta evangelium om riket skall bliva predikat i hela världen, till ett vittnesbörd för alla folk.
Och sedan skall änden komma.
När I nu fån se 'förödelsens styggelse', om vilken är talat genom profeten Daniel, stå på helig plats -- den som läser detta, han give akt därpå --
då må de som äro i Judeen fly bort till bergen,
och den som är på taket må icke stiga ned för att hämta vad som finnes i hans hus,
och den som är ute på marken må icke vända tillbaka för att hämta sin mantel.
Och ve dem som äro havande, eller som giva di på den tiden!
Men bedjen att eder flykt icke må ske om vintern eller på sabbaten.
Ty då skall det bliva 'en stor vedermöda, vars like icke har förekommit allt ifrån världens begynnelse intill nu', ej heller någonsin skall förekomma.
Och om den tiden icke bleve förkortad, så skulle intet kött bliva frälst; men för de utvaldas skull skall den tiden bliva förkortad.
Om någon då säger till eder: 'Se här är Messias', eller: 'Där är han', så tron det icke.
Ty människor som falskeligen säga sig vara Messias skola uppstå, så ock falska profeter, och de skola göra stora tecken och under, för att, om möjligt förvilla jämväl de utvalda.
Jag har nu sagt eder det förut.
Därför, om man säger till eder: 'Se, han är i öknen', så gån icke ditut, eller: 'Se, han är inne i huset', så tron det icke.
Ty såsom ljungelden, när den går ut från öster, synes ända till väster, så skall Människosonens tillkommelse vara. --
Där åteln är, dit skola rovfåglarna församla sig.
Men strax efter den tidens vedermöda skall solen förmörkas och månen upphöra att giva sitt sken, och stjärnorna skola falla ifrån himmelen, och himmelens makter skola bäva.
Och då skall Människosonens tecken visa sig på himmelen, och alla släkter på jorden skola då jämra sig.
Och man skall få se 'Människosonen komma på himmelens skyar' med stor makt och härlighet.
Och han skall sända ut sina änglar med starkt basunljud, och de skola församla hans utvalda från de fyra väderstrecken, från himmelens ena ända till den andra.
Ifrån fikonträdet mån I här hämta en liknelse.
När dess kvistar begynna att få save och löven spricka ut, då veten I att sommaren är nära.
Likaså, när I sen allt detta, då kunnen I ock veta att han är nära och står för dörren.
Sannerligen säger jag eder: Detta släkte skall icke förgås, förrän allt detta sker.
Himmel och jord skola förgås, men mina ord skola aldrig förgås.
Men om den dagen och den stunden vet ingen något, icke ens änglarna i himmelen, ingen utom Fadern allena.
Ty såsom det skedde på Noas tid, så skall det ske vid Människosonens tillkommelse.
Såsom människorna levde på den tiden, före floden: de åto och drucko, män togo sig hustrur, och hustrur gåvos åt män, ända till den dag då Noa gick in i arken;
och de visste av intet, förrän floden kom och tog dem allasammans bort -- så skall det ske vid Människosonens tillkommelse.
Då skola två män vara tillsammans ute på marken; en skall bliva upptagen, och en skall lämnas kvar.
Två kvinnor skola mala på samma kvarn; en skall bliva upptagen, och en skall lämnas kvar.
Vaken fördenskull; ty I veten icke vilken dag vår Herre kommer.
Men det förstån I väl, att om husbonden visste under vilken nattväkt tjuven skulle komma, så vakade han och tillstadde icke att någon bröt sig in i hans hus.
Varen därför ock I redo; ty i en stund då I icke vänten det skall Människosonen komma.
Finnes nu någon trogen och förståndig tjänare, som av sin herre har blivit satt över hans husfolk för att giva dem mat i rätt tid --
salig är då den tjänaren, om hans herre, när han kommer, finner honom göra så.
Sannerligen säger jag eder: Han skall sätta honom över allt vad han äger.
Men om så är, att tjänaren är en ond man, som säger i sitt hjärta: 'Min herre kommer icke så snart',
och han begynner slå sina medtjänare och äter och dricker med dem som äro druckna,
då skall den tjänarens herre komma på en dag då han icke väntar det, och i en stund då han icke tänker sig det,
och han skall låta hugga honom i stycken och låta honom få sin del med skrymtare.
Där skall vara gråt och tandagnisslan.»
»Då skall det vara med himmelriket, såsom när tio jungfrur togo sina lampor och gingo ut för att möta brudgummen.
Men fem av dem voro oförståndiga, och fem voro förståndiga.
De oförståndiga togo väl sina lampor, men togo ingen olja med sig.
De förståndiga åter togo olja i sina kärl, tillika med lamporna.
Då nu brudgummen dröjde, blevo de alla sömniga och somnade.
Men vid midnattstiden ljöd ett anskri: 'Se brudgummen kommer!
Gån ut och möten honom.'
Då stodo alla jungfrurna upp och redde till sina lampor.
Och de oförståndiga sade till de förståndiga: 'Given oss av eder olja, ty våra lampor slockna.'
Men de förståndiga svarade och sade: 'Nej, den skulle ingalunda räcka till för både oss och eder.
Gån hellre bort till dem som sälja, och köpen åt eder.'
Men när de gingo bort för att köpa, kom brudgummen, och de som voro redo gingo in med honom till bröllopet, och dörren stängdes igen.
Omsider kommo ock de andra jungfrurna och sade: 'Herre, herre, låt upp för oss.'
Men han svarade och sade: 'Sannerligen säger jag eder: Jag känner eder icke.'
Vaken fördenskull; ty I veten icke dagen, ej heller stunden.
Ty det skall ske, likasom när en man som ville fara utrikes kallade till sig sina tjänare och överlämnade åt dem sina ägodelar;
åt en gav han fem pund, åt en annan två och åt en tredje ett pund, åt var och en efter hans förmåga, och for utrikes.
Strax gick då den som hade fått de fem punden bort och förvaltade dem så, att han med dem vann andra fem pund.
Den som hade fått de två punden vann på samma sätt andra två.
Men den som hade fått ett pund gick bort och grävde en grop i jorden och gömde där sin herres penningar.
En lång tid därefter kom tjänarnas herre hem och höll räkenskap med dem.
Då trädde den fram, som hade fått de fem punden, och bar fram andra fem pund och sade: 'Herre, du överlämnade åt mig fem pund; se, andra fem pund har jag vunnit.'
Hans herre svarade honom: 'Rätt så, du gode och trogne tjänare!
När du var satt över det som ringa är, var du trogen; jag skall sätta dig över mycket.
Gå in i din herres glädje.'
Så trädde ock den fram, som hade fått de två punden, och sade: 'Herre, du överlämnade åt mig två pund; se, andra två pund har jag vunnit.'
Hans herre svarade honom: 'Rätt så, du gode och trogne tjänare!
När du var satt över det som ringa är, var du trogen; jag skall sätta dig över mycket.
Gå in i din herres glädje.'
Sedan trädde ock den fram, som hade fått ett pund, och sade: 'Herre, jag hade lärt känna dig såsom en sträng man, som vill skörda, där du icke har sått, och inbärga, där du icke har utstrött;
och av fruktan för dig gick jag bort och gömde ditt pund i jorden.
Se här har du vad dig tillhör.'
Då svarade hans herre och sade till honom: 'Du onde och late tjänare, du visste att jag vill skörda, där jag icke har sått, och inbärga, där jag icke har utstrött?
Då borde du också hava satt in mina penningar i en bank, så att jag hade fått igen mitt med ränta, när jag kom hem.
Tagen därför ifrån honom hans pund, och given det åt den som har de tio punden.
Ty var och en som har, åt honom skall varda givet, så att han får över nog; men den som icke har, från honom skall tagas också det han har.
Och kasten den oduglige tjänaren ut i mörkret härutanför.'
Där skall vara gråt och tandagnisslan.
Men när Människosonen kommer i sin härlighet, och alla änglar med honom, då skall han sätta sig på sin härlighets tron.
Och inför honom skola församlas alla folk och han skall skilja dem från varandra, såsom en herde skiljer fåren ifrån getterna.
Och fåren skall han ställa på sin högra sida, och getterna på den vänstra.
Därefter skall Konungen säga till dem som stå på hans högra sida: 'Kommen, I min Faders välsignade, och tagen i besittning det rike som är tillrett åt eder från världens begynnelse.
Ty jag var hungrig, och I gåven mig att äta; jag var törstig, och I gåven mig att dricka; jag var husvill, och I gåven mig härbärge,
naken, och I klädden mig; jag var sjuk, och I besökten mig; jag var i fängelse, och I kommen till mig.'
Då skola de rättfärdiga svara honom och säga: 'Herre, när sågo vi dig hungrig och gåvo dig mat, eller törstig och gåvo dig att dricka?
Och när sågo vi dig husvill och gåvo dig härbärge, eller naken och klädde dig?
Och när sågo vi dig sjuk eller i fängelse och kommo till dig?'
Då skall Konungen svara och säga till dem: 'Sannerligen säger jag eder: Vadhelst I haven gjort mot en av dessa mina minsta bröder, det haven I gjort mot mig.'
Därefter skall han ock säga till dem som stå på hans vänstra sida: 'Gån bort ifrån mig, I förbannade, till den eviga elden, som är tillredd åt djävulen och hans änglar.
Ty jag var hungrig, och I gåven mig icke att äta; jag var törstig, och I gåven mig icke att dricka;
jag var husvill, och I gåven mig icke härbärge, naken, och I klädden mig icke, sjuk och i fängelse, och I besökten mig icke.'
Då skola också de svara och säga: 'Herre, när sågo vi dig hungrig eller törstig eller husvill eller naken eller sjuk eller i fängelse och tjänade dig icke?'
Då skall han svara dem och säga: 'Sannerligen säger jag eder: Vadhelst I icke haven gjort mot en av dessa minsta, det haven I ej heller gjort mot mig.'
Och dessa skola då då bort till evigt straff, men de rättfärdiga till evigt liv.»
När nu Jesus hade talat allt detta till slut, sade han till sina lärjungar:
»I veten att det två dagar härefter är påsk; då skall Människosonen bliva förrådd och utlämnad till att korsfästas.»
Därefter församlade sig översteprästerna och folkets äldste hos översteprästen, som hette Kaifas, i hans hus,
och rådslogo om att låta gripa Jesus med list och döda honom.
Men de sade: »Icke under högtiden, för att ej oroligheter skola uppstå bland folket.»
Men när Jesus var i Betania, i Simon den spetälskes hus,
framträdde till honom en kvinna som hade med sig en alabasterflaska med dyrbar smörjelse; denna göt hon ut över hans huvud, där han låg till bords.
Då lärjungarna sågo detta, blevo de misslynta och sade: »Varför skulle detta förspillas?
Man hade ju kunnat sälja det för mycket penningar och giva dessa åt de fattiga.»
När Jesus märkte detta, sade han till dem: »Varför oroen I kvinnan?
Det är en god gärning som hon har gjort mot mig.
De fattiga haven I ju alltid ibland eder, men mig haven I icke alltid.
När hon göt ut denna smörjelse på min kropp, gjorde hon det såsom en tillredelse till min begravning.
Sannerligen säger jag eder: Varhelst i hela världen detta evangelium bliver predikat, där skall ock det som hon nu har gjort bliva omtalat, henne till åminnelse.»
Därefter gick en av de tolv, den som hette Judas Iskariot, bort till översteprästerna
och sade: »Vad viljen I giva mig för att jag skall överlämna honom åt eder?»
Då vägde de upp åt honom trettio silverpenningar.
Och från den stunden sökte han efter lägligt tillfälle att förråda honom.
Men på första dagen i det osyrade brödets högtid trädde lärjungarna fram till Jesus och frågade: »Var vill du att vi skola reda till åt dig att äta påskalammet?»
Han svarade: »Gån in i staden till den och den och sägen till honom: 'Mästaren låter säga: Min tid är nära; hos dig vill jag hålla påskhögtid med mina lärjungar.'»
Och lärjungarna gjorde såsom Jesus hade befallt dem och redde till påskalammet.
När det nu hade blivit afton, lade han sig till bords med de tolv.
Och medan de åto, sade han: »Sannerligen säger jag eder: En av eder skall förråda mig.»
Då blevo de mycket bedrövade och begynte fråga honom, var efter annan: »Icke är det väl jag, Herre?»
Då svarade han och sade: »Den som jämte mig nu doppade handen i fatet, han skall förråda mig.
Människosonen skall gå bort, såsom det är skrivet om honom; men ve den människa genom vilken Människosonen bliver förrådd!
Det hade varit bättre för den människan, om hon icke hade blivit född.»
Judas, han som förrådde honom, tog då till orda och frågade: »Rabbi, icke är det väl jag?»
Han svarade honom: »Du har själv sagt det.»
Medan de nu åto, tog Jesus ett bröd och välsignade det och bröt det och gav åt lärjungarna och sade: »Tagen och äten; detta är min lekamen.»
Och han tog en kalk och tackade Gud och gav åt dem och sade: »Dricken härav alla;
ty detta är mitt blod, förbundsblodet, som varder utgjutet för många till syndernas förlåtelse.
Och jag säger eder: Härefter skall jag icke mer dricka av det som kommer från vinträd, förrän på den dag då jag dricker det nytt med eder i min Faders rike.»
När de sedan hade sjungit lovsången, gingo de ut till Oljeberget.
Då sade Jesus till dem: »I denna natt skolen I alla komma på fall för min skull, ty det är skrivet: 'Jag skall slå herden, och fåren i hjorden skola förskingras.'
Men efter min uppståndelse skall jag före eder gå till Galileen.»
Då svarade Petrus och sade till honom: »Om än alla andra komma på fall för din skull, så skall dock jag aldrig komma på fall.»
Jesus sade till honom: »Sannerligen säger jag dig: I denna natt, förrän hanen har galit, skall du tre gånger förneka mig.»
Petrus svarade honom: »Om jag än måste dö med dig, så skall jag dock förvisso icke förneka dig.»
Sammalunda sade ock alla de andra lärjungarna.
Därefter kom Jesus med dem till ett ställe som hette Getsemane.
Och han sade till lärjungarna: »Bliven kvar här, medan jag går dit bort och beder.»
Och han tog med sig Petrus och Sebedeus' två söner; och han begynte bedrövas och ängslas.
Då sade han till dem: »Min själ är djupt bedrövad, ända till döds; stannen kvar här och vaken med mig.»
Därefter gick han litet längre bort och föll ned på sitt ansikte och bad och sade: »Min Fader, om det är möjligt, så gånge denna kalk ifrån mig.
Dock icke såsom jag vill, utan såsom du vill!»
Sedan kom han tillbaka till lärjungarna och fann dem sovande.
Då sade han till Petrus: »Så litet förmådden I då vaka en kort stund med mig!
Vaken, och bedjen att I icke mån komma i frestelse.
Anden är villig, men köttet är svagt.»
Åter gick han bort, för andra gången, och bad och sade: »Min Fader, om detta icke kan gå ifrån mig, utan jag måste dricka denna kalk, så ske din vilja.»
När han sedan kom tillbaka, fann han dem åter sovande, ty deras ögon voro förtyngda.
Då lät han dem vara och gick åter bort och bad, för tredje gången, och sade återigen samma ord.
Därefter kom han tillbaka till lärjungarna och sade till dem: »Ja, I soven ännu alltjämt och vilen eder!
Se, stunden är nära då Människosonen skall bliva överlämnad i syndares händer.
Stån upp, låt oss gå; se, den är nära, som förråder mig.»
Och se, medan han ännu talade, kom Judas, en av de tolv, och jämte honom en stor folkskara, med svärd och stavar, utsänd från översteprästerna och folkets äldste.
Men förrädaren hade givit dem ett tecken; han hade sagt: »Den som jag kysser, den är det; honom skolen I gripa.»
Och han trädde nu strax fram till Jesus och sade: »Hell dig, rabbi!» och kysste honom häftigt.
Jesus sade till honom: »Min vän, gör vad du är här för att göra.»
Då stego de fram och grepo Jesus och togo honom fången.
Men en av dem som voro med Jesus förde handen till sitt svärd och drog ut det och högg till översteprästens tjänare och högg så av honom örat.
Då sade Jesus till honom: »Stick ditt svärd tillbaka i skidan: ty alla som taga till svärd skola förgöras genom svärd.
Eller menar du att jag icke kunde utbedja mig av min Fader, att han nu sände till min tjänst mer än tolv legioner änglar?
Men huru bleve då skrifterna fullbordade, som säga att så måste ske?»
I samma stund sade Jesus till folkskaran: »Såsom mot en rövare haven I gått ut med svärd och stavar för att fasttaga mig.
Var dag har jag suttit i helgedomen och undervisat, utan att I haven gripit mig.
Men allt detta har skett, för att profeternas skrifter skola fullbordas.»
Då övergåvo alla lärjungarna honom och flydde.
Men de som hade gripit Jesus förde honom bort till översteprästen Kaifas, hos vilken de skriftlärde och de äldste hade församlat sig.
Och Petrus följde honom på avstånd ända till översteprästens gård; där gick han in och satte sig bland rättstjänarna för att se vad slutet skulle bliva.
Och översteprästerna och hela Stora rådet sökte efter något falskt vittnesbörd mot Jesus, för att kunna döda honom;
men fastän många falska vittnen trädde fram, funno de likväl intet.
Slutligen trädde dock två män fram
och sade: »Denne har sagt: 'Jag kan bryta ned Guds tempel och på tre dagar bygga upp det igen.'»
Då stod översteprästen upp och sade till honom: »Svarar du intet?
Huru är det med det som dessa vittna mot dig?»
Men Jesus teg.
Då sade översteprästen till honom: »Jag besvär dig vid den levande Guden, att du säger oss om du är Messias, Guds Son.»
Jesus svarade honom: »Du har själv sagt det.
Men jag säger eder: Härefter skolen I få se Människosonen sitta på Maktens högra sida och komma på himmelens skyar.»
Då rev översteprästen sönder sina kläder och sade: »Han har hädat.
Vad behöva vi mer några vittnen?
I haven nu hört hädelsen.
Vad synes eder?»
De svarade och sade: »Han är skyldig till döden.»
Därefter spottade man honom i ansiktet och slog honom på kinderna, den ene med knytnäven, den andre med flata handen,
och sade: »Profetera för oss, Messias: vem var det som slog dig?»
Men Petrus satt utanför på gården.
Då kom en tjänstekvinna fram till honom och sade: »Också du var med Jesus från Galileen.»
Men han nekade inför alla och sade: »Jag förstår icke vad du menar.»
När han sedan hade kommit ut i porten, fick en annan kvinna se honom och sade till dem som voro där: »Denne var med Jesus från Nasaret.»
Åter nekade han med en ed och sade: »Jag känner icke den mannen.»
Litet därefter kommo de kringstående fram och sade till Petrus: »Förvisso är också du en av dem; redan ditt uttal röjer dig ju.»
Då begynte han förbanna sig och svärja: »Jag känner icke den mannen.»
Och i detsamma gol hanen.
Då kom Petrus ihåg Jesu ord, huru han hade sagt: »Förrän hanen gal, skall du tre gånger förneka mig.»
Och han gick ut och grät bitterligen.
Men när det hade blivit morgon, fattade alla översteprästerna och folkets äldste det beslutet angående Jesus, att de skulle döda honom.
Och de läto binda honom och förde honom bort och överlämnade honom åt Pilatus, landshövdingen.
När då Judas, som hade förrått honom, såg att han var dömd, ångrade han sig och bar de trettio silverpenningarna tillbaka till översteprästerna och de äldste
och sade: »Jag har syndat därigenom att jag har förrått oskyldigt blod.»
Men de svarade: »Vad kommer det oss vid?
Du får själv svara därför.»
Då kastade han silverpenningarna i templet och gick sin väg.
Sedan gick han bort och hängde sig.
Men översteprästerna togo silverpenningarna och sade: »Det är icke lovligt att lägga dem i offerkistan, eftersom det är blodspenningar.»
Och sedan de hade fattat sitt beslut, köpte de för dem Krukmakaråkern till begravningsplats för främlingar.
Därför kallas den åkern ännu i dag Blodsåkern.
Så fullbordades det som var sagt genom profeten Jeremias, när han sade: »Och jag tog de trettio silverpenningarna -- priset för den man vilkens värde hade blivit bestämt, den som israelitiska män hade värderat --
och jag gav dem till betalning för Krukmakaråkern, i enlighet med Herrens befallning till mig.»
Men Jesus ställdes fram inför landshövdingen.
Och landshövdingen frågade honom och sade: »Är du judarnas konung?»
Jesus svarade honom: »Du säger det själv.»
Men när översteprästerna och de äldste framställde sina anklagelser mot honom, svarade han intet.
Då sade Pilatus till honom: »Hör du icke huru mycket de hava att vittna mot dig?»
Men han svarade honom icke på en enda fråga, så att landshövdingen mycket förundrade sig.
Nu var det sed att landshövdingen vid högtiden gav folket en fånge lös, vilken de ville.
Och man hade då en beryktad fånge, som hette Barabbas.
När de nu voro församlade, frågade Pilatus dem: »Vilken viljen I att jag skall giva eder lös, Barabbas eller Jesus, som kallas Messias?»
Han visste nämligen att det var av avund som man hade dragit Jesus inför rätta.
Och medan han satt på domarsätet, hade hans hustru sänt bud till honom och låtit säga: »Befatta dig icke med denne rättfärdige man; ty jag har i natt lidit mycket i drömmen för hans skull.»
Men översteprästerna och de äldste hade övertalat folket att begära Barabbas och låta förgöra Jesus.
När alltså landshövdingen nu frågade dem och sade: »Vilken av de två viljen I att jag skall giva eder lös?», så svarade de: »Barabbas.»
Då frågade Pilatus dem: »Vad skall jag då göra med Jesus, som kallas Messias?»
De svarade alla: »Låt korsfästa honom.»
Men han frågade: »Vad ont har han då gjort?»
Då skriade de ännu ivrigare: »Låt korsfästa honom.»
När nu Pilatus såg att han intet kunde uträtta, utan att larmet blev allt starkare, lät han hämta vatten och tvådde sina händer i folkets åsyn och sade: »Jag är oskyldig till denne mans blod.
I fån själva svara därför.»
Och allt folket svarade och sade: »Hans blod komme över oss och över våra barn.»
Då gav han dem Barabbas lös; men Jesus lät han gissla och utlämnade honom sedan till att korsfästas.
Då togo landshövdingens krigsmän Jesus med sig in i pretoriet och församlade hela den romerska vakten omkring honom.
Och de togo av honom hans kläder och satte på honom en röd mantel
och vredo samman en krona av törnen och satte den på hans huvud, och i hans högra hand satte de ett rör.
Sedan böjde de knä inför honom och begabbade honom och sade: »Hell dig, judarnas konung!»
Och de spottade på honom och togo röret och slogo honom därmed i huvudet.
Och när de så hade begabbat honom, klädde de av honom manteln och satte på honom hans egna kläder och förde honom bort till att korsfästas.
Då de nu voro på väg ditut, träffade de på en man från Cyrene, som hette Simon.
Honom tvingade de att gå med och bära hans kors.
Och när de hade kommit till en plats som kallades Golgata (det betyder huvudskalleplats),
räckte de honom vin att dricka, blandat med galla; men då han hade smakat därpå, ville han icke dricka det.
Och när de hade korsfäst honom, delade de hans kläder mellan sig genom att kasta lott om dem.
Sedan sutto de där och höllo vakt om honom.
Och över hans huvud hade man satt upp en överskrift, som angav vad han var anklagad för, och den lydde så: »Denne är Jesus, judarnas konung.»
Med honom korsfästes då ock två rövare, den ene på högra sidan och den andre på vänstra.
Och de som gingo där förbi bespottade honom och skakade huvudet
och sade: »Du som bryter ned templet och inom tre dagar bygger upp det igen, hjälp dig nu själv, om du är Guds Son, och stig ned från korset.»
Sammalunda talade ock översteprästerna, jämte de skriftlärde och de äldste, begabbande ord och sade:
»Andra har han hjälpt; sig själv kan han icke hjälpa.
Han är ju Israels konung; han stige nu ned från korset, så vilja vi tro på honom.
Han har satt sin förtröstan på Gud, må nu han frälsa honom, om han har behag till honom, han har ju sagt: 'Jag är Guds Son.'»
På samma sätt smädade honom också rövarna som voro korsfästa med honom.
Men vid sjätte timmen kom över hela landet ett mörker, som varade ända till nionde timmen.
Och vid nionde timmen ropade Jesus med hög röst och sade: »Eli, Eli, lema sabaktani?»; det betyder: »Min Gud, min Gud, varför har du övergivit mig?»
Men när några av dem som stodo där borde detta, sade de: »Han kallar på Elias.»
Och strax skyndade en av dem fram och tog en svamp och fyllde den med ättikvin och satte den på ett rör och gav honom att dricka.
Men de andra sade: »Låt oss se om Elias kommer och hjälper honom.»
Åter ropade Jesus med hög röst och gav upp andan.
Och se, då rämnade förlåten i templet i två stycken, uppifrån och ända ned, och jorden skalv, och klipporna rämnade,
och gravarna öppnades, och många avsomnade heligas kroppar stodo upp.
De gingo ut ur sina gravar och kommo efter hans uppståndelse in i den heliga staden och uppenbarade sig för många.
Men när hövitsmannen och de som med honom höllo vakt om Jesus sågo jordbävningen och det övriga som skedde, blevo de mycket förskräckta och sade: »Förvisso var denne Guds Son.»
Och många kvinnor som hade följt Jesus från Galileen och tjänat honom, stodo där på avstånd och sågo vad som skedde.
Bland dessa voro Maria från Magdala och den Maria som var Jakobs och Joses' moder, så ock Sebedeus' söners moder.
Men när det hade blivit afton, kom en rik man från Arimatea, vid namn Josef, som ock hade blivit en Jesu lärjunge;
denne gick till Pilatus och utbad sig att få Jesu kropp.
Då bjöd Pilatus att man skulle lämna ut den åt honom.
Och Josef tog hans kropp och svepte den i en ren linneduk
och lade den i den nya grav som han hade låtit hugga ut åt sig i klippan; och sedan han hade vältrat en stor sten för ingången till graven, gick han därifrån.
Men Maria från Magdala och den andra Maria voro där, och de sutto gent emot graven.
Följande dag, som var dagen efter tillredelsedagen, församlade sig översteprästerna och fariséerna och gingo till Pilatus
och sade: »Herre, vi hava dragit oss till minnes att den villoläraren sade, medan han ännu levde: 'Efter tre dagar skall jag uppstå.'
Bjud fördenskull att man skyddar graven intill tredje dagen, så att hans lärjungar icke komma och stjäla bort honom, och sedan säga till folket att han har uppstått från de döda.
Då bliver den sista villan värre än den första.»
Pilatus svarade dem: »Där haven I vakt; gån åstad och skydden graven så gott I kunnen.»
Och de gingo åstad och skyddade graven, i det att de icke allenast satte ut vakten, utan ock förseglade stenen.
När sabbaten hade gått till ända, i gryningen till första veckodagen, kommo Maria från Magdala och den andra Maria för att se graven.
Då blev det en stor jordbävning; ty en Herrens ängel steg ned från himmelen och gick fram och vältrade bort stenen och satte sig på den.
Och han var att skåda såsom en ljungeld, och hans kläder voro vita såsom snö.
Och väktarna skälvde av förskräckelse för honom och blevo såsom döda.
Men ängeln talade och sade till kvinnorna: »Varen I icke förskräckta; jag vet att I söken Jesus, den korsfäste.
Han är icke här, ty han är uppstånden, såsom han hade förutsagt.
Kommen hit, och sen platsen där han har legat.
Och gån så åstad med hast, och sägen till hans lärjungar att han är uppstånden från de döda.
Och han skall före eder gå till Galileen; där skolen I få se honom.
Jag har nu sagt eder det.»
Och de gingo med hast bort ifrån graven, under fruktan och med stor glädje, och skyndade åstad för att omtala det för hans lärjungar.
Men se, då kom Jesus emot dem och sade: »Hell eder!»
Och de gingo fram och fattade om hans fötter och tillbådo honom.
Då sade Jesus till dem: »Frukten icke; gån åstad och omtalen detta för mina bröder, på det att de må gå till Galileen; där skola de få se mig.»
Men under det att de voro på vägen, kommo några av väktarna till staden och underrättade översteprästerna om allt det som hade hänt.
Då församlade sig dessa jämte de äldste; och sedan de hade fattat sitt beslut, gåvo de en ganska stor summa penningar åt krigsmännen
och sade: »Så skolen I säga: 'Hans lärjungar kommo om natten och stulo bort honom, medan vi sovo.'
Och om saken kommer för landshövdingens öron, så skola vi ställa honom till freds och sörja för, att I kunnen vara utan bekymmer.»
Och de togo emot penningarna och gjorde såsom man hade lärt dem.
Och det talet utspriddes bland judarna och är gängse bland dem ännu i denna dag.
Men de elva lärjungarna begåvo sig till det berg i Galileen, dit Jesus hade bjudit dem att gå.
Och när de fingo se honom, tillbådo de honom.
Dock funnos några som tvivlade.
Då trädde Jesus fram och talade till dem och sade: »Mig är given all makt i himmelen och på jorden.
Gån fördenskull ut och gören alla folk till lärjungar, döpande dem i Faderns och Sonens och den helige Andes namn,
lärande dem att hålla allt vad jag har befallt eder.
Och se, jag är med eder alla dagar intill tidens ände.»
Detta är begynnelsen av evangelium om Jesus Kristus, Guds Son.
Så är skrivet hos profeten Esaias: »Se, jag sänder ut min ängel framför dig, och han skall bereda vägen för dig.
Hör rösten av en som ropar i öknen: 'Bereden vägen för Herren, gören stigarna jämna för honom.'»
I enlighet härmed uppträdde Johannes döparen i öknen och predikade bättringens döpelse till syndernas förlåtelse.
Och hela judiska landet och alla Jerusalems invånare gingo ut till honom och läto döpa sig av honom i floden Jordan, och bekände därvid sina synder.
Och Johannes hade kläder av kamelhår och bar en lädergördel om sina länder och levde av gräshoppor och vildhonung.
Och han predikade och sade: »Efter mig kommer den som är starkare än jag; jag är icke ens värdig att böja mig ned för att upplösa hans skorem.
Jag döper eder med vatten, men han skall döpa eder med helig ande.»
Och det hände sig vid den tiden att Jesus kom från Nasaret i Galileen.
Och han lät döpa sig i Jordan av Johannes.
Och strax då han steg upp ur vattnet, såg han himmelen dela sig och Anden såsom en duva sänka sig ned över honom.
Och en röst kom från himmelen: »Du är min älskade Son; i dig har jag funnit behag.»
Strax därefter förde Anden honom ut i öknen.
Och han var i öknen i fyrtio dagar och frestades av Satan och levde bland vilddjuren; och änglarna betjänade honom.
Men sedan Johannes hade blivit satt i fängelse, kom Jesus till Galileen och predikade Guds evangelium
och sade: »Tiden är fullbordad, och Guds rike är nära; gören bättring, och tron evangelium.»
När han nu gick fram utmed Galileiska sjön, fick han se Simon och Simons broder Andreas kasta ut nät i sjön, ty de voro fiskare.
Och Jesus sade till dem: »Följen mig, så skall jag göra eder till människofiskare.»
Strax lämnade de näten och följde honom.
När han hade gått litet längre fram, fick han se Jakob, Sebedeus' son, och Johannes, hans broder, där de sutto i båten, också de, och ordnade sina nät.
Och strax kallade han dem till sig; och de lämnade sin fader Sebedeus med legodrängarna kvar i båten och följde honom.
Sedan begåvo de sig in i Kapernaum; och strax, på sabbaten, gick han in i synagogan och undervisade.
Och folket häpnade över hans förkunnelse; ty han förkunnade sin lära för dem med makt och myndighet, och icke såsom de skriftlärde.
Strax härefter befann sig i deras synagoga en man som var besatt av en oren ande.
Denne ropade
och sade: »Vad har du med oss att göra, Jesus från Nasaret?
Har du kommit för att förgöra oss?
Jag vet vem du är, du Guds Helige.»
Men Jesus tilltalade honom strängt och sade: »Tig, och far ut ur honom.»
Då slet och ryckte den orene anden honom och ropade med hög röst och for ut ur honom.
Och alla häpnade, så att de begynte fråga varandra och säga: »Vad är detta?
Det är ju en ny lära, med makt och myndighet.
Till och med de orena andarna befaller han, och de lyda honom.»
Och ryktet om honom gick strax ut överallt i hela den kringliggande trakten av Galileen.
Och strax då de hade kommit ut ur synagogan, begåvo de sig med Jakob och Johannes till Simons och Andreas' hus.
Men Simons svärmoder låg sjuk i feber, och de talade strax med honom om henne.
Då gick han fram och tog henne vid handen och reste upp henne; och febern lämnade henne, och hon betjänade dem.
Men när solen hade gått ned och det hade blivit afton, förde man till honom alla som voro sjuka eller besatta;
och hela staden var församlad utanför dörren.
Och han botade många som ledo av olika slags sjukdomar; och han drev ut många onda andar, men tillstadde icke de onda andarna att tala, eftersom de kände honom.
Och bittida om morgonen, medan det ännu var mörkt, stod han upp och gick åstad bort till en öde trakt, och bad där.
Men Simon och de som voro med honom skyndade efter honom.
Och när de funno honom, sade de till honom: »Alla fråga efter dig.»
Då sade han till dem: »Låt oss draga bort åt annat håll, till de närmaste småstäderna, för att jag också där må predika; ty därför har jag begivit mig ut.»
Och han gick åstad och predikade i hela Galileen, i deras synagogor, och drev ut de onda andarna.
Och en spetälsk man kom fram till honom och föll på knä och bad honom och sade till honom: »Vill du, så kan du göra mig ren.»
Då förbarmade han sig och räckte ut handen och rörde vid honom och sade till honom: »Jag vill; bliv ren.»
Och strax vek spetälskan ifrån honom, och han blev ren.
Sedan vände Jesus strax bort honom med stränga ord
och sade till honom: »Se till, att du icke säger något härom för någon; men gå bort och visa dig för prästen, och frambär för din rening det offer som Moses har påbjudit, till ett vittnesbörd för dem.»
Men när han kom ut, begynte han ivrigt förkunna och utsprida vad som hade skett, så att Jesus icke mer kunde öppet gå in i någon stad, utan måste hålla sig ute i öde trakter; och dit kom man till honom från alla håll.
Några dagar därefter kom han åter till Kapernaum; och när det spordes att han var hemma,
församlade sig så mycket folk, att icke ens platsen utanför dörren mer kunde rymma dem; och han förkunnade ordet för dem.
Då kommo de till honom med en lam man, som bars dit av fyra män.
Och då de för folkets skull icke kunde komma fram till honom med mannen, togo de bort taket över platsen där han var; och sedan de så hade gjort en öppning, släppte de ned sängen, som den lame låg på.
När Jesus såg deras tro, sade han till den lame: »Min son, dina synder förlåtas dig.»
Nu sutto där några skriftlärde, och dessa tänkte i sina hjärtan:
»Huru kan denne tala så?
Han hädar ju.
Vem kan förlåta synder, utom Gud allena?»
Strax förnam då Jesus i sin ande att de tänkte så vid sig själva; och han sade till dem: »Huru kunnen I tänka sådant i edra hjärtan?
Vilket är lättare, att säga till den lame: 'Dina synder förlåtas dig' eller att säga: 'Stå upp, tag din säng och gå'?
Men för att I skolen veta att Människosonen har makt här på jorden att förlåta synder,
så säger jag dig» (och härmed vände han sig till den lame): »Stå upp, tag din säng och gå hem.»
Då stod han upp och tog strax sin säng och gick ut i allas åsyn, så att de alla uppfylldes av häpnad och prisade Gud och sade: »Sådant hava vi aldrig sett.»
Åter begav han sig ut och gick längs med sjön.
Och allt folket kom till honom, och han undervisade dem.
När han nu gick där fram, fick han se Levi, Alfeus' son, sitta vid tullhuset.
Och han sade till denne: »Följ mig.»
Då steg han upp och följde honom.
När Jesus därefter låg till bords i hans hus, voro där såsom bordsgäster, jämte Jesus och hans lärjungar, också många publikaner och syndare; ty många sådana funnos bland dem som följde honom.
Men när de skriftlärde bland fariséerna sågo att han åt med publikaner och syndare, sade de till hans lärjungar: »Huru kan han äta med publikaner och syndare?»
När Jesus hörde detta, sade han till dem: »Det är icke de friska som behöva läkare, utan de sjuka.
Jag har icke kommit för att kalla rättfärdiga, utan för att kalla syndare.»
Och Johannes' lärjungar och fariséerna höllo fasta.
Och man kom och sade till honom: »Varför fasta icke dina lärjungar, då Johannes' lärjungar och fariséernas lärjungar fasta?»
Jesus svarade dem: »Kunna väl bröllopsgästerna fasta, medan brudgummen ännu är hos dem?
Nej, så länge de hava brudgummen hos sig, kunna de icke fasta.
Men den tid skall komma, då brudgummen tages ifrån dem, och då, på den tiden, skola de fasta. --
Ingen syr en lapp av okrympt tyg på en gammal mantel; om någon så gjorde, skulle det isatta nya stycket riva bort ännu mer av den gamla manteln, och hålet skulle bliva värre.
Ej heller slår någon nytt vin i gamla skinnläglar; om någon så gjorde, skulle vinet spränga sönder läglarna, så att både vinet och läglarna fördärvades.
Nej, nytt vin slår man i nya läglar.»
Och det hände sig på sabbaten att han tog vägen genom ett sädesfält; och hans lärjungar begynte rycka av axen, medan de gingo.
Då sade fariséerna till honom: »Se!
Huru kunna de på sabbaten göra vad som icke är lovligt?»
Han svarade dem: »Haven I aldrig läst vad David gjorde, när han själv och de som följde honom kommo i nöd och blevo hungriga:
huru han då, på den tid Abjatar var överstepräst, gick in i Guds hus och åt skådebröden -- fastän det ju icke är lovligt för andra än för prästerna att äta sådant bröd -- och huru han jämväl gav åt dem som följde honom?»
Därefter sade han till dem: »Sabbaten blev gjord för människans skull, och icke människan för sabbatens skull.
Så år då Människosonen herre också över sabbaten.»
Och han gick åter in i en synagoga.
Där var då en man som hade en förvissnad hand.
Och de vaktade på honom, för att se om han skulle bota denne på sabbaten; de ville nämligen få något att anklaga honom för.
Då sade han till mannen som hade den förvissnade handen: »Stå upp, och kom fram.»
Sedan sade han till dem: »Vilketdera är lovligt på sabbaten: att göra vad gott är, eller att göra vad ont är, att rädda någons liv, eller att döda?»
Men de tego.
Då såg han sig omkring på dem med vrede, bedrövad över deras hjärtans förstockelse, och sade till mannen: »Räck ut din hand.»
Och han räckte ut den; och hans hand blev frisk igen. --
Då gingo fariséerna bort och fattade strax, tillsammans med herodianerna, det beslutet att de skulle förgöra honom.
Och Jesus drog sig med sina lärjungar undan till sjön, och en stor hop folk följde honom från Galileen.
Och från Judeen och Jerusalem och Idumeen och från landet på andra sidan Jordan och från trakterna omkring Tyrus och Sidon kom en stor hop folk till honom, när de fingo höra huru stora ting han gjorde.
Och han tillsade sina lärjungar att en båt skulle hållas tillreds åt honom, för folkets skull, för att de icke skulle tränga sig inpå honom.
Ty han botade många och blev därför överlupen av alla som hade någon plåga och fördenskull ville röra vid honom.
Och när de orena andarna sågo honom, föllo de ned för honom och och ropade och sade: »Du är Guds Son.»
Men han förbjöd dem strängeligen, åter och åter, att röja honom.
Och han gick upp på berget och kallade till sig några som han själv utsåg; och de kommo till honom.
Så förordnade han tolv som skulle följa honom, och som han ville sända ut till att predika,
och de skulle hava makt att bota sjuka och driva ut onda andar.
Han förordnade alltså dessa tolv: Simon, åt vilken han gav tillnamnet Petrus;
vidare Jakob, Sebedeus' son, och Johannes, Jakobs broder, åt vilka han gav tillnamnet Boanerges (det betyder tordönsmän);
vidare Andreas och Filippus och Bartolomeus och Matteus och Tomas och Jakob, Alfeus' son, och Taddeus och Simon ivraren
och Judas Iskariot, densamme som förrådde honom.
Och när han kom hem, församlade sig folket åter, så att de icke ens fingo tillfälle att äta.
Då nu hans närmaste fingo höra härom, gingo de åstad för att taga vara på honom; ty de menade att han var från sina sinnen.
Och de skriftlärde som hade kommit ned från Jerusalem sade att han var besatt av Beelsebul, och att det var med de onda andarnas furste som han drev ut de onda andarna.
Då kallade han dem till sig och sade till dem i liknelser: »Huru skulle Satan kunna driva ut Satan?
Om ett rike har kommit i strid med sig självt, så kan det riket ju icke hava bestånd;
och om ett hus har kommit i strid med sig självt, så skall icke heller det huset kunna äga bestånd.
Om alltså Satan har satt sig upp mot sig själv och kommit i strid med sig själv, så kan han icke äga bestånd, utan det är då ute med honom. --
Nej, ingen kan gå in i en stark mans hus och plundra honom på hans bohag, såframt han icke förut har bundit den starke.
Först därefter kan han plundra hans hus.
Sannerligen säger jag eder: Alla andra synder skola bliva människors barn förlåtna, ja ock alla andra hädelser, huru hädiskt de än må tala;
men den som hädar den helige Ande, han får icke någonsin förlåtelse, utan är skyldig till evig synd.»
De hade ju nämligen sagt att han var besatt av en oren ande.
Så kommo nu hans moder och hans bröder; och de stannade därutanför och sände bud in till honom för att kalla honom ut.
Och mycket folk satt där omkring honom; och man sade till honom: »Se, din moder och dina bröder stå härutanför och fråga efter dig.»
Då svarade han dem och sade: Vilken är min moder, och vilka äro mina bröder?»
Och han såg sig omkring på dem som sutto där runt omkring honom, och han sade: »Se här är min moder, och här äro mina bröder!
Den som gör Guds vilja, den är min broder och min syster och min moder.»
Och han begynte åter undervisa vid sjön.
Och där församlade sig en stor hop folk omkring honom.
Därför steg han i en båt; och han satt i den ute på sjön, under det att allt folket stod på land utmed sjön.
Och han undervisade dem mycket i liknelser och sade till dem i sin undervisning:
»Hören!
En såningsman gick ut för att så.
Då hände sig, när han sådde, att somt föll vid vägen, och fåglarna kommo och åto upp det.
Och somt föll på stengrund, där det icke hade mycket jord, och det kom strax upp, eftersom det icke hade djup jord;
men när solen hade gått upp, förbrändes det, och eftersom det icke hade någon rot, torkade det bort.
Och somt föll bland törnen, och törnena sköto upp och förkvävde det, så att det icke gav någon frukt.
Men somt föll i god jord, och det sköt upp och växte och gav frukt och bar trettiofalt och sextiofalt och hundrafalt.»
Och han tillade: »Den som har öron till att höra, han höre.»
När han sedan hade dragit sig undan ifrån folket, frågade honom de tolv, och med dem de andra som följde honom, om liknelserna.
Då sade han till dem: »Åt eder är Guds rikes hemlighet given, men åt dem som stå utanför meddelas alltsammans i liknelser,
för att de 'med seende ögon skola se, och dock intet förnimma, och med hörande öron höra, och dock intet förstå, så att de icke omvända sig och undfå förlåtelse'.»
Sedan sade han till dem: »Förstån I icke denna liknelse, huru skolen I då kunna fatta alla de andra liknelserna? --
Vad såningsmannen sår är ordet.
Och att säden såddes vid vägen, det är sagt om dem i vilka ordet väl bliver sått, men när de hava hört det, kommer strax Satan ock tager bort ordet som såddes i dem.
Sammalunda förhåller det sig med det som sås på stengrunden: det är sagt om dem, som när de få höra ordet, väl strax taga emot det med glädje,
men icke hava någon rot i sig, utan bliva beståndande allenast till en tid; när sedan bedrövelse eller förföljelse påkommer för ordets skull, då komma de strax på fall.
Annorlunda förhåller det sig med det som sås bland törnena: det är sagt om dem som väl höra ordet,
men låta tidens omsorger och rikedomens bedrägliga lockelse, och begärelser efter andra ting, komma därin och förkväva ordet, så att det bliver utan frukt.
Men att det såddes i den goda jorden, det är sagt om dem som både höra ordet och taga emot det, och som bära frukt, trettiofalt och sextiofalt och hundrafalt.»
Och han sade till dem: »Icke tager man väl fram ett ljus, för att det skall sättas under skäppan eller under bänken; man gör det ju, för att det skall sättas på ljusstaken.
Ty intet är fördolt, utom för att det skall bliva uppenbarat; ej heller har något blivit undangömt, utom för att det skall komma i dagen.
Om någon har öron till att höra, så höre han.»
Och han sade till dem: »Akten på vad I hören.
Med det mått som I mäten med skall ock mätas åt eder, och ännu mer skall bliva eder tilldelat.
Ty den som har, åt honom skall varda givet; men den som icke har, från honom skall tagas också det han har.»
Och han sade: »Så är det med Guds rike, som när en man sår säd i jorden;
och han sover, och han vaknar, och nätter och dagar gå, och säden skjuter upp och växer i höjden, han vet själv icke huru.
Av sig själv bär jorden frukt, först strå och sedan ax, och omsider finnes fullbildat vete i axet.
När så frukten är mogen, låter han strax lien gå, ty skördetiden är då inne.»
Och han sade: »Vad skola vi likna Guds rike vid, eller med vilken liknelse skola vi framställa det?
Det är såsom ett senapskorn, som när det lägges ned i jorden, är minst av alla frön på jorden;
men sedan det är nedlagt, skjuter det upp och bliver störst bland alla kryddväxter och får så stora grenar, att himmelens fåglar kunna bygga sina nästen i dess skugga.»
I många sådana liknelser förkunnade han ordet för dem, efter deras förmåga att fatta det;
och utan liknelse talade han icke till dem.
Men för sina lärjungar uttydde han allt, när de voro allena.
Samma dag, om aftonen, sade han till dem: »Låt oss fara över till andra stranden.»
Så läto de folket gå och togo honom med i båten, där han redan förut var; och jämväl andra båtar följde med honom.
Då kom en häftig stormvind, och vågorna slogo in i båten, så att båten redan begynte fyllas.
Men han själv låg i bakstammen och sov, lutad mot huvudgärden.
Då väckte de honom och sade till honom: »Mästare, frågar du icke efter att vi förgås?»
När han så hade vaknat, näpste han vinden och sade till sjön: »Tig, var stilla.»
Och vinden lade sig, och det blev alldeles lugnt.
Därefter sade han till dem: »Varför rädens I?
Haven I ännu ingen tro?»
Och de hade blivit mycket häpna och sade till varandra: »Vem är då denne, eftersom både vinden och sjön äro honom lydiga?»
Så kommo de över till gerasenernas land, på andra sidan sjön.
Och strax då han hade stigit ur båten, kom en man, som var besatt av en oren ande, emot honom från gravarna där;
han hade nämligen sitt tillhåll bland gravarna.
Och icke ens med kedjor kunde man numera fängsla honom;
ty väl hade han många gånger blivit fängslad med fotbojor och kedjor, men han hade slitit itu kedjorna och brutit sönder fotbojorna, och ingen kunde få makt med honom.
Och han vistades alltid, dag och natt, bland gravarna och på bergen och skriade och sargade sig själv med stenar.
När denne nu fick se Jesus på avstånd, skyndade han fram och föll ned för honom
och ropade med hög röst och sade: »Vad har du med mig att göra, Jesus, du Guds, den Högstes, Son?
Jag besvär dig vid Gud, plåga mig icke.»
Jesus skulle nämligen just säga till honom: »Far ut ur mannen, du orena ande.»
Då frågade han honom: »Vad är ditt namn?»
Han svarade honom: »Legion är mitt namn, ty vi äro många.»
Och han bad honom enträget att icke driva dem bort ifrån den trakten.
Nu gick där vid berget en stor svinhjord i bet.
Och de bådo honom och sade: »Sänd oss åstad in i svinen; låt oss få fara in i dem.»
Och han tillstadde dem det.
Då gåvo sig de orena andarna åstad och foro in i svinen.
Och hjorden, vid pass två tusen svin, störtade sig utför branten ned i sjön och drunknade i sjön.
Men de som vaktade dem flydde och berättade härom i staden och på landsbygden; och folket gick åstad för att se vad det var som hade skett.
När de då kommo till Jesus, fingo de se den som hade varit besatt, mannen som hade haft legionen i sig, sitta där klädd och vid sina sinnen; och de betogos av häpnad.
Och de som hade åsett händelsen förtäljde för dem vad som hade vederfarits den besatte, och vad som hade skett med svinen.
Då begynte folket bedja honom att han skulle gå bort ifrån deras område.
När han sedan steg i båten, bad honom mannen som hade varit besatt, att han skulle få följa honom.
Men han tillstadde honom det icke, utan sade till honom: »Gå hem till de dina, och berätta för dem huru stora ting Herren har gjort med dig, och huru han har förbarmat sig över dig.»
Då gick han åstad och begynte förkunna i Dekapolis huru stora ting Jesus hade gjort med honom; och alla förundrade sig.
Och när Jesus hade farit över i båten, tillbaka till andra stranden, församlade sig mycket folk omkring honom, där han stod vid sjön.
Då kom en synagogföreståndare, vid namn Jairus, dit; och när denne fick se honom, föll han ned för hans fötter
och bad honom enträget och sade: »Min dotter ligger på sitt yttersta.
Kom och lägg händerna på henne, så att hon bliver hulpen och får leva.»
Då gick han med mannen; och honom följde mycket folk, som trängde sig inpå honom.
Nu var där en kvinna som hade haft blodgång i tolv år,
och som hade lidit mycket hos många läkare och kostat på sig allt vad hon ägde, utan att det hade varit henne till något gagn; snarare hade det blivit värre med henne.
Hon hade fått höra om Jesus och kom nu i folkhopen, bakom honom, och rörde vid hans mantel.
Ty hon tänkte: »Om jag åtminstone får röra vid hans kläder, så bliver jag hulpen.»
Och strax uttorkade hennes blods källa, och hon kände i sin kropp att hon var botad från sin plåga.
Men strax då Jesus inom sig förnam vilken kraft som hade gått ut ifrån honom, vände han sig om i folkhopen och frågade: »Vem rörde vid mina kläder?»
Hans lärjungar sade till honom: »Du ser huru folket tränger på, och ändå frågar du: 'Vem rörde vid mig?'»
Då såg han sig omkring för att få se den som hade gjort detta.
Men kvinnan fruktade och bävade, ty hon visste vad som hade skett med henne; och hon kom fram och föll ned för honom och sade honom hela sanningen.
Då sade han till henne: »Min dotter, din tro har hjälpt dig.
Gå i frid, och var botad från din plåga.»
Medan han ännu talade, kommo några från synagogföreståndarens hus och sade: »Din dotter är död; du må icke vidare göra mästaren omak.»
Men när Jesus märkte vad som talades, sade han till synagogföreståndaren: »Frukta icke, tro allenast.»
Och han tillstadde ingen att följa med, utom Petrus och Jakob och Johannes, Jakobs broder.
Så kommo de till synagogföreståndarens hus, och han fick där se en hop människor som höjde klagolåt och gräto och jämrade sig högt.
Och han gick in och sade till dem: »Varför klagen I och gråten?
Flickan är icke död, hon sover.»
Då hånlogo de åt honom.
Men han visade ut dem allasammans; och han tog med sig allenast flickans fader och moder och dem som hade fått följa med honom, och gick in dit där flickan låg.
Och han tog flickan vid handen och sade till henne: »Talita, kum» (det betyder: »Flicka, jag säger dig, stå upp»).
Och strax stod flickan upp och begynte gå omkring (hon var nämligen tolv år gammal); och de blevo strax uppfyllda av stor häpnad.
Men han förbjöd dem strängeligen att låta någon få veta vad som hade skett.
Därefter tillsade han att man skulle giva henne något att äta.
Och han gick bort därifrån och begav sig till sin fädernestad; och hans lärjungar följde honom.
Och när det blev sabbat, begynte han undervisa i synagogan.
Och folket häpnade, när de hörde honom; de sade: »Varifrån har han fått detta?
Och vad är det för vishet som har blivit honom given?
Och dessa stora kraftgärningar som göras genom honom, varifrån komma de?
Är då denne icke timmermannen, han som är Marias son och broder till Jakob och Joses och Judas och Simon?
Och bo icke hans systrar här hos oss?»
Så blev han för dem en stötesten.
Då sade Jesus till dem: »En profet är icke föraktad utom i sin fädernestad och bland sina fränder och i sitt eget hus.»
Och han kunde icke där göra någon kraftgärning, utom att han botade några få sjuka, genom att lägga händerna på dem.
Och han förundrade sig över deras otro.
Sedan gick han omkring i byarna, från den ena byn till den andra, och undervisade.
Och han kallade till sig de tolv och sände så ut dem, två och två, och gav dem makt över de orena andarna.
Och han bjöd dem att icke taga något med sig på vägen, utom allenast en stav: icke bröd, icke ränsel, icke penningar i bältet.
Sandaler finge de dock hava på fötterna, men de skulle icke bära dubbla livklädnader.
Och han sade till dem: »När I haven kommit in i något hus, så stannen där, till dess I lämnen den orten.
Och om man på något ställe icke tager emot eder och icke hör på eder, så gån bort därifrån, och skudden av stoftet som är under edra fötter, till ett vittnesbörd mot dem.»
Och de gingo ut och predikade att man skulle göra bättring;
och de drevo ut många onda andar och smorde många sjuka med olja och botade dem.
Och konung Herodes fick höra om honom, ty hans namn hade blivit känt.
Man sade: »Det är Johannes döparen, som har uppstått från de döda, och därför verka dessa krafter i honom.»
Men andra sade: »Det är Elias.»
Andra åter sade: »Det är en profet, lik de andra profeterna.»
Men när Herodes hörde detta, sade han: »Det är Johannes, den som jag lät halshugga.
Han bar uppstått från de döda.»
Herodes hade nämligen sänt åstad och låtit gripa Johannes och binda honom och sätta honom i fängelse, för Herodias', sin broder Filippus' hustrus, skull.
Ty henne hade Herodes tagit till äkta,
och Johannes hade då sagt till honom: »Det är icke lovligt för dig att hava din broders hustru.»
Därför hyste nu Herodes agg till honom och ville döda honom, men han hade icke makt därtill.
Ty Herodes förstod att Johannes var en rättfärdig och helig man, och han fruktade för honom och gav honom sitt beskydd.
Och när han hade hört honom, blev han betänksam i många stycken; och han hörde honom gärna.
Men så kom en läglig dag, i det att Herodes på sin födelsedag gjorde ett gästabud för sina stormän och för krigsöverstarna och de förnämsta männen i Galileen.
Då gick Herodias' dotter ditin och dansade; och hon behagade Herodes och hans bordsgäster.
Och konungen sade till flickan: »Begär av mig vadhelst du vill, så skall jag giva dig det.»
Ja, han lovade henne detta med ed och sade: »Vadhelst du begär av mig, det skall jag giva dig, ända till hälften av mitt rike.»
Då gick hon ut och frågade sin moder: »Vad skall jag begära?»
Hon svarade: »Johannes döparens huvud.»
Och strax skyndade hon in till konungen och framställde sin begäran och sade: »Jag vill att du nu genast giver mig på ett fat Johannes döparens huvud.»
Då blev konungen mycket bekymrad, men för edens och för bordsgästernas skull ville han icke avvisa henne.
Alltså sände konungen strax en drabant med befallning att hämta hans huvud.
Och denne gick åstad och halshögg honom i fängelset
och bar sedan fram hans huvud på ett fat och gav det åt flickan, och flickan gav det åt sin moder.
Men när hans lärjungar fingo höra härom, kommo de och togo hans döda kropp och lade den i en grav.
Och apostlarna församlade sig hos Jesus och omtalade för honom allt vad de hade gjort, och allt vad de hade lärt folket.
Då sade han till dem: »Kommen nu I med mig bort till en öde trakt, där vi få vara allena, och vilen eder något litet.»
Ty de fingo icke ens tid att äta; så många voro de som kommo och gingo.
De foro alltså i båten bort till en öde trakt, där de kunde vara allena.
Men man såg dem fara sin väg, och många fingo veta det; och från alla städer strömmade då människor tillsammans dit landvägen och kommo fram före dem.
När han så steg i land, fick han se att där var mycket folk.
Då ömkade han sig över dem, eftersom de voro »lika får som icke hade någon herde»; och han begynte undervisa dem i mångahanda stycken.
Men när det redan var långt lidet på dagen, trädde hans lärjungar fram till honom och sade: »Trakten är öde, och det är redan långt lidet på dagen.
Låt dem skiljas åt, så att de kunna gå bort i gårdarna och byarna häromkring och köpa sig något att äta.»
Men han svarade och sade till dem: »Given I dem att äta.»
De svarade honom: »Skola vi då gå bort och köpa bröd för två hundra silverpenningar och giva dem att äta?»
Men han sade till dem: »Huru många bröd haven I?
Gån och sen efter.»
Sedan de hade gjort så, svarade de: »Fem, och därtill två fiskar.»
Då befallde han dem att låta alla i skilda matlag lägga sig ned i gröna gräset.
Och de lägrade sig där i skilda hopar, hundra eller femtio i var.
Därefter tog han de fem bröden och de två fiskarna och såg upp till himmelen och välsignade dem.
Och han bröt bröden och gav dem åt lärjungarna, för att de skulle lägga fram åt folket; också de två fiskarna delade han mellan dem alla.
Och de åto alla och blevo mätta.
Sedan samlade man upp överblivna brödstycken, tolv korgar fulla, därtill ock kvarlevor av fiskarna.
Och det var fem tusen män som hade ätit.
Strax därefter nödgade han sina lärjungar att stiga i båten och i förväg fara över till Betsaida på andra stranden, medan han själv tillsåg att folket skildes åt.
Och när han hade tagit avsked av folket, gick han därifrån upp på berget för att bedja.
När det så hade blivit afton, var båten mitt på sjön, och han var ensam kvar på land.
Och han såg dem vara hårt ansatta, där de rodde fram, ty vinden låg emot dem.
Vid fjärde nattväkten kom han då till dem, gående på sjön, och skulle just gå förbi dem.
Men när de fingo se honom gå på sjön, trodde de att det var en vålnad och ropade högt;
ty de sågo honom alla och blevo förfärade.
Men han begynte strax tala med dem och sade till dem: »Varen vid gott mod; det är jag, varen icke förskräckta.»
Därefter steg han upp till dem i båten, och vinden lade sig.
Och de blevo uppfyllda av stor häpnad;
ty de hade icke kommit till förstånd genom det som hade skett med bröden, utan deras hjärtan voro förstockade.
När de hade farit över till andra stranden, kommo de till Gennesarets land och lade till där.
Och när de stego ur båten, kände man strax igen honom;
och man skyndade omkring med bud i hela den trakten, och folket begynte då överallt bära de sjuka på sängar dit där man hörde att han var.
Och varhelst han gick in i någon by eller någon stad eller någon gård, där lade man de sjuka på de öppna platserna.
Och de bådo honom att åtminstone få röra vid hörntofsen på hans mantel; och alla som rörde vid den blevo hulpna.
Och fariséerna, så ock några skriftlärde som hade kommit från Jerusalem, församlade sig omkring honom;
och de fingo då se några av hans lärjungar äta med »orena», det är otvagna, händer.
Nu är det så med fariséerna och alla andra judar, att de icke äta något utan att förut, till åtlydnad av de äldstes stadgar, noga hava tvagit sina händer,
likasom de icke heller, när de komma från torget, äta något utan att förut hava tvagit sig; många andra stadgar finnas ock, som de av ålder pläga hålla, såsom att skölja bägare och träkannor och kopparskålar.
Därför frågade honom nu fariséerna och de skriftlärde: »Varför vandra icke dina lärjungar efter de äldstes stadgar, utan äta med orena händer?»
Men han svarade dem: »Rätt profeterade Esaias om eder, I skrymtare, såsom det är skrivet: 'Detta folk ärar mig med sina läppar, men deras hjärtan äro långt ifrån mig;
och fåfängt dyrka de mig, eftersom de läror de förkunna äro människobud.'
I sätten Guds bud å sido och hållen människors stadgar.»
Ytterligare sade han till dem: »Rätt så; I upphäven Guds bud för att hålla edra egna stadgar!
Moses har ju sagt: 'Hedra din fader och din moder' och 'Den som smädar sin fader eller sin moder, han skall döden dö.'
Men I sägen: om en son säger till sin fader eller sin moder: 'Vad du av mig kunde hava fått till hjälp, det giver jag i stället såsom korban' (det betyder offergåva),
då kunnen I icke tillstädja honom att vidare göra något för sin fader eller sin moder.
På detta sätt gören I Guds budord om intet genom edra fäderneärvda stadgar.
Och mycket annat sådant gören I.»
Därefter kallade han åter folket till sig och sade till dem: »Hören mig alla och förstån.
Intet som utifrån går in i människan kan orena henne, men vad som går ut ifrån människan, detta är det som orenar henne.»
245490
När han sedan hade lämnat folket och kommit inomhus, frågade hans lärjungar honom om detta bildliga tal.
Han svarade dem: »Ären då också I så utan förstånd?
Insen I icke att intet som utifrån går in i människan kan orena henne,
eftersom det icke går in i hennes hjärta, utan ned i buken, och har sin naturliga utgång?»
Härmed förklarade han all mat för ren.
Och han tillade: »Vad som går ut ifrån människan, detta är det som orenar människan.
Ty inifrån, från människornas hjärtan, utgå deras onda tankar, otukt, tjuveri, mord,
äktenskapsbrott, girighet, ondska, svek, lösaktighet, avund, hädelse, övermod, oförsynt väsende.
Allt detta onda går inifrån ut, och det orenar människan.»
Och han stod upp och begav sig bort därifrån till Tyrus' område.
Där gick han in i ett hus och ville icke att någon skulle få veta det.
Dock kunde han icke förbliva obemärkt,
utan en kvinna, vilkens dotter var besatt av en oren ande, kom, strax då hon hade fått höra om honom, och föll ned för hans fötter;
det var en grekisk kvinna av syrofenicisk härkomst.
Och hon bad honom att han skulle driva ut den onde anden ur hennes dotter.
Men han sade till henne: »Låt barnen först bliva mättade; det är ju otillbörligt att taga brödet från barnen och kasta det åt hundarna.»
Hon svarade och sade till honom: »Ja, Herre; också äta hundarna under bordet allenast av barnens smulor.»
Då sade han till henne: »För det ordets skull säger jag dig: Gå; den onde anden har farit ut ur din dotter.»
Och när hon kom hem, fann hon flickan ligga på sängen och såg att den onde anden hade farit ut.
Sedan begav han sig åter bort ifrån Tyrus' område och tog vägen över Sidon och kom, genom Dekapolis' område, till Galileiska sjön.
Och man förde till honom en som var döv och nästan stum och bad honom att lägga handen på denne.
Då tog han honom avsides ifrån folket och satte sina fingrar i hans öron och spottade och rörde vid hans tunga
och såg upp till himmelen, suckade och sade till honom: »Effata» (det betyder: »Upplåt dig»).
Då öppnades hans öron, och hans tungas band löstes, och han talade redigt och klart.
Och Jesus förbjöd dem att omtala detta för någon; men ju mer han förbjöd dem, dess mer förkunnade de det.
Och folket häpnade övermåttan och sade: »Allt har han väl beställt: de döva låter han höra och de stumma tala.»
Då vid samma tid åter mycket folk hade kommit tillstädes, och de icke hade något att äta, kallade han sina lärjungar till sig och sade till dem:
»Jag ömkar mig över folket, ty det är redan tre dagar som de hava dröjt kvar hos mig, och de hava intet att äta.
Om jag nu låter dem fastande gå ifrån mig hem, så uppgivas de på vägen; somliga av dem hava ju kommit långväga ifrån.»
Då svarade hans lärjungar honom: »Varifrån skall man här i en öken kunna få bröd till att mätta dessa med?»
Han frågade dem: »Huru många bröd haven I?»
De svarade: »Sju.»
Då tillsade han folket att lägra sig på marken.
Ock han tog de sju bröden, tackade Gud och bröt dem och gav åt sina lärjungar, för att de skulle lägga fram dem; och de lade fram åt folket.
De hade ock några få småfiskar; och när han hade välsignat dessa, bjöd han att man likaledes skulle lägga fram dem.
Så åto de och blevo mätta.
Och man samlade sedan upp sju korgar med överblivna stycken.
Men antalet av dem som voro tillstädes var vid pass fyra tusen.
Sedan lät han dem skiljas åt.
Och strax därefter steg han i båten med sina lärjungar och for till trakten av Dalmanuta.
Och fariséerna kommo ditut och begynte disputera med honom; de ville sätta honom på prov och begärde av honom något tecken från himmelen.
Då suckade han ur sin andes djup och sade: »Varför begär detta släkte ett tecken?
Sannerligen säger jag eder: Åt detta släkte skall intet tecken givas.»
Så lämnade han dem och steg åter i båten och for över till andra stranden.
Och de hade förgätit att taga med sig bröd; icke mer än ett enda bröd hade de med sig i båten.
Och han bjöd dem och sade: »Sen till, att I tagen eder till vara för fariséernas surdeg och för Herodes' surdeg.»
Då talade de med varandra om att de icke hade bröd med sig.
Men när han märkte detta, sade han till dem: »Varför talen I om att I icke haven bröd med eder?
Fatten och förstån I då ännu ingenting?
Äro edra hjärtan så förstockade?
I haven ju ögon; sen I då icke?
I haven ju öron; hören I då icke?
Och kommen I icke ihåg huru många korgar fulla av stycken I samladen upp, när jag bröt de fem bröden åt de fem tusen?»
De svarade honom: »Tolv.»
»Och när jag bröt de sju bröden åt de fyra tusen, huru många korgar fulla av stycken samladen I då upp?»
De svarade: »Sju.»
Då sade han till dem: »Förstån I då ännu ingenting?»
Därefter kommo de till Betsaida.
Och man förde till honom en som var blind och bad honom att han skulle röra vid denne.
Då tog han den blinde vid handen och ledde honom utanför byn; sedan spottade han på hans ögon och lade händerna på honom och frågade honom: »Ser du något?»
Han såg då upp och svarade: »Jag kan urskilja människorna; jag ser dem gå omkring, men de likna träd.»
Därefter lade han åter händerna på hans ögon, och nu såg han tydligt och var botad och kunde jämväl på långt håll se allting klart.
Och Jesus bjöd honom gå hem och sade: »Gå icke ens in i byn.»
Och Jesus gick med sina lärjungar bort till byarna vid Cesarea Filippi.
På vägen dit frågade han sina lärjungar och sade till dem: »Vem säger folket mig vara?»
De svarade och sade: »Johannes döparen; andra säga dock Elias, andra åter säga: 'Det är en av profeterna.'»
Då frågade han dem: »Vem sägen då I mig vara?»
Petrus svarade och sade till honom: »Du är Messias.»
Då förbjöd han dem strängeligen att för någon säga detta om honom.
Sedan begynte han undervisa dem om att Människosonen måste lida mycket, och att han skulle bliva förkastad av de äldste och översteprästerna och de skriftlärde, och att han skulle bliva dödad, men att han tre dagar därefter skulle uppstå igen.
Och han talade detta i oförtäckta ordalag.
Då tog Petrus honom avsides och begynte ivrigt motsäga honom.
Men han vände sig om, och när han då såg sina lärjungar, talade han strängt till Petrus och sade: »Gå bort, Satan, och stå mig icke i vägen; ty dina tankar äro icke Guds tankar, utan människotankar.»
Och han kallade till sig folket jämte sina lärjungar och sade till dem: »Om någon vill efterfölja mig, så försake han sig själv och tage sitt kors på sig; så följe han mig.
Ty den som vill bevara sitt liv, han skall mista det; men den som mister sitt liv, för min och för evangelii skull, han skall bevara det.
Och vad hjälper det en människa, om hon vinner hela världen, men förlorar sin själ?
Och vad kan en människa giva till lösen för sin själ?
Den som blyges för mig och för mina ord, i detta trolösa och syndiga släkte, för honom skall ock Människosonen blygas, när han kommer i sin Faders härlighet med de heliga änglarna.»
Ytterligare sade han till dem: »Sannerligen säger jag eder: Bland dem som här stå finnas några som icke skola smaka döden, förrän de få se Guds rike vara kommet i sin kraft.»
Sex dagar därefter tog Jesus med sig Petrus och Jakob och Johannes och förde dem ensamma upp på ett högt berg, där de voro allena.
Och hans utseende förvandlades inför dem;
och hans kläder blevo glänsande och mycket vita, så att ingen valkare på jorden kan göra kläder så vita.
Och för dem visade sig Elias jämte Moses, och dessa samtalade med Jesus.
Då tog Petrus till orda och sade till Jesus: »Rabbi, här är oss gott att vara; låt oss göra tre hyddor, åt dig en och åt Moses en och åt Elias en.»
Han visste nämligen icke vad han skulle säga; så stor var deras förskräckelse.
Då kom en sky som överskyggde dem, och ur skyn kom en röst: »Denne är min älskade Son; hören honom.»
Och plötsligt märkte de, när de sågo sig omkring, att där icke mer fanns någon hos dem utom Jesus allena.
Då de sedan gingo ned från berget, bjöd han dem att de icke, förrän Människosonen hade uppstått från de döda, skulle för någon omtala vad de hade sett.
Och de lade märke till det ordet och begynte tala med varandra om vad som kunde menas med att han skulle uppstå från de döda.
Och de frågade honom och sade: »De skriftlärde säga ju att Elias först måste komma?»
Han svarade dem: »Elias måste visserligen först komma och upprätta allt igen.
Men huru kan det då vara skrivet om Människosonen att han skall lida mycket och bliva föraktad?
Dock, jag säger eder att Elias redan har kommit; och de förforo mot honom alldeles såsom de ville, och såsom det var skrivet att det skulle gå honom.»
När de därefter kommo till lärjungarna, sågo de att mycket folk var samlat omkring dem, och att några skriftlärde disputerade med dem.
Och strax då allt folket fick se honom, blevo de mycket häpna och skyndade fram och hälsade honom.
Då frågade han dem: »Varom disputeren I med dem?»
Och en man i folkhopen svarade honom: »Mästare, jag har fört till dig min son, som är besatt av en stum ande.
Och varhelst denne får fatt i honom kastar han omkull honom, och fradgan står gossen om munnen, och han gnisslar med tänderna och bliver såsom livlös.
Nu bad jag dina lärjungar att de skulle driva ut honom, men de förmådde det icke.»
Då svarade han dem och sade: »O du otrogna släkte, huru länge måste jag vara hos eder?
Huru länge måste jag härda ut med eder?
Fören honom till mig.»
Och de förde honom till Jesus.
Och strax då han fick se Jesus, slet och ryckte anden honom, och han föll ned på jorden och vältrade sig, under det att fradgan stod honom om munnen.
Jesus frågade då hans fader: »Huru länge har det varit så med honom?»
Han svarade: »Alltsedan han var ett litet barn;
och det har ofta hänt att han har kastat honom än i elden, än i vattnet, för att förgöra honom.
Men om du förmår något, så förbarma dig över oss och hjälp oss.»
Då sade Jesus till honom: »Om jag förmår, säger du.
Allt förmår den som tror.»
Strax ropade gossens fader och sade: »Jag tror!
Hjälp min otro.»
Men när Jesus såg att folk strömmade tillsammans dit, tilltalade han den orene anden strängt och sade till honom: »Du stumme och döve ande, jag befaller dig: Far ut ur honom, och kom icke mer in i honom.»
Då skriade han och slet och ryckte gossen svårt och for ut; och gossen blev såsom död, så att folket menade att han verkligen var död.
Men Jesus tog honom vid handen och reste upp honom; och han stod då upp.
När Jesus därefter hade kommit inomhus, frågade hans lärjungar honom, då de nu voro allena: »Varför kunde icke vi driva ut honom?»
Han svarade dem: »Detta slag kan icke drivas ut genom något annat än bön och fasta.»
Och de gingo därifrån och vandrade genom Galileen; men han ville icke att någon skulle få veta det.
Han undervisade nämligen sina lärjungar och sade till dem: »Människosonen skall bliva överlämnad i människors händer, och man skall döda honom; men tre dagar efter det att han har blivit dödad skall han uppstå igen.»
Och de förstodo icke vad han sade, men de fruktade att fråga honom.
Och de kommo till Kapernaum.
Och när han hade kommit dit där han bodde, frågade han dem: »Vad var det I samtaladen om på vägen?»
Men de tego, ty de hade på vägen talat med varandra om vilken som vore störst.
Då satte han sig ned och kallade till sig de tolv och sade till dem: »Om någon vill vara den förste, så vare han den siste av alla och allas tjänare.»
Och han tog ett barn och ställde det mitt ibland dem; sedan tog han det upp i famnen och sade till dem:
»Den som tager emot ett sådant barn i mitt namn, han tager emot mig, och den som tager emot mig, han tager icke emot mig, utan honom som har sänt mig.»
Johannes sade till honom: »Mästare, vi sågo huru en man som icke följer oss drev ut onda andar genom ditt namn; och vi ville hindra honom, eftersom han icke följde oss.»
Men Jesus sade: »Hindren honom icke; ty ingen som genom mitt namn har gjort en kraftgärning kan strax därefter tala illa om mig.
Ty den som icke är emot oss, han är för oss.
Ja, den som giver eder en bägare vatten att dricka, därför att I hören Kristus till -- sannerligen säger jag eder: Han skall ingalunda gå miste om sin lön.
Och den som förför en av dessa små som tro, för honom vore det bättre, om en kvarnsten hängdes om hans hals och han kastades i havet.
Om nu din hand är dig till förförelse, så hugg av den.
Det är bättre för dig att ingå i livet lytt, än att hava båda händerna i behåll och komma till Gehenna, till den eld som icke utsläckes.
246520
Och om din fot är dig till förförelse, så hugg av den.
Det är bättre för dig att ingå i livet halt, än att hava båda fötterna i behåll och kastas i Gehenna.
246540
Och om ditt öga är dig till förförelse, så riv ut det.
Det är bättre för dig att ingå i Guds rike enögd, än att hava båda ögonen i behåll och kastas i Gehenna,
där 'deras mask icke dör och elden icke utsläckes'.
Ty var människa måste saltas med eld.
Saltet är en god sak; men om saltet mister sin sälta, varmed skolen I då återställa dess kraft? -- Haven salt i eder och hållen frid inbördes.»
Och han stod upp och begav sig därifrån, genom landet på andra sidan Jordan, till Judeens område.
Och mycket folk församlades åter omkring honom, och åter undervisade han dem, såsom hans sed var.
Då ville några fariséer snärja honom, och de trädde fram och frågade honom om det vore lovligt för en man att skilja sig från sin hustru.
Men han svarade och sade till dem: »Vad har Moses bjudit eder?»
De sade: »Moses tillstadde att en man fick skriva skiljebrev åt sin hustru och så skilja sig från henne.»
Då sade Jesus till dem: »För edra hjärtans hårdhets skull skrev han åt eder detta bud.
Men redan vid världens begynnelse 'gjorde Gud dem till man och kvinna'.
'Fördenskull skall en man övergiva sin fader och sin moder.
Och de tu skola varda ett kött.'
Så äro de icke mer två, utan ett kött.
Vad nu Gud har sammanfogat, det må människan icke åtskilja.»
När de sedan hade kommit hem, frågade hans lärjungar honom åter om detsamma.
Och han svarade dem: »Den som skiljer sig från sin hustru och tager sig en annan hustru, han begår äktenskapsbrott mot henne.
Och om en hustru skiljer sig från sin man och tager sig en annan man, då begår hon äktenskapsbrott.
Och man bar fram barn till honom, för att han skulle röra vid dem; men lärjungarna visade bort dem.
När Jesus såg detta, blev han misslynt och sade till dem: »Låten barnen komma till mig, och förmenen dem det icke; ty Guds rike hör sådana till.
Sannerligen säger jag eder: Den som icke tager emot Guds rike såsom ett barn, han kommer aldrig ditin.»
Och han tog dem upp i famnen och lade händerna på dem och välsignade dem.
När han sedan begav sig åstad för att fortsätta sin väg, skyndade en man fram och föll på knä för honom och frågade honom: »Gode Mästare, vad skall jag göra för att få evigt liv till arvedel?»
Jesus sade till honom: »Varför kallar du mig god?
Ingen är god utom Gud allena.
Buden känner du: 'Du skall icke dräpa', 'Du skall icke begå äktenskapsbrott', 'Du skall icke stjäla', 'Du skall icke bära falskt vittnesbörd', 'Du skall icke undanhålla någon vad honom tillkommer', Hedra din fader och din moder.'»
Då svarade han honom: »Mästare, allt detta har jag hållit från min ungdom.»
Då såg Jesus på honom och fick kärlek till honom och sade till honom: »Ett fattas dig: gå bort och sälj allt vad du äger och giv åt de fattiga; då skall du få en skatt i himmelen.
Och kom sedan och följ mig.»
Men han blev illa till mods vid det talet och gick bedrövad bort, ty han hade många ägodelar.
Då såg Jesus sig omkring och sade till sina lärjungar: »Huru svårt är det icke för dem som hava penningar att komma in i Guds rike!»
Men lärjungarna häpnade vid hans ord.
Då tog Jesus åter till orda och sade till dem: »Ja, mina barn, huru svårt är det icke att komma in i Guds rike!
Det är lättare för en kamel att komma igenom ett nålsöga, än för den som är rik att komma in i Guds rike.»
Då blevo de ännu mer häpna och sade till varandra: »Vem kan då bliva frälst?»
Jesus såg på dem och sade: »För människor är det omöjligt, men icke för Gud, ty för Gud är allting möjligt.»
Då tog Petrus till orda och sade till honom: »Se, vi hava övergivit allt och följt dig.»
Jesus svarade: »Sannerligen säger jag eder: Ingen som för min och evangelii skull har övergivit hus, eller bröder eller systrar, eller moder eller fader, eller barn, eller jordagods,
ingen sådan finnes, som icke skall få hundrafalt igen: redan här i tiden hus, och bröder och systrar, och mödrar och barn, och jordagods, mitt under förföljelser, och i den tillkommande tidsåldern evigt liv.
Men många som äro de första skola bliva de sista, medan de sista bliva de första.»
Och de voro på vägen upp till Jerusalem.
Och Jesus gick före dem, och de gingo där bävande; och de som följde med dem voro uppfyllda av fruktan.
Då tog han åter till sig de tolv och begynte tala till dem om vad som skulle övergå honom:
»Se, vi gå nu upp till Jerusalem, och Människosonen skall bliva överlämnad åt översteprästerna och de skriftlärde, och de skola döma honom till döden och överlämna honom åt hedningarna,
och dessa skola begabba honom och bespotta honom och gissla honom och döda honom; men tre dagar därefter skall han uppstå igen.»
Då trädde Jakob och Johannes, Sebedeus' söner, fram till honom och sade till honom: »Mästare, vi skulle vilja att du läte oss få vad vi nu tänka begära av dig.»
Han frågade dem: »Vad viljen I då att jag skall låta eder få?»
De svarade honom: »Låt den ene av oss i din härlighet få sitta på din högra sida, och den andre på din vänstra.»
Men Jesus sade till dem: »I veten icke vad I begären.
Kunnen I dricka den kalk som jag dricker, eller genomgå det dop som jag genomgår?»
De svarade honom: »Det kunna vi.»
Då sade Jesus till dem: »Ja, den kalk jag dricker skolen I få dricka, och det dop jag genomgår skolen I genomgå,
men platsen på min högra sida och platsen på min vänstra tillkommer det icke mig att bortgiva, utan de skola tillfalla dem för vilka så är bestämt.»
När de tio andra hörde detta, blevo de misslynta på Jakob och Johannes.
Då kallade Jesus dem till sig och sade till dem: »I veten att de som räknas för folkens furstar uppträda mot dem såsom herrar, och att deras mäktige låta dem känna sin myndighet.
Men så är det icke bland eder; utan den som vill bliva störst bland eder, han vare de andras tjänare,
och den som vill vara främst bland eder, han vare allas dräng.
Också Människosonen har ju kommit, icke för att låta tjäna sig, utan för att tjäna och giva sitt liv till lösen för många.»
Och de kommo till Jeriko.
Men när han åter gick ut ifrån Jeriko, följd av sina lärjungar och en ganska stor hop folk, satt där vid vägen en blind tiggare, Bartimeus, Timeus' son.
När denne hörde att det var Jesus från Nasaret, begynte han ropa och säga: »Jesus, Davids son, förbarma dig över mig.»
Och många tillsade honom strängeligen att han skulle tiga; men han ropade ännu mycket mer: »Davids son, förbarma dig över mig.»
Då stannade Jesus och sade: »Kallen honom hit.»
Och de kallade på den blinde och sade till honom: »Var vid gott mod, stå upp; han kallar dig till sig.»
Då kastade han av sig sin mantel och stod upp med hast och kom fram till Jesus.
Och Jesus talade till honom och sade: »Vad vill du att jag skall göra dig?»
Den blinde svarade honom: »Rabbuni, låt mig få min syn.»
Jesus sade till honom: »Gå; din tro har hjälpt dig.»
Och strax fick han sin syn och följde honom på vägen.
När de nu nalkades Jerusalem och voro nära Betfage och Betania vid Oljeberget, sände han åstad två av sina lärjungar
och sade till dem: »Gån in i byn som ligger mitt framför eder, så skolen I, strax då I kommen ditin, finna en åsnefåle stå där bunden, som ännu ingen människa har suttit på; lösen den och fören den hit.
Och om någon frågar eder varför I gören detta, så skolen I svara: 'Herren behöver den, men han skall strax sända den tillbaka hit.»
Då gingo de åstad och funno en åsnefåle stå där bunden utanför en port vid vägen, och de löste den.
Och några som stodo där bredvid sade till dem: »Vad gören I?
Varför lösen I fålen?»
Men de svarade dem såsom Jesus hade bjudit.
Då lät man dem vara.
Och de förde fålen till Jesus och lade sina mantlar på den, och han satte sig upp på den.
Och många bredde ut sina mantlar på vägen, andra åter skuro av kvistar och löv på fälten och strödde på vägen.
Och de som gingo före och de som följde efter ropade: »Hosianna!
Välsignad vare han som kommer, i Herrens namn.
Välsignat vare vår fader Davids rike, som nu kommer.
Hosianna i höjden!»
Så drog han in i Jerusalem och kom in i helgedomen; och när han hade sett sig omkring överallt och det redan var sent på dagen, gick han med de tolv ut till Betania.
När de dagen därefter voro på väg tillbaka från Betania, blev han hungrig.
Och då han på avstånd fick se ett fikonträd som hade löv, gick han dit för att se om han till äventyrs skulle finna något därpå; men när han kom fram till det, fann han intet annat än löv, det var icke då fikonens tid.
Då talade han och sade till trädet: »Aldrig någonsin mer äte någon frukt av dig.»
Och hans lärjungar hörde detta.
När de sedan kommo fram till Jerusalem, gick han in i helgedomen och begynte driva ut dem som sålde och köpte i helgedomen.
Och han stötte omkull växlarnas bord och duvomånglarnas säten;
han tillstadde icke heller att man bar någonting genom helgedomen.
Och han undervisade dem och sade: »Det är ju skrivet: 'Mitt hus skall kallas ett bönehus för alla folk.'
Men I haven gjort det till en rövarkula.»
Då översteprästerna och de skriftlärde fingo höra härom, sökte de efter tillfälle att förgöra honom; ty de fruktade för honom, eftersom allt folket häpnade över hans undervisning.
När det blev afton, begåvo de sig ut ur staden.
Men då de nu på morgonen åter gingo där fram, fingo de se fikonträdet vara förtorkat ända från roten.
Då kom Petrus ihåg vad som hade skett och sade till honom: »Rabbi, se, fikonträdet som du förbannade är förtorkat.»
Jesus svarade och sade till dem: »Haven tro på Gud.
Sannerligen säger jag eder: Om någon säger till detta berg: 'Häv dig upp, och kasta dig i havet' och därvid icke tvivlar i sitt hjärta, utan tror att det han säger skall ske, då skall det ske honom så.
Därför säger jag eder: Allt vad I bedjen om och begären, tron att det är eder givet; och det skall ske eder så.
Och när I stån och bedjen, så förlåten, om I haven något emot någon, för att också eder Fader, som är i himmelen, må förlåta eder edra försyndelser.»
247360
Så kommo de åter till Jerusalem.
Och medan han gick omkring i helgedomen, kommo översteprästerna och de skriftlärde och de äldste fram till honom;
och de sade till honom: »Med vad myndighet gör du detta?
Och vem har givit dig myndighet att göra detta?»
Jesus svarade dem: »Jag vill ställa en fråga till eder; svaren mig på den, så skall ock jag säga eder med vad myndighet jag gör detta.
Johannes' döpelse, var den från himmelen eller från människor?
Svaren mig härpå.»
Då överlade de med varandra och sade: »Om vi svara: 'Från himmelen', så frågar han: 'Varför trodden I honom då icke?'
Eller skola vi svara: 'Från människor'?» -- det vågade de icke av fruktan för folket, ty alla höllo före att Johannes verkligen var en profet.
De svarade alltså Jesus och sade: »Vi veta det icke.»
Då sade Jesus till dem: »Så säger icke heller jag eder med vad myndighet jag gör detta.»
Och han begynte tala till dem i liknelser: »En man planterade en vingård och satte stängsel däromkring och högg ut ett presskar och byggde ett vakttorn; därefter lejde han ut den åt vingårdsmän och for utrikes.
När sedan rätta tiden var inne, sände han en tjänare till vingårdsmännen, för att denne av vingårdsmännen skulle uppbära någon del av vingårdens frukt.
Men de togo fatt på honom och misshandlade honom och läto honom gå tomhänt tillbaka.
Åter sände han till dem en annan tjänare.
Honom slogo de i huvudet och skymfade.
Sedan sände han åstad ännu en annan, men denne dräpte de.
Likaså gjorde de med många andra: somliga misshandlade de, och andra dräpte de.
Nu hade han ock en enda son, vilken han älskade.
Honom sände han slutligen åstad till dem, ty han tänkte: 'De skola väl hava försyn för min son.'
Men vingårdsmännen sade till varandra: 'Denne är arvingen; kom, låt oss dräpa honom, så bliver arvet vårt.'
Och de togo fatt på honom och dräpte honom och kastade honom ut ur vingården. --
Vad skall nu vingårdens herre göra?
Jo, han skall komma och förgöra vingårdsmännen och lämna vingården åt andra.
Haven I icke läst detta skriftens ord: 'Den sten som byggningsmännen förkastade, den har blivit en hörnsten;
av Herren har den blivit detta, och underbar är den i våra ögon'?»
De hade nu gärna velat gripa honom, men de fruktade för folket; ty de förstodo att det var om dem som han hade talat i denna liknelse.
Så läto de honom vara och gingo sin väg.
Därefter sände de till honom några fariséer och herodianer, för att dessa skulle fånga honom genom något hans ord.
Dessa kommo nu och sade till honom: »Mästare, vi veta att du är sannfärdig och icke frågar efter någon, ty du ser icke till personen, utan lär om Guds väg vad sant är.
Är det lovligt att giva kejsaren skatt, eller är det icke lovligt?
Skola vi giva skatt, eller icke giva?»
Men han förstod deras skrymteri och sade till dem: »Varför söken I att snärja mig?
Tagen hit en penning, så att jag får se den.»
Då lämnade de fram en sådan.
Därefter frågade han dem: »Vems bild och överskrift är detta?»
De svarade honom: »Kejsarens.»
Då sade Jesus till dem: »Så given kejsaren vad kejsaren tillhör, och Gud vad Gud tillhör.»
Och de förundrade sig högeligen över honom.
Sedan kommo till honom några av sadducéerna, vilka mena att det icke gives någon uppståndelse.
Dessa frågade honom och sade:
»Mästare, Moses har givit oss den föreskriften, att om någon har en broder som dör, och som efterlämnar hustru, men icke lämnar barn efter sig, så skall han taga sin broders hustru till äkta och skaffa avkomma åt sin broder.
Nu voro här sju bröder.
Den förste tog sig en hustru, men dog utan att lämna någon avkomma efter sig.
Då tog den andre i ordningen henne, men också han dog utan att lämna någon avkomma efter sig; sammalunda den tredje.
Så skedde med alla sju: ingen av dem lämnade någon avkomma efter sig.
Sist av alla dog ock hustrun.
Vilken av dem skall nu vid uppståndelsen, när de uppstå, få henne till hustru?
De hade ju alla sju tagit henne till hustru.»
Jesus svarade dem: »Visar icke eder fråga att I faren vilse och varken förstån skrifterna, ej heller Guds kraft?
Efter uppståndelsen från de döda taga män sig icke hustrur, ej heller givas hustrur åt män, utan de äro då såsom änglarna i himmelen.
Men vad nu det angår, att de döda uppstå, haven I icke läst i Moses' bok, på det ställe där det talas om törnbusken, huru Gud sade till honom så: 'Jag är Abrahams Gud och Isaks Gud och Jakobs Gud'?
Han är en Gud icke för döda, utan för levande.
I faren mycket vilse.»
Då trädde en av de skriftlärde fram, en som hade hört deras ordskifte och förstått att han hade svarat dem väl.
Denne frågade honom: »Vilket är det förnämsta av alla buden?»
Jesus svarade: »Det förnämsta är detta: 'Hör, Israel!
Herren, vår Gud, Herren är en.
Och du skall älska Herren, din Gud, av allt ditt hjärta och av all din själ och av allt ditt förstånd och av all din kraft.'
Därnäst kommer detta: 'Du skall älska din nästa såsom dig själv.'
Intet annat bud är större än dessa.»
Då svarade den skriftlärde honom: »Mästare, du har i sanning rätt i vad du säger, att han är en, och att ingen annan är än han.
Och att älska honom av allt sitt hjärta och av allt sitt förstånd och av all sin kraft och att älska sin nästa såsom sig själv, det är 'förmer än alla brännoffer och slaktoffer'.»
Då nu Jesus märkte att han hade svarat förståndigt, sade han till honom: »Du är icke långt ifrån Guds rike.»
Sedan dristade sig ingen att vidare ställa någon fråga på honom.
Medan Jesus undervisade i helgedomen, framställde han denna fråga: »Huru kunna de skriftlärde säga att Messias är Davids son?
David själv har ju sagt genom den helige Andes ingivelse: 'Herren sade till min herre: Sätt dig på min högra sida, till dess jag har lagt dina fiender dig till en fotapall.'
Så kallar nu David själv honom 'herre'; huru kan han då vara hans son?»
Och folkskarorna hörde honom gärna.
Och han undervisade dem och sade till dem: »Tagen eder till vara för de skriftlärde, som gärna gå omkring i fotsida kläder och gärna vilja bliva hälsade på torgen
och gärna sitta främst i synagogorna och på de främsta platserna vid gästabuden --
detta under det att de utsuga änkors hus, medan de för syns skull hålla långa böner.
De skola få en dess hårdare dom.»
Och han satte sig mitt emot offerkistorna och såg huru folket lade ned penningar i offerkistorna.
Och många rika lade dit mycket.
Men en fattig änka kom och lade ned två skärvar, det är ett öre.
Då kallade han sina lärjungar till sig och sade till dem: »Sannerligen säger jag eder: Denna fattiga änka lade dit mer än alla de andra som lade något i offerkistorna.
Ty dessa lade alla dit av sitt överflöd, men hon lade dit av sitt armod allt vad hon hade, så mycket som fanns i hennes ägo.»
Då han nu gick ut ur helgedomen, sade en av hans lärjungar till honom: »Mästare, se hurudana stenar och hurudana byggnader!»
Jesus svarade honom: »Ja, du ser nu dessa stora byggnader; men här skall förvisso icke lämnas sten på sten; allt skall bliva nedbrutet.»
När han sedan satt på Oljeberget, mitt emot helgedomen, frågade honom Petrus och Jakob och Johannes och Andreas, då de voro allena:
»Säg oss när detta skall ske, och vad som bliver tecknet till att tiden är inne, då allt detta skall gå i fullbordan.»
Då begynte Jesus tala till dem och sade: »Sen till, att ingen förvillar eder.
Många skola komma under mitt namn och säga: 'Det är jag' och skola förvilla många.
Men när I fån höra krigslarm och rykten om krig, så förloren icke besinningen; sådant måste komma, men därmed är ännu icke änden inne.
Ja, folk skall resa sig upp mot folk och rike mot rike, och det skall bliva jordbävningar på den ena orten efter den andra, och hungersnöd skall uppstå; detta är begynnelsen till 'födslovåndorna'.
Men tagen I eder till vara.
Man skall då draga eder inför domstolar, och I skolen bliva gisslade i synagogor och ställas fram inför landshövdingar och konungar, för min skull, till ett vittnesbörd för dem.
Men evangelium måste först bliva predikat för alla folk.
När man nu för eder åstad och drager eder inför rätta, så gören eder icke förut bekymmer om vad I skolen tala; utan vad som bliver eder givet i den stunden, det mån I tala.
Ty det är icke I som skolen tala, utan den helige Ande.
Och den ene brodern skall då överlämna den andre till att dödas, ja ock fadern sitt barn; och barn skola sätta sig upp mot sina föräldrar och skola döda dem.
Och I skolen bliva hatade av alla, för mitt namns skull.
Men den som är ståndaktig intill änden, han skall bliva frälst.
Men när I fån se 'förödelsens styggelse' stå där han icke borde stå -- den som läser detta, han give akt därpå -- då må de som äro i Judeen fly bort till bergen,
och den som är på taket må icke stiga ned och gå in för att hämta något ur sitt hus,
och den som är ute på marken må icke vända tillbaka för att hämta sin mantel.
Och ve de som äro havande, eller som giva di på den tiden!
Men bedjen att det icke må ske om vintern.
Ty den tiden skall bliva 'en tid av vedermöda, så svår att dess like icke har förekommit allt ifrån världens begynnelse, från den tid då Gud skapade världen, intill nu', ej heller någonsin skall förekomma.
Och om Herren icke förkortade den tiden, så skulle intet kött bliva frälst; men för de utvaldas skull, för de människors skull, som han har utvalt, har han förkortat den tiden.
Och om någon då säger till eder: 'Se här är Messias', eller: 'Se där är han', så tron det icke.
Ty människor som falskeligen säga sig vara Messias skola uppstå, så ock falska profeter, och de skola göra tecken och under, för att, om möjligt, förvilla de utvalda.
Men tagen I eder till vara.
Jag har nu sagt eder allt förut.
Men på den tiden, efter den vedermödan, skall solen förmörkas och månen upphöra att giva sitt sken,
och stjärnorna skola falla ifrån himmelen, och makterna i himmelen skola bäva.
Och då skall man få se 'Människosonen komma i skyarna' med stor makt och härlighet.
Och han skall då sända ut sina änglar och församla sina utvalda från de fyra väderstrecken, från jordens ända till himmelens ända.
Ifrån fikonträdet mån I här hämta en liknelse.
När dess kvistar begynna att få save och löven spricka ut, då veten I att sommaren är nära.
Likaså, när I sen detta ske, då kunnen I ock veta att han är nära och står för dörren.
Sannerligen säger jag eder: Detta släkte skall icke förgås, förrän allt detta sker.
Himmel och jord skola förgås, men mina ord skola icke förgås.
Men om den dagen och den stunden vet ingen något, icke änglarna i himmelen, icke ens Sonen -- ingen utom Fadern.
Tagen eder till vara, vaken; ty I veten icke när tiden är inne.
Såsom när en man reser utrikes och lämnar sitt hus och giver sina tjänare makt och myndighet däröver, åt var och en hans särskilda syssla, och därvid ock bjuder portvaktaren att vaka.
likaså bjuder jag eder: Vaken; ty I veten icke när husets herre kommer, om han kommer på aftonen eller vid midnattstiden eller i hanegället eller på morgonen;
vaken, så att han icke finner eder sovande, när han oförtänkt kommer.
Men vad jag säger till eder, det säger jag till alla: Vaken!»
Två dagar därefter var det påsk och det osyrade brödets högtid.
Och översteprästerna och de skriftlärde sökte efter tillfälle att gripa honom med list och döda honom.
De sade nämligen: »Icke under högtiden, för att ej oroligheter skola uppstå bland folket.»
Men när han var i Betania, i Simon den spetälskes hus, och där låg till bords, kom en kvinna som hade med sig en alabasterflaska med smörjelse av dyrbar äkta nardus.
Och hon bröt sönder flaskan och göt ut smörjelsen över hans huvud.
Några som voro där blevo då misslynta och sade till varandra: »Varför skulle denna smörjelse förspillas?
Man hade ju kunnat sälja den för mer än tre hundra silverpenningar och giva dessa åt de fattiga.»
Och de talade hårda ord till henne.
Men Jesus sade: »Låten henne vara.
Varför oroen I henne?
Det är en god gärning som hon har gjort mot mig.
De fattiga haven I ju alltid ibland eder, och närhelst I viljen kunnen I göra dem gott, men mig haven I icke alltid.
Vad hon kunde, det gjorde hon.
Hon har i förväg smort min kropp såsom en tillredelse till min begravning.
Och sannerligen säger jag eder: Varhelst i hela världen evangelium bliver predikat, där skall ock det som hon nu har gjort bliva omtalat, henne till åminnelse.»
Och Judas Iskariot, han som var en av de tolv, gick bort till översteprästerna och ville förråda honom åt dem.
När de hörde detta, blevo de glada och lovade att giva honom en summa penningar.
Sedan sökte han efter tillfälle att förråda honom, då lägligt var.
På första dagen i det osyrade brödets högtid, när man slaktade påskalammet, sade hans lärjungar till honom: »Vart vill du att vi skola gå och reda till, så att du kan äta påskalammet?»
Då sände han åstad två av sina lärjungar och sade till dem: »Gån in i staden; där skolen I möta en man som bär en kruka vatten.
Följen honom.
Och sägen till husbonden i det hus där han går in: 'Mästaren frågar: Var finnes härbärget där jag skall äta påskalammet med mina lärjungar?'
Då skall han visa eder en stor sal i övre våningen, tillredd och ordnad för måltid; reden till åt oss där.»
Och lärjungarna begåvo sig i väg och kommo in i staden och funno det så som han hade sagt dem; och de redde till påskalammet.
När det sedan hade blivit afton, kom han dit med de tolv.
Och medan de lågo till bords och åto, sade Jesus: »Sannerligen säger jag eder: En av eder skall förråda mig, 'den som äter med mig'.»
Då begynte de bedrövas och fråga honom, den ene efter den andre: »Icke är det väl jag?»
Och han sade till dem: »Det är en av de tolv, den som jämte mig doppar i fatet.
Ja, Människosonen skall gå bort, såsom det är skrivet om honom; men ve den människa genom vilken Människosonen bliver förrådd!
Det hade varit bättre för den människan, om hon icke hade blivit född.»
Medan de nu åto, tog han ett bröd och välsignade det och bröt det och gav åt dem och sade: »Tagen detta; detta är min lekamen.»
Och han tog en kalk och tackade Gud ock gav åt dem; och de drucko alla därav.
Och han sade till dem: »Detta är mitt blod, förbundsblodet, som varder utgjutet för många.
Sannerligen säger jag eder: Jag skall icke mer dricka av det som kommer från vinträd, förrän på den dag då jag dricker det nytt i Guds rike.»
När de sedan hade sjungit lovsången, gingo de ut till Oljeberget.
Då sade Jesus till dem: »I skolen alla komma på fall; ty det är skrivet: 'Jag skall slå herden, och fåren skola förskingras.'
Men efter min uppståndelse skall jag före eder gå till Galileen.»
Då svarade Petrus honom: »Om än alla andra komma på fall, så skall dock jag det icke.»
Jesus sade till honom: »Sannerligen säger jag dig: Redan i denna natt, förrän hanen har galit två gånger, skall du tre gånger förneka mig.»
Då försäkrade han ännu ivrigare: »Om jag än måste dö med dig, så skall jag dock icke förneka dig.»
Sammalunda sade ock alla de andra.
Och de kommo till ett ställe som kallades Getsemane.
Då sade han till sina lärjungar: »Bliven kvar här, medan jag beder.»
Och han tog med sig Petrus och Jakob och Johannes; och han begynte bäva och ängslas.
Och han sade till dem: »Min själ är djupt bedrövad, ända till döds; stannen kvar här och vaken.»
Därefter gick han litet längre bort och föll ned på jorden och bad, att om möjligt vore, den stunden skulle bliva honom besparad.
Och han sade: »Abba, Fader, allt är möjligt för dig.
Tag denna kalk ifrån mig.
Dock icke vad jag vill, utan vad du vill!»
Sedan kom han tillbaka och fann dem sovande.
Då sade han till Petrus: »Simon, sover du?
Förmådde du då icke vaka en kort stund?
Vaken, och bedjen att I icke mån komma i frestelse.
Anden är villig, men köttet är svagt.»
Och han gick åter bort och bad och sade samma ord.
När han sedan kom tillbaka, fann han dem åter sovande, ty deras ögon voro förtyngda.
Och de visste icke vad de skulle svara honom.
För tredje gången kom han tillbaka och sade då till dem: »Ja, I soven ännu alltjämt och vilen eder!
Det är nog.
Stunden är kommen.
Människosonen skall nu bliva överlämnad i syndarnas händer.
Stån upp, låt oss gå; se, den som förråder mig är nära.»
Och i detsamma, medan han ännu talade, kom Judas, en av de tolv, och jämte honom en folkskara med svärd och stavar, utsänd från översteprästerna och de skriftlärde och de äldste.
Men förrädaren hade kommit överens med dem om ett tecken och sagt: »Den som jag kysser, den är det; honom skolen I gripa och föra bort under säker bevakning.»
Och när han nu kom dit, trädde han strax fram till honom och sade: »Rabbi!» och kysste honom häftigt.
Då grepo de Jesus och togo honom fången.
Men en av dem som stodo där bredvid drog sitt svärd och högg till översteprästens tjänare och högg så av honom örat.
Och Jesus talade till dem och sade: »Såsom mot en rövare haven I gått ut med svärd och stavar för att fasttaga mig.
Var dag har jag varit ibland eder i helgedomen och undervisat, utan att I haven gripit mig.
Men skrifterna skulle ju fullbordas.»
Då övergåvo de honom alla och flydde.
Och bland dem som hade följt med honom var en ung man, höljd i ett linnekläde, som var kastat över blotta kroppen; honom grepo de.
Men han lämnade linneklädet kvar och flydde undan naken.
Så förde de nu Jesus bort till översteprästen, och där församlade sig alla översteprästerna och de äldste och de skriftlärde.
Och Petrus följde honom på avstånd ända in på översteprästens gård; där satt han sedan tillsammans med tjänarna och värmde sig vid elden.
Och översteprästerna och hela Stora rådet sökte efter något vittnesbörd mot Jesus, för att kunna döda honom; men de funno intet.
Ty väl vittnade många falskt mot honom, men vittnesbörden stämde icke överens.
Och några stodo upp och vittnade falskt mot honom och sade:
»Vi hava själva hört honom säga: 'Jag skall bryta ned detta tempel, som är gjort med händer, och skall sedan på tre dagar bygga upp ett annat, som icke är gjort med händer.'»
Men icke ens i det stycket stämde deras vittnesbörd överens.
Då stod översteprästen upp ibland dem och frågade Jesus och sade: »Svarar du intet?
Huru är det med det som dessa vittna mot dig?»
Men han teg och svarade intet.
Åter frågade översteprästen honom och sade till honom: »Är du Messias, den Högtlovades Son?»
Jesus svarade: »Jag är det.
Och I skolen få se Människosonen sitta på Maktens högra sida och komma med himmelens skyar.»
Då rev översteprästen sönder sina kläder och sade: »Vad behöva vi mer några vittnen?
I hörden hädelsen.
Vad synes eder?»
Då dömde de alla honom skyldig till döden.
Och några begynte spotta på honom; och sedan de hade höljt över hans ansikte, slogo de honom på kinderna med knytnävarna och sade till honom: »Profetera.»
Också rättstjänarna slogo honom på kinderna.
Medan nu Petrus befann sig därnere på gården, kom en av översteprästens tjänstekvinnor dit.
Och när hon fick se Petrus, där han satt och värmde sig, såg hon på honom och sade: »Också du var med nasaréen, denne Jesus.»
Men han nekade och sade: »Jag varken vet eller förstår vad du menar.»
Sedan gick han ut på den yttre gården.
När tjänstekvinnan då fick se honom där, begynte hon åter säga till dem som stodo bredvid: »Denne är en av dem.»
Då nekade han åter.
Litet därefter sade återigen de som stodo där bredvid till Petrus: »Förvisso är du en av dem; du är ju också en galilé.»
Då begynte han förbanna sig och svärja: »Jag känner icke den man som I talen om.»
Och i detsamma gol hanen för andra gången.
Då kom Petrus ihåg Jesu ord, huru han hade sagt till honom: »Förrän hanen har galit två gånger, skall du tre gånger förneka mig.»
Och han brast ut i gråt.
Sedan nu översteprästerna, tillsammans med de äldste och de skriftlärde, hela Stora rådet, på morgonen hade fattat sitt beslut, läto de strax binda Jesus och förde honom bort och överlämnade honom åt Pilatus.
Då frågade Pilatus honom: »Är du judarnas konung?»
Han svarade honom och sade: »Du säger det själv.»
Och översteprästerna framställde många anklagelser mot honom.
Pilatus frågade honom då åter och sade: »Svarar du intet?
Du hör ju huru mycket det är som de anklaga dig för.»
Men Jesus svarade intet mer, så att Pilatus förundrade sig.
Nu plägade han vid högtiden giva dem en fånge lös, den som de begärde.
Och där fanns då en man, han som kallades Barabbas, vilken satt fängslad jämte de andra som hade gjort upplopp och under upploppet begått dråp.
Folket kom ditupp och begynte begära att han skulle göra åt dem såsom han plägade göra.
Pilatus svarade dem och sade: »Viljen I att jag skall giva eder 'judarnas konung' lös?»
Han förstod nämligen att det var av avund som översteprästerna hade dragit Jesus inför rätta.
Men översteprästerna uppeggade folket till att begära att han hellre skulle giva dem Barabbas lös.
När alltså Pilatus åter tog till orda och frågade dem: »Vad skall jag då göra med den som I kallen 'judarnas konung'?»,
så skriade de åter: »Korsfäst honom!»
Men Pilatus frågade dem: »Vad ont har han då gjort?»
Då skriade de ännu ivrigare: »Korsfäst honom!»
Och eftersom Pilatus ville göra folket till viljes, gav han dem Barabbas lös; men Jesus lät han gissla och utlämnade honom sedan till att korsfästas.
Och krigsmännen förde honom in i palatset, eller pretoriet, och kallade tillhopa hela den romerska vakten.
Och de klädde på honom en purpurfärgad mantel och vredo samman en krona av törnen och satte den på honom.
Sedan begynte de hälsa honom: »Hell dig, judarnas konung!»
Och de slogo honom i huvudet med ett rör och spottade på honom; därvid böjde de knä och gåvo honom sin hyllning.
Och när de hade begabbat honom, klädde de av honom den purpurfärgade manteln och satte på honom hans egna kläder och förde honom ut för att korsfästa honom.
Och en man som kom utifrån marken gick där fram, Simon från Cyrene, Alexanders och Rufus' fader; honom tvingade de att gå med och bära hans kors.
Och de förde honom till Golgataplatsen (det betyder huvudskalleplatsen).
Och de räckte honom vin, blandat med myrra, men han tog icke emot det.
Och de korsfäste honom och delade sedan hans kläder mellan sig, genom att kasta lott om vad var och en skulle få.
Och det var vid tredje timmen som de korsfäste honom.
Och den överskrift som man hade satt upp över honom, för att angiva vad han var anklagad för, hade denna lydelse: »Judarnas konung.»
Och de korsfäste med honom två rövare, den ene på hans högra sida och den andre på hans vänstra.
249240
Och de som gingo där förbi bespottade honom och skakade huvudet och sade: »Tvi dig, du som 'bryter ned templet och bygger upp det igen inom tre dagar'!
Hjälp dig nu själv, och stig ned från korset.»
Sammalunda talade ock översteprästerna, jämte de skriftlärde, begabbande ord med varandra och sade: »Andra har han hjälpt; sig själv kan han icke hjälpa.
Han som är Messias, Israels konung, han stige nu ned från korset, så att vi få se det och tro.»
Också de män som voro korsfästa med honom smädade honom.
Men vid sjätte timmen kom över hela landet ett mörker, som varade ända till nionde timmen.
Och vid nionde timmen ropade Jesus med hög röst: »Eloi, Eloi, lema sabaktani?»; det betyder: »Min Gud, min Gud, varför har du övergivit mig?»
Då några av dem som stodo där bredvid hörde detta, sade de: »Hör, han kallar på Elias.»
Men en av dem skyndade fram och fyllde en svamp med ättikvin och satte den på ett rör och gav honom att dricka, i det han sade: »Låt oss se om Elias kommer och tager honom ned.»
Men Jesus ropade med hög röst och gav upp andan.
Då rämnade förlåten i templet i två stycken, uppifrån och ända ned.
Men när hövitsmannen, som stod där mitt emot honom, såg att han på sådant sätt gav upp andan, sade han: »Förvisso var denne man Guds Son.»
Också några kvinnor stodo där på avstånd och sågo vad som skedde.
Bland dessa voro jämväl Maria från Magdala och den Maria som var Jakob den yngres och Joses' moder, så ock Salome
-- vilka hade följt honom och tjänat honom, medan han var i Galileen -- därtill många andra kvinnor, de som med honom hade vandrat upp till Jerusalem.
Det var nu tillredelsedag (det är dagen före sabbaten), och det hade blivit afton.
Josef från Arimatea, en ansedd rådsherre och en av dem som väntade på Guds rike, tog därför nu mod till sig och gick in till Pilatus och utbad sig att få Jesu kropp.
Då förundrade sig Pilatus över att Jesus redan skulle vara död, och han kallade till sig hövitsmannen och frågade honom om det var länge sedan han hade dött.
Och när han av hövitsmannen hade fått veta huru det var, skänkte han åt Josef hans döda kropp.
Denne köpte då en linneduk och tog honom ned och svepte honom i linneduken och lade honom i en grav som var uthuggen i en klippa; sedan vältrade han en sten för ingången till graven.
Men Maria från Magdala och den Maria som var Joses' moder sågo var han lades.
Och när sabbaten var förliden, köpte Maria från Magdala och den Maria som var Jakobs moder och Salome välluktande kryddor, för att sedan gå åstad och smörja honom.
Och bittida om morgonen på första veckodagen kommo de till graven, redan vid soluppgången.
Och de sade till varandra: »Vem skall åt oss vältra bort stenen från ingången till graven?»
Men när de sågo upp, fingo de se att stenen redan var bortvältrad.
Den var nämligen mycket stor.
Och när de hade kommit in i graven, fingo de se en ung man sitta där på högra sidan, klädd i en vit fotsid klädnad; och de blevo förskräckta.
Men han sade till dem: »Varen icke förskräckta.
I söken Jesus från Nasaret, den korsfäste.
Han är uppstånden, han är icke här.
Se där är platsen där de lade honom.
Men gån bort och sägen till hans lärjungar, och särskilt till Petrus: 'Han skall före eder gå till Galileen; där skolen I få se honom, såsom han bar sagt eder.'»
Då gingo de ut och flydde bort ifrån graven, ty bävan och bestörtning hade kommit över dem.
Och i sin fruktan sade de intet till någon.
n efter sin uppståndelse visade han sig på första veckodagens morgon först för Maria från Magdala, ur vilken han hade drivit ut sju onda andar.
Hon gick då och omtalade det för dem som hade följt med honom, och som nu sörjde och gräto.
Men när dessa hörde sägas att han levde och hade blivit sedd av henne, trodde de det icke.
Därefter uppenbarade han sig i en annan skepnad för två av dem, medan de voro stadda på vandring utåt landsbygden.
Också dessa gingo bort och omtalade det för de andra; men icke heller dem trodde man.
Sedan uppenbarade han sig också för de elva, när de lågo till bords; och han förebrådde dem då deras otro och deras hjärtans hårdhet, i det att de icke hade trott dem som hade sett honom vara uppstånden.
Och han sade till dem: »Gån ut i hela världen och prediken evangelium för allt skapat.
Den som tror och bliver döpt, han skall bliva frälst; men den som icke tror, han skall bliva fördömd.
Och dessa tecken skola åtfölja dem som tro: genom mitt namn skola de driva ut onda andar, de skola tala nya tungomål,
ormar skola de taga i händerna, och om de dricka något dödande gift, så skall det alls icke skada dem; på sjuka skola de lägga händerna, och de skola då bliva friska.»
Därefter, sedan Herren Jesus hade talat med dem, blev han upptagen i himmelen och satte sig på Guds högra sida.
Men de gingo ut och predikade allestädes.
Och Herren verkade med dem och stadfäste ordet genom de tecken som åtföljde det.]
Alldenstund många andra hava företagit sig att om de händelser, som bland oss hava timat, avfatta berättelser,
i enlighet med vad som har blivit oss meddelat av dem som själva voro åsyna vittnen och ordets tjänare,
så har ock jag, sedan jag grundligt har efterforskat allt ända ifrån begynnelsen, beslutit mig för att i följd och ordning skriva därom till dig, ädle Teofilus,
så att du kan inse huru tillförlitliga de stycken äro, i vilka du har blivit undervisad.
På den tid då Herodes var konung över Judeen levde en präst vid namn Sakarias, av Abias' »dagsavdelning».
Denne hade till hustru en av Arons döttrar som hette Elisabet.
De voro båda rättfärdiga inför Gud och vandrade ostraffligt efter alla Herrens bud och stadgar.
Men de hade inga barn, ty Elisabet var ofruktsam; och båda voro de komna till hög ålder.
Medan han nu en gång, när ordningen kom till hans avdelning, gjorde prästerlig tjänst inför Gud,
hände det sig, vid den övliga lottningen om de prästerliga sysslorna, att det tillföll honom att gå in i Herrens tempel och tända rökelsen.
Och hela menigheten stod utanför och bad, medan rökoffret förrättades.
Då visade sig för honom en Herrens ängel, stående på högra sidan om rökelsealtaret.
Och när Sakarias såg honom, blev han förskräckt, och fruktan föll över honom.
Men ängeln sade till honom: »Frukta icke, Sakarias; ty din bön är hörd, och din hustru Elisabet skall föda dig en son, och honom skall du giva namnet Johannes.
Och han skall bliva dig till glädje och fröjd, och många skola glädja sig över hans födelse.
Ty han skall bliva stor inför Herren.
Vin och starka drycker skall han icke dricka, och redan i sin moders liv skall han bliva uppfylld av helig ande.
Och många av Israels barn skall han omvända till Herren, deras Gud.
Han skall gå framför honom i Elias' ande och kraft, för att 'vända fädernas hjärtan till barnen' och omvända de ohörsamma till de rättfärdigas sinnelag, så att han skaffar åt Herren ett välberett folk.»
Då sade Sakarias till ängeln: »Varav skall jag veta detta?
Jag är ju själv gammal, och min hustru är kommen till hög ålder.»
Ängeln svarade och sade till honom: »Jag är Gabriel, som står inför Gud, och jag är utsänd för att tala till dig och förkunna dig detta glada budskap.
Och se, ända till den dag då detta sker skall du vara mållös och icke kunna tala, därför att du icke trodde mina ord, vilka dock i sin tid skola fullbordas.»
Och folket stod och väntade på Sakarias och förundrade sig över att han så länge dröjde i templet;
och när han kom ut, kunde han icke tala till dem.
Då förstodo de att han hade sett någon syn i templet.
Och han tecknade åt dem och förblev stum.
Och när tiden för hans tjänstgöring hade gått till ända, begav han sig hem.
Men efter den tiden blev hans hustru Elisabet havande och höll sig dold i fem månader;
och hon sade: »Så har Herren gjort med mig nu, då han har sett till min smälek bland människorna, för att borttaga den.»
I sjätte månaden blev ängeln Gabriel sänd av Gud till en stad i Galileen som hette Nasaret,
till en jungfru som var trolovad med en man vid namn Josef, av Davids hus; och jungfruns namn var Maria.
Och ängeln kom in till henne och sade: »Hell dig, du högtbenådade!
Herren är med dig.»
Men hon blev mycket förskräckt vid hans ord och tänkte på vad denna hälsning månde innebära.
Då sade ängeln till henne: »Frukta icke, Maria; ty du har funnit nåd för Gud.
Se, du skall bliva havande och föda en son, och honom skall du giva namnet Jesus.
Han skall bliva stor och kallas den Högstes Son, och Herren Gud skall giva honom hans fader Davids tron.
Och han skall vara konung över Jakobs hus till evig tid, och på hans rike skall ingen ände vara.»
Då sade Maria till ängeln: »Huru skall detta ske?
Jag vet ju icke av någon man.»
Ängeln svarade och sade till henne: »Helig ande skall komma över dig, och kraft från den Högste skall överskygga dig; därför skall ock det heliga som varder fött kallas Guds Son.
Och se, jämväl din fränka Elisabet har blivit havande och skall föda en son, nu på sin ålderdom; och detta är sjätte månaden för henne, som säges vara ofruktsam.
Ty för Gud kan intet vara omöjligt.»
Då sade Maria: »Se, jag är Herrens tjänarinna; ske mig såsom du har sagt.»
Och ängeln lämnade henne.
En av de närmaste dagarna stod Maria upp och begav sig skyndsamt till en stad i Judeen, uppe i bergsbygden.
Och hon trädde in i Sakarias' hus och hälsade Elisabet.
När då Elisabet hörde Marias hälsning, spratt barnet till i hennes liv; och Elisabet blev fylld av helig ande
och brast ut och ropade högt och sade: »Välsignad vare du bland kvinnor, och välsignad din livsfrukt!
Men varför sker mig detta, att min Herres moder kommer till mig?
Se, när ljudet av din hälsning nådde mina öron, spratt barnet till av fröjd i mitt liv.
Och salig är du, som trodde att det skulle fullbordas, som blev dig sagt från Herren.»
Då sade Maria: »Min själ prisar storligen Herren,
och min ande fröjdar sig i Gud, min Frälsare.
Ty han har sett till sin tjänarinnas ringhet; och se, härefter skola alla släkten prisa mig salig.
Ty den Mäktige har gjort stora ting med mig, och heligt är hans namn.
Hans barmhärtighet varar från släkte till släkte över dem som frukta honom.
Han har utfört väldiga gärningar med sin arm, han har förskingrat dem som tänkte övermodiga tankar i sina hjärtan.
Härskare har han störtat från deras troner, och ringa män har han upphöjt;
hungriga har han mättat med sitt goda, och rika har han skickat bort med tomma händer.
Han har tagit sig an sin tjänare Israel och tänkt på att bevisa barmhärtighet
mot Abraham och mot hans säd till evig tid, efter sitt löfte till våra fäder.»
Och Maria stannade hos henne vid pass tre månader och vände därefter hem igen.
Så var nu för Elisabet tiden inne, då hon skulle föda; och hon födde en son.
Och när hennes grannar och fränder fingo höra att Herren hade bevisat henne så stor barmhärtighet, gladde de sig med henne.
Och på åttonde dagen kommo de för att omskära barnet; och de ville kalla honom Sakarias, efter hans fader.
Men hans moder tog till orda och sade: »Ingalunda; han skall heta Johannes.»
Då sade de till henne: »I din släkt finnes ju ingen som har det namnet.»
Och de frågade hans fader genom tecken vad han ville att barnet skulle heta.
Då begärde han en tavla och skrev dessa ord: »Johannes är hans namn.»
Och alla förundrade sig.
Men i detsamma öppnades hans mun, och hans tunga löstes, och han talade och lovade Gud.
Och deras grannar betogos alla av häpnad, och ryktet om allt detta gick ut över Judeens hela bergsbygd.
Och alla som hörde det lade märke därtill och sade: »Vad månde väl varda av detta barn?»
Också var ju Herrens hand med honom.
Och hans fader Sakarias blev uppfylld av helig ande och profeterade och sade:
»Lovad vare Herren, Israels Gud, som har sett till sitt folk och berett det förlossning,
och som har upprättat åt oss ett frälsningens horn i sin tjänare Davids hus,
såsom han hade lovat genom sin forntida heliga profeters mun.
Ty han ville frälsa oss från våra ovänner och ur alla våra motståndares hand,
och så göra barmhärtighet med våra fäder och tänka på sitt heliga förbund,
vad han med ed hade lovat för vår fader Abraham,
Han ville beskära oss att få tjäna honom utan fruktan, frälsta ur våra ovänners hand,
ja, att göra tjänst inför honom i helighet och rättfärdighet i alla våra dagar.
Och du, barn, skall bliva kallad den Högstes profet, ty du skall gå framför Herren och bereda vägar för honom,
till att giva hans folk kunskap om frälsning, i det att deras synder bliva dem förlåtna.
Så skall ske för vår Guds förbarmande kärleks skull, som skall låta ett ljus gå upp och skåda ned till oss från höjden,
för att 'skina över dem som sitta i mörker och dödsskugga' och så styra våra fötter in på fridens väg.»
Och barnet växte upp och blev allt starkare i anden.
Och han vistades i öknen, intill den dag då han skulle träda fram för Israel.
Och det hände sig vid den tiden att från kejsar Augustus utgick ett påbud att hela världen skulle skattskrivas.
Detta var den första skattskrivningen, och den hölls, när Kvirinius var landshövding över Syrien.
Då färdades alla var och en till sin stad, för att låta skattskriva sig.
Så gjorde ock Josef; och eftersom han var av Davids hus och släkt, for han från staden Nasaret i Galileen upp till Davids stad, som heter Betlehem, i Judeen,
för att låta skattskriva sig jämte Maria, sin trolovade, som var havande.
Medan de voro där, hände sig att tiden var inne, då hon skulle föda.
Och hon födde sin förstfödde son och lindade honom och lade honom i en krubba, ty det fanns icke rum för dem i härbärget.
I samma nejd voro då några herdar ute på marken och höllo vakt om natten över sin hjord.
Då stod en Herrens ängel framför dem, och Herrens härlighet kringstrålade dem; och de blevo mycket förskräckta.
Men ängeln sade till dem: »Varen icke förskräckta.
Se, jag bådar eder en stor glädje, som skall vederfaras allt folket.
Ty i dag har en Frälsare blivit född åt eder i Davids stad, och han är Messias, Herren.
Och detta skall för eder vara tecknet: I skolen finna ett nyfött barn, som ligger lindat i en krubba.»
I detsamma sågs där jämte ängeln en stor hop av den himmelska härskaran, och de lovade Gud och sade:
»Ära vare Gud i höjden, och frid på jorden, bland människor till vilka han har behag!»
När så änglarna hade farit ifrån herdarna upp i himmelen, sade dessa till varandra: »Låt oss nu gå till Betlehem och se det som där har skett, och som Herren har kungjort för oss.»
Och de skyndade åstad dit och funno Maria och Josef, och barnet som låg i krubban.
Och när de hade sett det, omtalade de vad som hade blivit sagt till dem om detta barn.
Och alla som hörde det förundrade sig över vad herdarna berättade för dem.
Men Maria gömde och begrundade allt detta i sitt hjärta.
Och herdarna vände tillbaka och prisade och lovade Gud för allt vad de hade fått höra och se, alldeles såsom det blivit dem sagt.
När sedan åtta dagar hade gått till ända och han skulle omskäras, gavs honom namnet Jesus, det namn som hade blivit nämnt av ängeln, förrän han blev avlad i sin moders liv.
Och när deras reningsdagar hade gått till ända, de som voro föreskrivna i Moses' lag, förde de honom upp till Jerusalem för att bära honom fram inför Herren,
enligt den föreskriften i Herrens lag, att »allt mankön som öppnar moderlivet skall räknas såsom helgat åt Herren»,
så ock för att offra »ett par duvor eller två unga turturduvor», såsom stadgat var i Herrens lag.
I Jerusalem levde då en man, vid namn Simeon, en rättfärdig och from man, som väntade på Israels tröst; och helig ande var över honom.
Och av den helige Ande hade han fått den uppenbarelsen att han icke skulle se döden, förrän han hade fått se Herrens Smorde.
Han kom nu genom Andens tillskyndelse till helgedomen.
Och när föräldrarna buro in barnet Jesus, för att så göra med honom som sed var efter lagen,
då tog också han honom i sin famn och lovade Gud och sade:
»Herre, nu låter du din tjänare fara hädan i frid, efter ditt ord,
ty mina ögon hava sett din frälsning,
vilken du har berett till att skådas av alla folk:
ett ljus som skall uppenbaras för hedningarna, och en härlighet som skall givas åt ditt folk Israel.»
Och hans fader och moder förundrade sig över det som sades om honom.
Och Simeon välsignade dem och sade till Maria, hans moder: »Se, denne är satt till fall eller upprättelse för många i Israel, och till ett tecken som skall bliva motsagt.
Ja, också genom din själ skall ett svärd gå.
Så skola många hjärtans tankar bliva uppenbara.»
Där fanns ock en profetissa, Hanna, Fanuels dotter, av Asers stam.
Hon var kommen till hög ålder; i sju år hade hon levat med sin man, från den tid då hon var jungfru,
och hon var nu änka, åttiofyra år gammal.
Och hon lämnade aldrig helgedomen, utan tjänade där Gud med fastor och böner, natt och dag.
Hon kom också i samma stund tillstädes och prisade Gud och talade om honom till alla dem som väntade på förlossning för Jerusalem.
Och när de hade fullgjort allt som var stadgat i Herrens lag, vände de tillbaka till sin stad, Nasaret i Galileen.
Men barnet växte upp och blev allt starkare och uppfylldes av vishet; och Guds nåd var över honom.
Nu plägade hans föräldrar årligen vid påskhögtiden begiva sig till Jerusalem.
När han var tolv år gammal, gingo de också dit upp, såsom sed var vid högtiden.
Men när de hade varit med om alla högtidsdagarna och vände hem igen, stannade gossen Jesus kvar i Jerusalem, utan att hans föräldrar lade märke därtill.
De menade att han var med i ressällskapet och vandrade så en dagsled och sökte efter honom bland fränder och vänner.
När de då icke funno honom, vände de tillbaka till Jerusalem och sökte efter honom.
Och efter tre dagar funno de honom i helgedomen, där han satt mitt ibland lärarna och hörde på dem och frågade dem;
och alla som hörde honom blevo uppfyllda av häpnad över hans förstånd och hans svar.
När de nu fingo se honom där, förundrade de sig högeligen; och hans moder sade till honom: »Min son, varför gjorde du oss detta?
Se, din fader och jag hava sökt efter dig med stor oro.»
Då sade han till dem: »Varför behövden I söka efter mig?
Vissten I då icke att jag bör vara där min Fader bor?»
Men de förstodo icke det som han talade till dem.
Så följde han med dem och kom ned till Nasaret; och han var dem underdånig.
Och hans moder gömde allt detta i sitt hjärta.
Och Jesus växte till i ålder och vishet och nåd inför Gud och människor.
I femtonde året av kejsar Tiberius' regering, när Pontius Pilatus var landshövding i Judeen, och Herodes var landsfurste i Galileen, och hans broder Filippus landsfurste i Itureen och Trakonitis-landet, och Lysanias landsfurste i Abilene,
på den tid då Hannas var överstepräst jämte Kaifas -- då kom Guds befallning till Johannes, Sakarias' son, i öknen;
och han gick åstad och predikade i hela trakten omkring Jordan bättringens döpelse till syndernas förlåtelse.
Så uppfylldes vad som var skrivet i profeten Esaias' utsagors bok: »Hör rösten av en som ropar i öknen: Bereden vägen för Herren, gören stigarna jämna för honom.
Alla dalar skola fyllas och alla berg och höjder sänkas; vad krokigt är skall bliva rak väg, och vad oländigt är skall bliva släta stigar;
och allt kött skall se Guds frälsning.'»
Han sade nu till folket som kom ut för att låta döpa sig av honom: »I huggormars avföda, vem har ingivit eder att söka komma undan den tillstundande vredesdomen?
Bären då ock sådan frukt som tillhör bättringen.
Och sägen icke vid eder själva: 'Vi hava ju Abraham till fader'; Ty jag säger eder att Gud av dessa stenar kan uppväcka barn åt Abraham.
Redan är också yxan satt till roten på träden; så bliver då vart träd som icke bär god frukt avhugget och kastat på elden.
Och folket frågade honom och sade: »Vad skola vi då göra?»
Han svarade och sade till dem: »Den som har två livklädnader, han dele med sig åt den som icke har någon; och en som har matförråd, han göre sammalunda.»
Så kommo ock publikaner för att låta döpa sig, och de sade till honom: »Mästare, vad skola vi göra?»
Han svarade dem: »Kräven icke ut mer än vad som är eder föreskrivet.»
Också krigsmän frågade honom och sade: »Vad skola då vi göra?
Han svarade dem: »Tilltvingen eder icke penningar av någon, genom hot eller på annat otillbörligt sätt, utan låten eder nöja med eder sold.»
Och folket gick där i förbidan, och alla undrade i sina hjärtan om Johannes icke till äventyrs vore Messias.
Men Johannes tog till orda och sade: till dem alla: »Jag döper eder med vatten, men den som kommer, som är starkare än jag, den vilkens skorem jag icke är värdig att upplösa; han skall döpa eder i helig ande och eld.
Han har sin kastskovel i handen, ty han vill noga rensa sin loge och samla in vetet i sin lada; men agnarna skall han bränna upp i en eld som icke utsläckes.»
Så förmanade han folket också i många andra stycken och förkunnade evangelium för dem.
Men när han hade förehållit Herodes, landsfursten, hans synd i fråga om hans broders hustru Herodias och förehållit honom allt det onda som han eljest hade gjort,
lade Herodes till allt annat också det att han inspärrade Johannes i fängelse.
När nu allt folket lät döpa sig och jämväl Jesus blev döpt, så skedde därvid, medan han bad, att himmelen öppnades,
och den helige Ande sänkte sig ned över honom I lekamlig skepnad såsom en duva; och från himmelen kom en röst: »Du är min älskade Son; i dig har jag funnit behag.»
Och Jesus var vid pass trettio år gammal, när han begynte sitt verk.
Och man menade att han var son av Josef, som var son av Eli,
som var son av Mattat, som var son av Levi, som var son av Melki, som var son av Jannai, som var son av Josef,
som var son av Mattatias, som var son av Amos, som var son av Naum, som var son av Esli, som var son av Naggai,
som var son av Maat, som var son av Mattatias, som var son av Semein, som var son av Josek, som var son av Joda,
som var son av Joanan, som var son av Resa, som var son av Sorobabel, som var son av Salatiel, som var son av Neri,
som var son av Melki, som var son av Addi, som var son av Kosam, som var son av Elmadam, som var son av Er,
som var son av Jesus, som var son av Elieser, som var son av Jorim, som var son av Mattat, som var son av Levi,
som var son av Simeon, som var son av Judas, som var son av Josef, som var son av Jonam, som var son av Eljakim,
som var son av Melea, som var son av Menna, som var son av Mattata, som var son av Natam, som var son av David,
som var son av Jessai, som var son av Jobed, som var son av Boos, som var son av Sala, som var son av Naasson,
som var son av Aminadab, som var son av Admin, som var son av Arni, som var son av Esrom, som var son av Fares, som var son av Judas,
som var son av Jakob, som var son av Isak, som var son av Abraham, som var son av Tara, som var son av Nakor,
som var son av Seruk, som var son av Ragau, som var son av Falek, som var son av Eber, som var son av Sala,
som var son av Kainam, som var son av Arfaksad, som var son av Sem, som var son av Noa, som var son av Lamek,
som var son av Matusala, som var son av Enok, som var son av Jaret som var son av Maleleel, som var son av Kainan,
som var son av Enos, som var son av Set, som var son av Adam, som var son av Gud.
Sedan vände Jesus tillbaka från Jordan, full av helig ande, och fördes genom Anden omkring i öknen
och frestades av djävulen under fyrtio dagar.
Och under de dagarna åt han intet; men när de hade gått till ända, blev han hungrig.
Då sade djävulen till honom: »Är du Guds Son, så bjud denna sten att bliva bröd.»
Jesus svarade honom: »Det är skrivet: 'Människan skall leva icke allenast av bröd.'»
Och djävulen förde honom upp på en höjd och visade honom i ett ögonblick alla riken i världen
och sade till honom: »Åt dig vill jag giva makten över allt detta med dess härlighet; ty åt mig har den blivit överlämnad, och åt vem jag vill kan jag giva den.
Om du alltså tillbeder inför mig, så skall den hel och hållen höra dig till.»
Jesus svarade och sade till honom: »Det är skrivet: 'Herren, din Gud, skall du tillbedja, och honom allena skall du tjäna.'»
Och han förde honom till Jerusalem och ställde honom uppe på helgedomens mur och sade till honom: »Är du Guds Son, så kasta dig ned härifrån;
det är ju skrivet: 'Han skall giva sina änglar befallning om dig, att de skola väl bevara dig';
så ock: 'De skola bära dig på händerna, så att du icke stöter din fot mot någon sten.'»
Då svarade Jesus och sade till honom: »Det är sagt: 'Du skall icke fresta Herren, din Gud.'»
När djävulen så hade slutat med alla sina frestelser, vek han ifrån honom, intill läglig tid.
Och Jesus vände i Andens kraft tillbaka till Galileen; och ryktet om honom gick ut i hela den kringliggande trakten.
Och han undervisade i deras synagogor och blev prisad av alla.
Så kom han till Nasaret, där han var uppfödd.
Och på sabbatsdagen gick han, såsom hans sed var, in i synagogan: och där stod han upp till att föreläsa.
Då räckte man åt honom profeten Esaias' bok; och när han öppnade boken, fick han se det ställe där det stod skrivet:
»Herrens Ande är över mig, ty han har smort mig.
Han har satt mig till att förkunna glädjens budskap för de fattiga, till att predika frihet för de fångna och syn för de blinda, ja, till att giva de förtryckta frihet
och till att predika ett nådens år från Herren.»
Sedan lade han ihop boken och gav den tillbaka åt tjänaren och satte sig ned.
Och alla som voro i synagogan hade sina ögon fästa på honom.
Då begynte han tala och sade till dem: »I dag är detta skriftens ord fullbordat inför edra öron.»
Och de gåvo honom alla sitt vittnesbörd och förundrade sig över de nådens ord som utgingo från hans mun, och sade: »Är då denne icke Josefs son?»
Då sade han till dem: »Helt visst skolen I nu vända mot mig det ordet: 'Läkare, bota dig själv' och säga: 'Sådana stora ting som vi hava hört vara gjorda i Kapernaum, sådana må du göra också här i din fädernestad.'»
Och han tillade: »Sannerligen säger jag eder: Ingen profet bliver i sitt fädernesland väl mottagen.
Men jag säger eder, såsom sant är: I Israel funnos många änkor på Elias' tid då himmelen var tillsluten i tre år och sex månader, och stor hungersnöd kom över hela landet --
och likväl blev Elias icke sänd till någon av dessa, utan allenast till en änka i Sarepta i Sidons land.
Och många spetälska funnos i Israel på profeten Elisas tid; och likväl blev ingen av dessa gjord ren, utan allenast Naiman från Syrien.»
När de som voro i synagogan hörde detta, uppfylldes de alla av vrede
och stodo upp och drevo honom ut ur staden och förde honom ända fram till branten av det berg som deras stad var byggd på, och ville störta honom därutför.
Men han gick sin väg mitt igenom hopen och vandrade vidare.
Och han kom ned till Kapernaum, en stad i Galileen, och undervisade folket på sabbaten.
Och de häpnade över hans undervisning, ty han talade med makt och myndighet.
Och i synagogan var en man som var besatt av en oren ond ande.
Denne ropade med hög röst:
»Bort härifrån!
Vad har du med oss att göra, Jesus från Nasaret?
Har du kommit för att förgöra oss?
Jag vet vem du är, du Guds Helige.»
Men Jesus tilltalade honom strängt och sade: »Tig och far ut ur honom.»
Då kastade den onde anden omkull mannen mitt ibland dem och for ut ur honom, utan att hava gjort honom någon skada.
Och häpnad kom över dem alla, och de talade med varandra och sade: »Vad är det med dennes ord?
Med myndighet och makt befaller han ju de orena andarna, och de fara ut.»
Och ryktet om honom spriddes åt alla håll i den kringliggande trakten.
Men han stod upp och gick ut ur synagogan och kom in i Simons hus.
Och Simons svärmoder var ansatt av en svår feber, och de bådo honom för henne.
Då trädde han fram och lutade sig över henne och näpste febern, och den lämnade henne; och strax stod hon upp och betjänade dem.
Men när solen gick ned, förde alla till honom sina sjuka, sådana som ledo av olika slags sjukdomar.
Och han lade händerna på var och en av dem och botade dem.
Onda andar blevo ock utdrivna ur många, och de ropade därvid och sade: »Du är Guds Son.»
Men han tilltalade dem strängt och tillsade dem att icke säga något, eftersom de visste att han var Messias.
Och när det åter hade blivit dag, gick han åstad bort till en öde trakt.
Men folket sökte efter honom; och när de kommo fram till honom, ville de hålla honom kvar och hindra honom att gå sin väg.
Men han sade till dem: »Också för de andra städerna måste jag förkunna evangelium om Guds rike, ty därtill har jag blivit utsänd.»
Och han predikade i synagogorna i Judeen.
Då nu en gång folket, för att höra Guds ord, trängde sig inpå honom där han stod vid Gennesarets sjö,
fick han se två båtar ligga vid sjöstranden; men de som fiskade hade gått i land och höllo på att skölja sina nät.
Då steg han i en av båtarna, den som tillhörde Simon, och bad honom lägga ut något litet från land.
Sedan satte han sig ned och undervisade folket från båten.
Och när han hade slutat att tala, sade han till Simon: »Lägg ut på djupet; och kasten där ut edra nät till fångst.»
Då svarade Simon och sade: »Mästare, vi hava arbetat hela natten och fått intet; men på ditt ord vill jag kasta ut näten.»
Och när de hade gjort så, fingo de en stor hop fiskar i sina nät; och näten gingo sönder.
Då vinkade de åt sina kamrater i den andra båten, att dessa skulle komma och hjälpa dem.
Och de kommo och fyllde upp båda båtarna, så att de begynte sjunka.
När Simon Petrus såg detta, föll han ned för Jesu knän och sade: »Gå bort ifrån mig, Herre; jag är en syndig människa.»
Ty för detta fiskafänges skull hade han och alla som voro med honom betagits av häpnad,
jämväl Jakob och Johannes, Sebedeus' söner, som deltogo med Simon i fisket.
Men Jesus sade till Simon: »Frukta icke; härefter skall du fånga människor.»
Och de förde båtarna i land och lämnade alltsammans och följde honom.
Och medan han var i en av städerna, hände sig, att där kom en man som var full av spetälska.
När denne fick se Jesus, föll han ned på sitt ansikte och bad honom och sade: »Herre, vill du, så kan du göra mig ren.»
Då räckte han ut handen och rörde vid honom och sade: »Jag vill; bliv ren.»
Och strax vek spetälskan ifrån honom.
Och han förbjöd honom att omtala detta för någon, men tillade: »Gå åstad och visa dig för prästen och frambär för din rening ett offer, såsom Moses har påbjudit, till ett vittnesbörd för dem.»
Men ryktet om honom spridde sig dess mer; och mycket folk samlade sig för att höra honom och för att bliva botade från sina sjukdomar.
Men han drog sig undan till öde trakter och bad.
Nu hände sig en dag, då han undervisade folket, att där sutto några fariséer och laglärare -- sådana hade nämligen kommit dit från alla byar i Galileen och Judeen och från Jerusalem -- och Herrens kraft verkade, så att sjuka blevo botade av honom.
Då kommo några män dit med en lam man, som de buro på en säng; och de försökte komma in med honom för att lägga honom ned framför Jesus.
Men då de för folkets skull icke kunde finna något annat sätt att komma in med honom stego de upp på taket och släppte honom tillika med sängen ned genom tegelbeläggningen, mitt ibland dem, framför Jesus.
När han såg deras tro, sade han: »Min vän, dina synder äro dig förlåtna.»
Då begynte de skriftlärde och fariséerna tänka så: »Vad är denne för en, som talar så hädiska ord?
Vem kan förlåta synder utom Gud allena?»
Men Jesus förnam deras tankar och svarade och sade till dem: »Vad är det I tänken i edra hjärtan?
Vilket är lättare att säga: 'Dina synder äro dig förlåtna' eller att säga: 'Stå upp och gå'?
Men för att I skolen veta, att Människosonen har makt här på jorden att förlåta synder, så säger jag dig» (och härmed vände han sig till den lame): »Stå upp, tag din säng och gå hem.»
Då stod han strax upp i deras åsyn och tog sängen, som han hade legat på, och gick hem, prisande Gud.
Och de grepos alla av bestörtning och prisade Gud; och de sade, fulla av häpnad: »Vi hava i dag sett förunderliga ting.»
Sedan begav han sig därifrån.
Och han fick se en publikan, vid namn Levi, sitta vid tullhuset.
Och han sade till denne: »Följ mig.»
Då lämnade han allt och stod upp och följde honom.
Och Levi gjorde i sitt hus ett stort gästabud för honom; och en stor hop publikaner och andra voro bordsgäster där jämte dem.
Men fariséerna -- särskilt de skriftlärde bland dem -- knorrade mot hans lärjungar och sade: »Huru kunnen I äta och dricka med publikaner och syndare?»
Då svarade Jesus och sade till dem: »De är icke de friska som behöva läkare, utan de sjuka.
Jag har icke kommit för att kalla rättfärdiga, utan syndare, till bättring.
Och de sade till honom: »Johannes' lärjungar fasta ofta och hålla böner, sammalunda ock fariséernas; men dina lärjungar äta och dricka.»
Jesus svarade dem: »Icke kunnen I väl ålägga bröllopsgästerna att fasta, medan brudgummen ännu är hos dem?
Men en annan tid skall komma, och då, när brudgummen tages ifrån dem, då, på den tiden, skola de fasta.» --
Han framställde ock för dem denna liknelse: »Ingen river av en lapp från en ny mantel och sätter den på en gammal mantel; om någon så gjorde, skulle han icke allenast riva sönder den nya manteln, utan därtill komme, att lappen från den nya manteln icke skulle passa den gamla.
Ej heller slår någon nytt vin i gamla skinnläglar; om någon så gjorde, skulle det nya vinet spränga sönder läglarna, och vinet skulle spillas ut, jämte det att läglarna fördärvades.
Nej, nytt vin bör man slå i nya läglar. --
Och ingen som har druckit gammalt vin vill sedan gärna hava nytt; ty han tycker, att det gamla är bättre.»
Och det hände sig på en sabbat att han tog vägen genom ett sädesfält; och hans lärjungar ryckte av axen och gnuggade sönder dem med händerna och åto.
Då sade några av fariséerna; »Huru kunnen I göra vad som icke är lovligt att göra på sabbaten?
Jesus svarade och sade till dem: »Haven I icke läst om det som David gjorde, när han själv och de som följde honom blevo hungriga:
huru han då gick in i Guds hus och tog skådebröden och åt, och jämväl gav åt dem som följde honom, fastän det ju icke är lovligt för andra än allenast för prästerna att äta sådant bröd?»
Därefter sade han till dem: »Människosonen är herre över sabbaten.»
På en annan sabbat hände sig att han gick in i synagogan och undervisade.
Där var då en man vilkens högra hand var förvissnad.
Och de skriftlärde och fariséerna vaktade på honom, för att se om han botade någon på sabbaten; de ville nämligen finna något att anklaga honom för.
Men han förstod deras tankar och sade till mannen som hade den förvissnade handen: »Stå upp, och träd fram.»
Då stod han upp och trädde fram.
Sedan sade Jesus till dem: »Jag vill göra eder en fråga.
Vilketdera är lovligt på sabbaten: att göra vad gott är, eller att göra vad ont är, att rädda någons liv, eller att förgöra det?»
Och han såg sig omkring på dem alla och sade till mannen: »Räck ut din hand.»
Och han gjorde så; och hans hand blev frisk igen.
Men de blevo såsom ursinniga och talade med varandra om vad de skulle kunna företaga sig mot Jesus.
Så hände sig på den tiden att han gick åstad upp på berget för att bedja; och han blev kvar där över natten i bön till Gud.
Men när det blev dag, kallade han till sig sina lärjungar och utvalde bland dem tolv, som han ock benämnde apostlar:
Simon, vilken han ock gav namnet Petrus, och Andreas, hans broder; vidare Jakob och Johannes och Filippus och Bartolomeus
och Matteus och Tomas och Jakob, Alfeus' son, och Simon, som kallades ivraren;
vidare Judas, Jakobs son, och Judas Iskariot, den som blev en förrädare.
Dessa tog han nu med sig och steg åter ned och stannade på en jämn plats; och en stor skara av hans lärjungar var där församlad, så ock en stor hop folk ifrån hela Judeen och Jerusalem, och från kuststräckan vid Tyrus och Sidon.
Dessa hade kommit för att höra honom och för att bliva botade från sina sjukdomar.
Och jämväl de som voro kvalda av orena andar blevo botade.
Och allt folket sökte att få röra vid honom, ty kraft gick ut ifrån honom och botade alla.
Och han lyfte upp sina ögon och säg på sina lärjungar och sade: »Saliga ären I, som ären fattiga, ty eder hör Guds rike till.
Saliga ären I, som nu hungren, ty I skolen bliva mättade.
Saliga ären I, som nu gråten, ty I skolen le.
Saliga ären I, när människorna för Människosonens skull hata eder och förskjuta och smäda eder och kasta bort edert namn såsom något ont.
Glädjens på den dagen, ja, springen upp av fröjd, ty se, eder lön är stor i himmelen.
På samma satt gjorde ju deras fäder med profeterna.
Men ve eder, I som ären rika, ty I haven fått ut eder hugnad!
Ve eder, som nu ären mätta, ty I skolen hungra!
Ve eder, som nu len, ty I skolen sörja och gråta!
Ve eder, när alla människor tala väl om eder!
På samma sätt gjorde ju deras fader i fråga om de falska profeterna.
Men till eder, som hören mig, säger jag: Älsken edra ovänner, gören gott mot dem som hata eder,
välsignen dem som förbanna eder, bedjen för dem som förorätta eder.
Om någon slår dig på den ena kinden, så håll ock fram den andra åt honom; och om någon tager manteln ifrån dig, så förvägra honom icke heller livklädnaden.
Giv åt var och en som beder dig; och om någon tager ifrån dig vad som är ditt, så kräv det icke igen.
Såsom I viljen att människorna skola göra mot eder, så skolen I ock göra mot dem.
Om I älsken dem som älska eder, vad tack kunnen I få därför?
Också syndare älska ju dem av vilka de bliva älskade.
Och om I gören gott mot dem som göra eder gott, vad tack kunnen I få därför?
Också syndare göra ju detsamma.
Och om I lånen åt dem av vilka I kunnen hoppas att själva få något, vad tack kunnen I få därför?
Också syndare låna ju åt syndare för att få lika igen.
Nej, älsken edra ovänner, och gören gott och given lån utan att hoppas på någon gengäld.
Då skall eder lön bliva stor, och då skolen I vara den Högstes barn; ty han är mild mot de otacksamma och onda.
Varen barmhärtiga, såsom eder Fader är barmhärtig.
Dömen icke, så skolen I icke bliva dömda; fördömen icke, så skolen I icke bliva fördömda.
Förlåten, och eder skall bliva förlåtet.
Given, och eder skall bliva givet.
Ett gott mått, väl packat, skakat och överflödande, skall man giva eder i skötet; ty med det mått som I mäten med skall ock mätas åt eder igen.»
Han framställde ock för dem denna liknelse: »Kan väl en blind leda en blind?
Falla de icke då båda i gropen?
Lärjungen är icke förmer än sin mästare; när någon bliver fullärd, så bliver han allenast sin mästare lik.
Huru kommer det till, att du ser grandet i din broders öga, men icke bliver varse bjälken i ditt eget öga?
Huru kan du säga till din broder: 'Broder, låt mig taga ut grandet i ditt öga', du som icke ser bjälken i ditt eget öga?
Du skrymtare, tag först ut bjälken ur ditt eget öga; därefter må du se till, att du kan tala ut grandet i din broders öga.
Ty intet gott träd finnes, som bär dålig frukt, och lika litet finnes något dåligt träd som bär god frukt;
vart och ett träd kännes ju igen på sin frukt.
Icke hämtar man väl fikon ifrån törnen, ej heller skördar man vindruvor av törnbuskar.
En god människa bär ur sitt hjärtas goda förråd fram vad gott är, och en ond människa bär ur sitt onda förråd fram vad ont är; ty vad hennes hjärta är fullt av, det talar hennes mun. --
Men varför ropen I till mig: 'Herre, Herre', och gören dock icke vad jag säger?
Var och en som kommer till mig och hör mina ord och gör efter dem, vem han är lik, det skall jag visa eder.
Han är lik en man som ville bygga ett hus och som då grävde djupt och lade dess grund på hälleberget.
När sedan översvämning kom, störtade sig vattenströmmen mot det huset, men den förmådde dock icke skaka det, eftersom det var så byggt.
Men den som hör och icke gör, han är lik en man som byggde ett hus på blotta jorden, utan att lägga någon grund.
Och vattenströmmen störtade sig emot det, och strax föll det samman, och det husets fall blev stort.»
När han nu hade talat allt detta till slut inför folket, gick han in i Kapernaum.
Men där var en hövitsman som hade en tjänare, vilken låg sjuk och var nära döden; och denne var högt skattad av honom.
Då han nu fick höra om Jesus, sände han till honom några av judarnas äldste och bad honom komma och bota hans tjänare.
När dessa kommo till Jesus, bådo de honom enträget och sade: »Han är värd att du gör honom detta,
ty han har vårt folk kärt, och det är han som har byggt synagogan åt oss.»
Då gick Jesus med dem.
Men när han icke var långt ifrån hövitsmannens hus, sände denne några av sina vänner och lät säga till honom: »Herre, gör dig icke omak; ty jag är icke värdig att du går in under mitt tak.
Därför har jag ej heller aktat mig själv värdig att komma till dig Men säg ett ord, så bliver min tjänare frisk.
Jag är ju själv en man som står under andras befäl; jag har ock krigsmän under mig, och om jag säger till en av dem: 'Gå', så går han, eller till en annan: 'Kom', så kommer han, och om jag säger till min tjänare: 'Gör det', då gör han så.»
När Jesus hörde detta, förundrade han sig över honom och vände sig om och sade till folket som följde honom: »Jag säger eder: Icke ens i Israel har jag funnit så stor tro.»
Och de som hade blivit utsända gingo hem igen och funno tjänaren vara frisk.
Därefter begav han sig till en stad som hette Nain; och med honom gingo hans lärjungar och mycket folk.
Och se, då han kom nära stadsporten, bars där ut en död, och han var sin moders ende son, och hon var änka; och en ganska stor hop folk ifrån staden gick med henne.
När Herren fick se henne, ömkade han sig över henne och sade till henne: »Gråt icke.»
Och han gick fram och rörde vid båren, och de som buro stannade.
Och han sade: »Unge man, jag säger dig: Stå upp.»
Då satte sig den döde upp och begynte tala.
Och han gav honom åt hans moder.
Och alla betogos av häpnad och prisade Gud och sade: Den stor profet har uppstått ibland oss» och: »Gud har sett till sitt folk.»
Och detta tal om honom gick ut i hela Judeen och i hela landet däromkring.
Och allt detta fick Johannes höra berättas av sina lärjungar.
Då kallade Johannes till sig två av sina lärjungar och sände dem till Herren med denna fråga: »Är du den som skulle komma, eller skola vi förbida någon annan?»
När mannen kommo fram till honom, sade de: »Johannes döparen har sänt oss till dig och låter fråga: 'Är du den som skulle komma, eller skola vi förbida någon annan?'»
Just då höll Jesus på med att bota många som ledo av sjukdomar och plågor, eller som voro besatta av onda andar, och åt många blinda gav han deras syn.
Och han svarade och sade till männen: »Gån tillbaka och omtalen för Johannes vad I haven sett och hört: blinda få sin syn, halta gå, spetälska bliva rena, döva höra, döda uppstå, 'för fattiga förkunnas glädjens budskap'.
Och salig är den för vilken jag icke bliver en stötesten.»
När sedan Johannes' sändebud hade gått sin väg, begynte han tala till folket om Johannes: »Varför var det I gingen ut i öknen?
Var det för att se ett rör som drives hit och dit av vinden?
Eller varför gingen I ut?
Var det för att se en människa klädd i fina kläder?
De som bära präktiga kläder och leva i kräslighet, dem finnen I ju i konungapalatsen.
Varför gingen I då ut?
Var det för att se en profet?
Ja, jag säger eder: Ännu mer än en profet är han.
Han är den om vilken det är skrivet: 'Se, jag sänder ut min ängel framför dig, och han skall bereda vägen för dig.'
Jag säger eder: Bland dem som äro födda av kvinnor har ingen varit större än Johannes; men den som är minst i Guds rike är likväl större än han.
Så gav ock allt folket som hörde honom Gud rätt, jämväl publikanerna, och läto döpa sig med Johannes' dop.
Men fariséerna och de lagkloke föraktade Guds rådslut i fråga om dem själva och läto icke döpa sig av honom.
Vad skall jag då likna detta släktes människor vid?
Ja, vad äro de lika?
De äro lika barn som sitta på torget och ropa till varandra och säga: 'Vi hava spelat för eder, och I haven icke dansat; vi hava sjungit sorgesång, och I haven icke gråtit.'
Ty Johannes döparen har kommit, och han äter icke bröd och dricker ej heller vin, och så sägen I: 'Han är besatt av en ond ande.'
Människosonen har kommit, och han både äter och dricker, och nu sägen I: 'Se, vilken frossare och vindrinkare han är, en publikaners och syndares vän!'
Men Visheten har fått rätt av alla sina barn.»
Och en farisé inbjöd honom till en måltid hos sig; och han gick in i fariséens hus och lade sig till bords.
Nu fanns där i staden en synderska; och när denna fick veta att han låg till bords i fariséens hus, gick hon dit med en alabasterflaska med smörjelse
och stannade bakom honom vid hans fötter, gråtande, och begynte väta hans fötter med sina tårar och torkade dem med sitt huvudhår och kysste ivrigt hans fötter och smorde dem med smörjelsen.
Men när fariséen som hade inbjudit honom såg detta, sade han vid sig själv: »Vore denne en profet, så skulle han känna till, vilken och hurudan denna kvinna är, som rör vid honom; han skulle då veta att hon är en synderska.»
Då tog Jesus till orda och sade till honom: »Simon, jag har något att säga dig.»
Han svarade: »Mästare, säg det.
»En man som lånade ut penningar hade två gäldenärer.
Den ene var skyldig honom fem hundra silverpenningar, den andre femtio.
Men då de icke kunde betala, efterskänkte han skulden för dem båda.
Vilken av dem kommer nu att älska honom mest?»
Simon svarade och sade: »Jag menar den åt vilken han efterskänkte mest.»
Då sade han till honom: »Rätt dömde du»
Och så vände han sig åt kvinnan och sade till Simon: »Ser du denna kvinna?
När jag kom in i ditt hus, gav du mig intet vatten till mina fötter, men hon har vätt mina fötter med sina tårar och torkat dem med sitt hår.
Du gav mig ingen hälsningskyss, men ända ifrån den stund då jag kom hitin, har hon icke upphört att ivrigt kyssa mina fötter.
Du smorde icke mitt huvud med olja, men hon har smort mina fötter med smörjelse.
Fördenskull säger jag dig: Hennes många synder äro henne förlåtna; hon har ju ock visat mycken kärlek.
Men den som får litet förlåtet, han älskar ock litet.»
Sedan sade han till henne: »Dina synder äro dig förlåtna.»
Då begynte de som voro bordsgäster jämte honom att säga vid sig själva: »Vem är denne, som till och med förlåter synder?»
Men han sade till kvinnan: »Din tro har frälst dig.
Gå i frid.»
Därefter vandrade han igenom landet, från stad till stad och från by till by, och predikade och förkunnade evangelium om Guds rike.
Och med honom följde de tolv,
så ock några kvinnor som hade blivit befriade från onda andar och botade från sjukdomar: Maria, som kallades Magdalena, ur vilken sju onda andar hade blivit utdrivna,
och Johanna, hustru till Herodes' fogde Kusas, och Susanna och många andra som tjänade dem med sina ägodelar.
Då nu mycket folk kom tillhopa, i det att inbyggarna i de särskilda städerna begåvo sig ut till honom, sade han i en liknelse:
»En såningsman gick ut för att så sin säd.
Och när han sådde, föll somt vid vägen och blev nedtrampat, och himmelens fåglar åto upp det.
Och somt föll på stengrund, och när det hade vuxit upp, torkade det bort, eftersom det icke där hade någon fuktighet.
Och somt föll bland törnen, och törnena växte upp tillsammans därmed och förkvävde det.
Men somt föll i god jord, och när det hade vuxit upp, bar det hundrafaldig frukt.»
Sedan han hade talat detta, sade han med hög röst: »Den som har öron till att höra, han höre.»
Då frågade hans lärjungar honom vad denna liknelse betydde.
Han sade: »Eder är givet att lära känna Guds rikes hemligheter, men åt de andra meddelas de i liknelser, för att de med seende ögon intet skola se och med hörande öron intet förstå'.
Så är nu detta liknelsens mening: Säden är Guds ord.
Och att den såddes vid vägen, det är sagt om dem som hava hört ordet, men sedan kommer djävulen och tager bort det ur deras hjärtan, för att de icke skola komma till tro och bliva frälsta.
Och att den såddes på stengrunden det är sagt om dem, som när de få höra ordet, taga emot det med glädje, men icke hava någon rot; de tro allenast till en tid, och i frestelsens stund avfalla de.
Och att den föll bland törnena, det är sagt om dem, som när de hava hört ordet, gå bort och låta sig förkvävas av rikedomens omsorger och njutandet av livets goda och så icke föra något fram till mognad.
Men att den föll i den goda jorden, det är sagt om dem, som när de hava hört ordet, behålla det i rättsinniga och goda hjärtan och bära frukt i ståndaktighet.
Ingen tänder ett ljus och gömmer det sedan under ett kärl eller sätter det under en bänk, utan man sätter det på en ljusstake, för att de som komma in skola se skenet.
Ty intet är fördolt, som icke skall bliva uppenbart, ej heller är något undangömt, som icke skall bliva känt och komma i dagen.
Akten fördenskull på huru I hören.
Ty den som har, åt honom skall varda givet; men den som icke har, från honom skall tagas också det han menar sig hava.»
Och hans moder och hans bröder kommo och sökte honom, men för folkets skull kunde de icke komma in till honom.
Då sade man till honom: »Din moder och dina broder stå härutanför och vilja träffa dig.»
Men han svarade och sade till dem: »Min moder och mina bröder äro dessa, som höra Guds ord och göra det.»
En dag steg han med sina lärjungar i en båt och sade till dem: »Låt oss fara över sjön till andra sidan.»
Och de lade ut.
Och medan de seglade fram, somnade han.
Men en stormvind for ned över sjön, och deras båt begynte fyllas med vatten, så att de voro i fara.
Då gingo de fram och väckte upp honom och sade: »Mästare, Mästare, vi förgås.»
När han så hade vaknat, näpste han vinden och vattnets vågor, och de stillades, och det blev lugnt.
Därefter sade han till dem: »Var är eder tro?»
Men de hade blivit häpna och förundrade sig och sade till varandra: »Vem är då denne?
Han befaller ju både vindarna och vattnet, och de lyda honom.»
Så foro de över till gerasenernas land, som ligger mitt emot Galileen.
Och när han hade stigit i land, kom en man från staden emot honom, en som var besatt av onda andar, och som under ganska lång tid icke hade haft kläder på sig och icke bodde i hus, utan bland gravarna.
Då nu denne fick se Jesus, skriade han och föll ned för honom och sade med hög röst: »Vad har du med mig att göra, Jesus, du Guds, den Högstes, son?
Jag beder dig, plåga mig icke.»
Jesus skulle nämligen just bjuda den orene anden att fara ut ur mannen.
Ty i lång tid hade han farit svårt fram med mannen; och väl hade denne varit fängslad med kedjor och fotbojor och hållits i förvar, men han hade slitit sönder bojorna och hade av den onde anden blivit driven ut i öknarna.
Jesus frågade honom: »Vad är ditt namn?»
Han svarade: »Legion.»
Ty det var många onda andar som hade farit in i honom.
Och dessa bådo Jesus att han icke skulle befalla dem att fara ned i avgrunden.
Nu gick där en ganska stor svinhjord i bet på berget.
Och de bådo honom att han ville tillstädja dem att fara in i svinen.
Och han tillstadde dem det.
Då gåvo sig de onda andarna åstad ut ur mannen och foro in i svinen.
Och hjorden störtade sig utför branten ned i sjön och drunknade.
Men när herdarna sågo vad som hade skett, flydde de och berättade härom i staden och på landsbygden.
Och folket gick ut för att se vad som hade skett.
När de då kommo till Jesus, funno de mannen, ur vilken de onda andarna hade blivit utdrivna, sitta invid Jesu fötter, klädd och vid sina sinnen; och de betogos av häpnad.
Och de som hade sett händelsen omtalade för dem huru den besatte hade blivit botad.
Allt folket ifrån den kringliggande trakten av gerasenernas land bad då Jesus att han skulle gå bort ifrån dem, ty de voro gripna av stor förskräckelse.
Så steg han då i en båt för att vända tillbaka.
Och mannen, ur vilken de onda andarna hade blivit utdrivna, bad honom att få följa honom.
Men Jesus tillsade honom att gå, med de orden:
»Vänd tillbaka hem, och förtälj huru stora ting Gud har gjort med dig.»
Då gick han bort och förkunnade i hela staden huru stora ting Jesus hade gjort med honom.
När Jesus kom tillbaka, mottogs han av folket; ty alla väntade de på honom.
Då kom där en man, vid namn Jairus, som var föreståndare för synagogan.
Denne föll ned för Jesu fötter och bad honom att han skulle komma till hans hus;
ty han hade ett enda barn, en dotter, vid pass tolv år gammal, som låg för döden.
Men under det att han var på väg dit, trängde folket hårt på honom.
Nu var där en kvinna som hade haft blodgång i tolv år och icke hade kunnat botas av någon.
Hon närmade sig honom bakifrån och rörde vid hörntofsen på hans mantel, och strax stannade hennes blodgång
Men Jesus frågade: »Vem var det som rörde vid mig?»
Då alla nekade till att hava gjort det, sade Petrus: »Mästare, hela folkhopen trycker och tränger dig ju.»
Men Jesus sade: »Det var någon som rörde vid mig; ty jag kände att kraft gick ut ifrån mig.»
Då nu kvinnan såg att hon icke hade blivit obemärkt, kom hon fram bävande och föll ned för honom och omtalade inför allt folket varför hon hade rört vid honom, och huru hon strax hade blivit frisk.
Då sade han till henne: »Min dotter, din tro har hjälpt dig.
Gå i frid.»
Medan han ännu talade, kom någon från synagogföreståndarens hus och sade: »Din dotter är död; du må icke vidare göra mästaren omak.»
Men när Jesus hörde detta, sade han till honom: »Frukta icke; tro allenast, så får hon liv igen.»
Och när han hade kommit fram till hans hus, tillstadde han ingen att gå med ditin, utom Petrus och Johannes och Jakob och därtill flickans fader och moder.
Och alla gräto och jämrade sig över henne.
Men han sade: »Gråten icke; hon är icke död, hon sover.»
Då hånlogo de åt honom, ty de visste ju att hon var död.
Men han tog henne vid handen och sade med hög röst: »Flicka, stå upp.»
Då kom hennes ande igen, och hon stod strax upp.
Och han tillsade att man skulle giva henne något att äta.
Och hennes föräldrar blevo uppfyllda av häpnad; men han förbjöd dem att för någon omtala vad som hade skett.
Och han kallade tillhopa de tolv och gav dem makt och myndighet över alla onda andar, så ock makt att bota sjukdomar.
Och han sände ut dem till att predika Guds rike och till att bota sjuka.
Och han sade till dem: »Tagen intet med eder på vägen, varken stav eller ränsel eller bröd eller penningar, och haven icke heller dubbla livklädnader.
Och när I haven kommit in något hus, så stannen där, till dess I lämnen den orten.
Och om man någonstädes icke tager emot eder, så gån bort ifrån den staden, och skudden stoftet av edra fötter, till ett vittnesbörd mot dem.»
Och de gingo ut och vandrade igenom landet, från by till by, och förkunnade evangelium och botade sjuka allestädes.
Men när Herodes, landsfursten, fick höra om allt detta som skedde visste han icke vad han skulle tro.
Ty somliga sade: »Det är Johannes, som har uppstått från de döda.»
Men andra sade: »Det är Elias, som har visat sig.»
Andra åter sade: »Det är någon av de gamla profeterna, som har uppstått.»
Men Herodes själv sade: »Johannes har jag låtit halshugga.
Vem är då denne, som jag hör sådant om?»
Och han sökte efter tillfälle att få se honom.
Och apostlarna kommo tillbaka och förtäljde för Jesus huru stora ting de hade gjort.
De tog han dem med sig och drog sig undan till en stad som hette Betsaida, där de kunde vara allena.
Men när folket fick veta detta, gingo de efter honom.
Och han lät dem komma till sig och talade till dem om Guds rike; och dem som behövde botas gjorde han friska.
Men dagen begynte nalkas sitt slut.
Då trädde de tolv fram och sade till honom: »Låt folket skiljas åt, så att de kunna gå bort i byarna och gårdarna häromkring och skaffa sig härbärge och få mat; vi äro ju här i en öde trakt.»
Men han sade till dem: »Given I dem att äta.»
De svarade: »Vi hava icke mer än fem bröd och två fiskar, såframt vi icke skola gå bort och köpa mat åt allt detta folk.»
Där voro nämligen vid pass fem tusen män.
Då sade han till sina lärjungar: »Låten dem lägga sig ned i matlag, femtio eller så omkring i vart.»
Och de gjorde så och läto dem alla lägga sig ned.
Därefter tog han de fem bröden och de två fiskarna och säg upp till himmelen och välsignade dem.
Och han bröt bröden och gav åt lärjungarna, för att de skulle lägga fram åt folket.
Och de åto alla och blevo mätta. sedan samlade man upp de stycken som hade blivit över efter dem, tolv korgar.
När han en gång hade dragit sig undan och var stadd i byn, voro hans lärjungar hos honom.
Och han frågade dem och sade: »Vem säger folket mig vara?»
De svarade och sade: »Johannes döparen; dock säga andra Elias; andra åter säga: 'Det är någon av de gamla profeterna, som har uppstått.'»
Då frågade han dem: »Vem sägen då I mig vara?»
Petrus svarade och sade: »Guds Smorde.»
Då förbjöd han dem strängeligen att säga detta till någon.
Och han sade: »Människosonen måste lida mycket, och han skall bliva förkastad av de äldste och översteprästerna och de skriftlärda och skall bliva dödad, men på tredje dagen skall han uppstå igen.»
Och han sade till alla: »Om någon vill efterfölja mig, så försake han sig själv och tage sitt kors på sig var dag; så följe han mig.
Ty den som vill bevara sitt liv han skall mista det; men den som mister sitt liv, för min skull, han skall bevara det.
Och vad hjälper det en människa om hon vinner hela världen, men mister sig själv eller själv går förlorad?
Den som blyges för mig och för mina ord, för honom skall Människosonen blygas, när han kom mer i sin och min Faders och de heliga änglarnas härlighet.
Men sannerligen säger jag eder: Bland dem som här stå finnas några som icke skola smaka döden, förrän de få se Guds rike.»
Vid pass åtta dagar efter det att han hade talat detta tog han Petrus och Johannes och Jakob med sig och gick upp på berget för att bedja.
Och under det att han bad, blev hans ansikte förvandlat, och hans kläder blevo skinande vita.
Och de, två män stodo där och samtalade med honom, och dessa voro Moses och Elias.
De visade sig i härlighet och talade om hans bortgång, vilken han skulle fullborda i Jerusalem.
Men Petrus och de som voro med honom voro förtyngda av sömn; då de sedan vaknade, sågo de hans härlighet och de båda männen, som stodo hos honom.
När så dessa skulle skiljas ifrån honom, sade Petrus till Jesus: »Mästare, har är oss gott att vara; låt oss göra tre hyddor, en åt dig och en åt Moses och en åt Elias.»
Han visste nämligen icke vad han sade.
Medan han så talade, kom en sky och överskyggde dem; och de blevo förskräckta, när de trädde in i skyn.
Och ur skyn kom en röst som sade: »Denne är min Son, den utvalde; hören honom.»
Och i detsamma som rösten kom, funno de Jesus vara där allena. -- Och de förtego detta och omtalade icke för någon på den tiden något av vad de hade sett.
När de dagen därefter gingo ned från berget, hände sig att mycket folk kom honom till mötes.
Då ropade en man ur folkhopen och sade: »Mästare, jag beder dig, se till min son, ty han är mitt enda barn.
Det är så, att en ande plägar gripa fatt i honom, och strax skriar han då, och anden sliter och rycker honom, och fradgan står honom om munnen.
Och det är med knapp nöd han släpper honom, sedan han har sönderbråkat honom.
Nu bad jag dina lärjungar att de skulle driva ut honom, men de kunde det icke.»
Då svarade Jesus och sade: »O du otrogna och vrånga släkte, huru länge måste jag vara hos eder och härda ut med eder?
För hit din son.»
Men ännu medan denne var på väg fram, kastade den onde anden omkull honom och slet och ryckte honom.
Då tilltalade Jesus den orene anden strängt och gjorde gossen frisk och gav honom tillbaka åt hans fader.
Och alla häpnade över Guds stora makt.
Då nu alla förundrade sig över alla de gärningar som han gjorde, sade han till sina lärjungar:
»Tagen emot dessa ord med öppna öron: Människosonen skall bliva överlämnad i människors händer.
Men de förstodo icke detta som han sade, och det var förborgat för dem, så att de icke kunde fatta det; dock fruktade de att fråga honom om det som han hade sagt.
Och bland dem uppstod tanken på vilken av dem som vore störst.
Men Jesus förstod deras hjärtans tankar och tog ett barn och ställde det bredvid sig
och sade till dem: »Den som tager emot detta barn i mitt namn, han tager emot mig, och den som tager emot mig, han tager emot honom som har sänt mig.
Ty den som är minst bland eder alla, han är störst.
Och Johannes tog till orda och sade: »Mästare, sågo huru en man drev ut onda andar genom ditt namn; och du ville hindra honom, eftersom han icke följde med oss.»
Men Jesus sade till honom: »Hindren honom icke; ty den som icke är emot eder, han är för eder.»
Då nu tiden var inne att han skulle bliva upptagen, beslöt han att ställa sin färd till Jerusalem.
Och han sände budbärare framför sig; och de gingo åstad och kommo in i en samaritisk by för att reda till åt honom.
Men folket där tog icke emot honom, eftersom han var stadd på färd till Jerusalem.
När de båda lärjungarna Jakob i och Johannes förnummo detta, sade de: »Herre, vill du att vi skola bedja att eld kommer ned från himmelen och förtär dem?»
Då vände han sig om och tillrättavisade dem.
Och de gingo till en annan by.
Medan de nu färdades fram på vägen, sade någon till honom: »Jag vill följa dig, varthelst du går.
Då svarade Jesus honom: »Rävarna hava kulor, och himmelens fåglar hava nästen; men Människosonen har ingen plats där han kan vila sitt huvud.»
Och till en annan sade han: »Föl; mig.»
Men denne svarade: »Tillstäd mig att först gå bort och begrava min fader.»
Då sade han till honom: »Låt de döda begrava sina döda; men gå du åstad och förkunna Guds rike.»
Åter en annan sade: »Jag vill följa dig, Herre, men tillstäd mig att först taga avsked av dem som höra till mitt hus.»
Då svarade Jesus honom: »Ingen som ser sig tillbaka, sedan han har satt sin hand till plogen, är skickad för Guds rike.»
Därefter utsåg Herren sjuttiotvå andra och sände ut dem framför sig, två och två, till var stad och ort dit han själv tänkte komma
»Skörden är mycken, men arbetarna äro få.
Bedjen fördenskull skördens Herre att han sänder ut arbetare till sin skörd.
Gån åstad.
Se, jag sänder eder såsom lamm mitt in ibland ulvar.
Bären ingen penningpung, ingen ränsel, inga skor, och hälsen icke på någon under vägen.
Men när I kommen in i något hus, så sägen först: 'Frid vare över detta hus.'
Om då någon finnes därinne, som är frid värd, så skall den frid I tillönsken vila över honom; varom icke, så skall den vända tillbaka över eder själva.
Och stannen kvar i det huset, och äten och dricken vad de hava att giva, ty arbetaren är värd sin lön.
Gån icke ur hus i hus.
Och när I kommen in i någon stad där man tager emot eder, så äten vad som sättes fram åt eder,
och boten de sjuka som finnas där, och sägen till dem: 'Guds rike är eder nära.'
Men när I kommen in i någon stad där man icke tager emot eder, så gån ut på dess gator och sägen:
'Till och med det stoft som låder vid våra fötter ifrån eder stad skaka vi av oss åt eder.
Men det mån I veta, att Guds rike är nära.'
Jag säger eder att det för Sodom skall på 'den dagen' bliva drägligare än för den staden.
Ve dig, Korasin!
Ve dig, Betsaida!
Ty om de kraftgärningar som äro gjorda i eder hade blivit gjorda i Tyrus och Sidon, så skulle de för länge sedan hava suttit i säck och aska och gjort bättring.
Men också skall det vid domen bliva drägligare för Tyrus och Sidon än för eder.
Och du.
Kapernaum, skall väl du bliva upphöjt till himmelen?
Nej, ned till dödsriket måste du fara. --
Den som hör eder, han hör mig, och den som förkastar eder, han förkastar mig; men den som förkastar mig, han förkastar honom som har sänt mig.»
Och de sjuttiotvå kommo tillbaka, uppfyllda av glädje, och sade: »Herre, också de onda andarna äro oss underdåniga genom ditt namn.»
Då sade han till dem: »Jag såg Satan falla ned från himmelen såsom en ljungeld.
Se, jag har givit eder makt att trampa på ormar och skorpioner och att förtrampa all ovännens härsmakt, och han skall icke kunna göra eder någon skada.
Dock, glädjens icke över att änglarna äro eder underdåniga, utan glädjens över att edra namn äro skrivna i himmelen.»
I samma stund uppfylldes han av fröjd genom den helige Ande och sade: »Jag prisar dig, Fader, du himmelens och jordens Herre, för att du väl har dolt detta för de visa och kloka, men uppenbarat det för de enfaldiga.
Ja, Fader; så har ju varit ditt behag.
Allt har av min Fader blivit för trott åt mig.
Och ingen känner vem Sonen är utom Fadern, ej heller vem Fadern är, utom Sonen och den för vilken Sonen vill göra honom känd.»
Sedan vände han sig till lärjungarna, när han var allena med dem och sade: »Saliga äro de ögon som se det I sen.
Ty jag säger eder: Många profeter och konungar ville se det som I sen men fingo dock icke se det, och höra det som I hören, men fingo dock icke höra det.»
Men en lagklok stod upp och ville snärja honom och sade: »Mästare, vad skall jag göra för att få evigt liv till arvedel?»
Då sade han till honom: »Vad är skrivet i lagen?
Huru läser du?»
Han svarade och sade: »'Du skall älska Herren, din Gud, av allt ditt hjärta och av all din själ och av all din kraft och av allt ditt förstånd och din nästa såsom dig själv.'»
Han sade till honom: »Rätt svarade du.
Gör det, så får du leva,
Då ville han rättfärdiga sig och sade till Jesus: »Vilken är då min nästa?»
Jesus svarade och sade: »En man begav sig från Jerusalem ned till Jeriko, men råkade ut för rövare, som togo ifrån honom hans kläder och därtill slogo honom; därefter gingo de sin väg och läto honom ligga där halvdöd.
Så hände sig att en präst färdades samma väg; och när han fick se honom, gick han förbi.
Likaledes ock en levit: när denne kom till det stället och fick se honom, gick han förbi.
Men en samarit, som färdades samma väg, kom också dit där han låg; och när denne fick se honom, ömkade han sig över honom
och gick fram till honom och göt olja och vin i hans sår och förband dem.
Sedan lyfte han upp honom på sin åsna och förde honom till ett härbärge och skötte honom.
Morgonen därefter tog han fram två silverpenningar och gav dem åt värden och sade: 'Sköt honom och vad du mer kostar på honom skall jag betala dig, när jag kommer tillbaka.' --
Vilken av dessa tre synes dig nu hava visat sig vara den mannens nästa, som hade fallit i rövarhänder?»
Han svarade: »Den som bevisade honom barmhärtighet.»
Då sade Jesus till honom: »Gå du och gör sammalunda.»
När de nu voro på vandring, gick han in i en by, och en kvinna, vid namn Marta, tog emot honom i sitt hus.
Och hon hade en syster, som hette Maria; denna satte sig ned vid Herrens fötter och hörde på hans ord.
Men Marta var upptagen av mångahanda bestyr för att tjäna honom.
Och hon gick fram och sade: »Herre, frågar du icke efter att min syster har lämnat alla bestyr åt mig allena?
Säg nu till henne att hon hjälper mig.»
Då svarade Herren och sade till henne: »Marta, Marta, du gör dig bekymmer och oro för mångahanda,
men allenast ett är nödvändigt.
Maria har utvalt den goda delen, och den skall icke tagas ifrån henne.»
När han en gång uppehöll sig på ett ställe för att bedja och hade slutat sin bön, sade en av hans lärjungar till honom: »Herre, lär oss att bedja, såsom ock Johannes lärde sina lärjungar.»
Då sade han till dem: »När I bedjen, skolen I säga så: 'Fader, helgat varde ditt namn; tillkomme ditt rike;
vårt dagliga bröd giv oss var dag;
och förlåt oss våra synder, ty också vi förlåta var och en som är oss något skyldig; och inled oss icke i frestelse.'»
Ytterligare sade han till dem: »Om någon av eder har en vän och mitt i natten kommer till denne och säger till honom: 'Käre vän, låna mig tre bröd;
ty en av mina vänner har kommit resande till mig, och jag har intet att sätta fram åt honom'
så svarar kanske den andre inifrån huset och säger: 'Gör mig icke omak; dörren är redan stängd, och både jag och mina barn hava gått till sängs; jag kan icke stå upp och göra dig något.'
Men jag säger eder: Om han än icke, av det skälet att han är hans vän, vill stå upp och giva honom något, så kommer han likväl, därför att den andre är så påträngande, att stå upp och giva honom så mycket han behöver.
Likaså säger jag till eder: Bedjen, och eder skall varda givet; söken, och I skolen finna; klappen, och för eder skall varda upplåtet.
Ty var och en som beder, han får; och den som söker, han finner; och för den som klappar skall varda upplåtet.
Finnes bland eder någon fader, som när hans son beder honom om en fisk, i stallet för en fisk räcker honom en orm,
eller som räcker honom en skorpion, när han beder om ett ägg?
Om nu I, som ären onda, förstån att giva edra barn goda gåvor, huru mycket mer skall icke då den himmelske Fadern giva helig ande åt dem som bedja honom!»
Och han drev ut en ond ande som var dövstum.
Och när den onde anden hade blivit utdriven, talade den dövstumme; och folket förundrade sig.
Men några av dem sade: »Det är med Beelsebul, de onda andarnas furste, som han driver ut de onda andarna.»
Och några andra ville sätta honom på prov och begärde av honom ett tecken från himmelen.
Men han förstod deras tankar och sade till dem: »Vart rike som har kommit i strid med sig självt bliver förött, så att hus faller på hus.
Om nu Satan har kommit i strid med sig själv, huru kan då hans rike hava bestånd?
I sägen ju att det är med Beelsebul som jag driver ut de onda andarna.
Men om det är med Beelsebul som jag driver ut de onda andarna, med vem driva då edra egna anhängare ut dem?
De skola alltså vara edra domare.
Om det åter är med Guds finger som jag driver ut de onda andarna, så har ju Guds rike kommit till eder. --
När en stark man, fullt väpnad, bevakar sin gård, då äro hans ägodelar fredade.
Men om någon som är starkare än han angriper honom och övervinner honom, så tager denne ifrån honom alla vapnen, som han förtröstade på, och skiftar ut bytet efter honom.
Den som icke är med mig, han är emot mig, och den som icke församlar med mig, han förskingrar.
När en oren ande har farit ut ur en människa, vandrar han omkring i ökentrakter och söker efter ro.
Men då han icke finner någon, säger han: 'Jag vill vända tillbaka till mitt hus, som jag gick ut ifrån.'
Och när han kommer dit och finner det fejat och prytt,
då går han åstad och tager med sig sju andra andar, som äro värre än han själv, och de gå ditin och bo där; och så bliver för den människan det sista värre än det första.»
När han sade detta, hov en kvinna in folkhopen upp sin röst och ropade till honom: »Saligt är det moderssköte som har burit dig, och de bröst som du har diat.»
Men han svarade: »Ja, saliga är de som höra Guds ord och gömma det.»
Men när folket strömmade till tog han till orda och sade: »Detta släkte är ett ont släkte Det begär ett tecken, men intet annat tecken skall givas det än Jonas' tecken.
Ty såsom Jonas blev ett tecken för nineviterna, så skall ock Människosonen vara ett tecken för detta släkte.
Drottningen av Söderlandet skall vid domen träda fram tillsammans med detta släktes män och bliva dem till dom.
Ty hon kom från jordens ända för att höra Salomos visdom; och se, har är vad som är mer än Salomo.
Ninevitiska män skola vid domen träda fram tillsammans med detta släkte och bliva det till dom.
Ty de gjorde bättring vid Jonas' predikan; och se, här är vad som är mer än Jonas.
Ingen tänder ett ljus och sätter det på en undangömd plats eller under skäppan, utan man sätter det på ljusstaken, för att de som komma in skola se skenet.
Ditt öga är kroppens lykta.
När ditt öga är friskt, då har ock hela din kropp ljus; men när det är fördärvat, då är ock din kropp höljd i mörker.
Se därför till, att ljuset som du har i dig icke är mörker.
Om så hela din kropp får ljus och icke har någon del höljd i mörker, då har den ljus i sin helhet, såsom när en lykta lyser dig med sitt klara sken.»
Under det att han så talade, inbjöd en farisé honom till måltid hos sig; och han gick ditin och tog plats vid bordet.
Men när fariséen såg att han icke tvådde sig före måltiden, förundrade han sig.
Då sade Herren till honom: »I fariséer, I gören nu det yttre av bägaren och fatet rent, medan edert inre är fullt av rofferi och ondska.
I dårar, har icke han som har gjort det yttre också gjort det inre?
Given fastmer såsom allmosa vad inuti kärlet är; först då bliver allt hos eder rent.
Men ve eder, I fariséer, som given tionde av mynta och ruta och alla slags kryddväxter, men icke akten på rätten och på kärleken till Gud!
Det ena borden I göra, men icke underlåta det andra.
Ve eder, I fariséer, som gärna viljen sitta främst i synagogorna och gärna viljen bliva hälsade på torgen!
Ve eder, I som ären lika gravar som ingen kan märka, och över vilka människorna gå fram utan att veta det!»
Då tog en av de lagkloke till orda och sade till honom: »Mästare, när du så talar, skymfar du också oss.»
Han svarade: »Ja, ve ock eder, I lagkloke, som på människorna läggen bördor, svåra att bära, men själva icke viljen med ett enda finger röra vid de bördorna!
Ve eder, I som byggen upp profeternas gravar, deras som edra fäder dräpte!
Så bären I då vittnesbörd om edra fäders gärningar och gillen dem; ty om de dräpte profeterna, så byggen I upp deras gravar.
Därför har ock Guds vishet sagt: 'Jag skall sända till dem profeter och apostlar, och somliga av dem skola de dräpa, och andra skola de förfölja.
Och så skall av detta släkte utkrävas alla profeters blod, allt det som är utgjutet från världens begynnelse,
ända ifrån Abels blod intill Sakarias' blod, hans som förgjordes mellan altaret och templet.'
Ja, jag säger eder: Det skall utkrävas av detta släkte.
Ve eder, I lagkloke, som haven tagit bort nyckeln till kunskapen!
Själva haven I icke kommit ditin och för dem som ville komma dit haven I lagt hinder.»
När han inför allt folket sade detta till dem, blevo fariséerna och de lagkloke mycket förbittrade och gåvo sig i strid med honom om många stycken;
de sökte nämligen efter tillfälle att kunna anklaga honom.
Då nu otaligt mycket folk var församlat omkring honom, så att de trampade på varandra, tog han till orda och sade, närmast till sina lärjungar: »Tagen eder till vara för fariséernas surdeg, det är för skrymteri.
Intet är förborgat, som icke skall bliva uppenbarat, och intet är fördolt, som icke skall bliva känt.
Därför skall allt vad I haven sagt i mörkret bliva hört i ljuset, och vad I haven viskat i någons öra i kammaren, det skall bliva utropat på taken.
Men jag säger eder, mina vänner: Frukten icke för dem som väl kunna dräpa kroppen, men sedan icke hava makt att göra något mer.
Jag vill lära eder vem I skolen frukta: frukten honom som har makt att, sedan han har dräpt, också kasta i Gehenna.
Ja, jag säger eder: Honom skolen I frukta. --
Säljas icke fem sparvar för två skärvar?
Och icke en av dem är förgäten hos Gud.
Men på eder äro till och med huvudhåren allasammans räknade.
Frukten icke; I ären mer värda än många sparvar.
Och jag säger eder: Var och en som bekänner mig inför människorna, honom skall ock Människosonen kännas vid inför Guds änglar.
Men den som förnekar mig inför människorna, han skall ock bliva förnekad inför Guds änglar.
Och om någon säger något mot Människosonen, så skall det bliva honom förlåtet; men den som hädar den helige Ande, honom skall det icke bliva förlåtet.
Men när man drager eder fram inför synagogor och överheter och myndigheter, så gören eder icke bekymmer för huru eller varmed I skolen försvara eder, eller vad I skolen säga;
ty den helige Ande skall i samma stund lära eder vad I skolen säga.»
Och en man i folkhopen sade till honom: »Mästare, säg till min broder att han skiftar arvet med mig.»
Men han svarade honom: »Min vän, vem har satt mig till domare eller skiftesman över eder?»
Därefter sade han till dem: »Sen till, att I tagen eder till vara för allt slags girighet; ty en människas liv beror icke därpå att hon har överflöd på ägodelar.»
Och han framställde för dem en liknelse; han sade: »Det var en rik man vilkens åkrar buro ymniga skördar.
Och han tänkte vid sig själv och sade: 'Vad skall jag göra?
Jag har ju icke rum nog för att inbärga min skörd.'
Därefter sade han: 'Så vill jag göra: jag vill riva ned mina lador och bygga upp större, och i dem skall jag samla in all min gröda och allt mitt goda.
Sedan vill jag säga till min själ: Kära själ, du har mycket gott för varat för många år; giv dig nu ro, ät, drick och var glad.
Men Gud sade till honom: 'Du dåre, i denna natt skall din själ utkrävas av dig; vem skall då få vad du har samlat i förråd?' --
Så går det den som samlar skatter åt sig själv, men icke är rik inför Gud.»
Och han sade till sina lärjungar: »Därför säger jag eder: Gören eder icke bekymmer för edert liv, vad I skolen äta, ej heller för eder kropp, vad I skolen kläda eder med.
Livet är ju mer än maten, och kroppen mer än kläderna.
Given akt på korparna: de så icke, ej heller skörda de, och de hava varken visthus eller lada; och likväl föder Gud dem.
Huru mycket mer ären icke I än fåglarna!
Vilken av eder kan med allt sitt bekymmer lägga en aln till sin livslängd?
Förmån I nu icke ens det som minst är, varför gören I eder då bekymmer för det övriga?
Given akt på liljorna, huru de varken spinna eller väva; och likväl säger jag eder att icke ens Salomo i all sin härlighet var så klädd som en av dem.
Kläder nu Gud så gräset på marken, vilket i dag står och i morgon kastas i ugnen, huru mycket mer skall han då icke kläda eder, I klentrogne!
Söken därför icke heller I efter vad I skolen äta, eller vad I skolen dricka, och begären icke vad som är för högt.
Efter allt detta söka ju hedningarna i världen, och eder Fader vet att I behöven detta.
Nej, söken efter hans rike, så skall också detta andra tillfalla eder.
Frukta icke, du lilla hjord; ty det har behagat eder Fader att giva eder riket.
Säljen vad I ägen och given allmosor; skaffen eder penningpungar som icke nötas ut, en outtömlig skatt i himmelen, dit ingen tjuv når, och där man icke fördärvar.
Ty där eder skatt är, där komma ock edra hjärtan att vara.
Haven edra länder omgjordade och edra lampor brinnande.
Och varen I lika tjänare som vänta på att deras herre skall bryta upp från bröllopet, för att strax kunna öppna för honom, när han kommer och klappar.
Saliga äro de tjänare som deras herre finner vakande, när han kommer.
Sannerligen säger jag eder: Han skall fästa upp sin klädnad och låta dem taga plats vid bordet och själv gå fram och betjäna dem.
Och vare sig han kommer under den andra nattväkten eller under den tredje och finner dem så göra -- saliga äro de då.
Men det förstån I väl, att om husbonden visste vilken stund tjuven skulle komma, så tillstadde han icke att någon bröt sig in i hans hus.
Så varen ock I redo ty i en stund då I icke vänten det skall Människosonen komma.»
Då sade Petrus: »Herre, är det om oss som du talar i denna liknelse, eller är det om alla?»
Herren svarade: »Finnes någon trogen och förståndig förvaltare, som av sin herre kan sättas över hans husfolk, för att i rätt tid giva dem deras bestämda kost --
salig är då den tjänaren, om hans herre, när han kommer, finner honom göra så.
Sannerligen säger jag eder: Han skall sätta honom över allt vad han äger.
Men om så är, att tjänaren säger i sitt hjärta: 'Min herre kommer icke så snart', och han begynner att slå de andra tjänarna och tjänarinnorna och att äta och dricka så att han bliver drucken,
då skall den tjänarens herre komma på en dag då han icke väntar det, och i en stund då han icke tänker sig det, och han skall låta hugga honom i stycken och låta honom få sin del med de otrogna. --
Och den tjänare som hade fått veta sin herres vilja, men icke redde till eller gjorde efter hans vilja, han skall bliva straffad med många slag.
Men den som, utan att hava fått veta hans vilja, gjorde vad som val slag värt, han skall bliva straffad med allenast få slag.
Var och en åt vilken mycket är givet, av honom skall mycket varda utkrävt och den som har blivit betrodd med mycket, av honom skall man fordra dess mera.
Jag har kommit för att tända en eld på jorden; och huru gärna ville jag icke att den redan brunne!
Men jag måste genomgå ett dop; och huru ängslas jag icke, till dess att det är fullbordat!
Menen I att jag har kommit för att skaffa frid på jorden?
Nej, säger jag eder, fastmer söndring.
Ty om fem finnas i samma hus, skola de härefter vara söndrade från varandra, så att tre stå mot två Och två mot tre:
fadern mot sin son och sonen mot sin fader, modern mot sin dotter och dottern mot sin moder, svärmodern mot sin sonhustru och sonhustrun mot sin svärmoder.
Han hade också till folket: »När I sen ett moln stiga upp i väster, sägen I strax: 'Nu kommer regn'; och det sker så.
Och när I sen sunnanvind blåsa, sägen I: 'Nu kommer stark hetta'; och detta sker.
I skrymtare, jordens och himmelens utseende förstån I att tyda; huru kommer det då till, att I icke kunnen tyda denna tiden?
Varför låten I icke edert eget inre döma om vad rätt är?
När du går till en överhetsperson med din motpart, så gör dig under vägen all möda att bliva förlikt med denne, så att han icke drager dig fram inför domaren; då händer att domaren överlämnar dig åt rättstjänaren, och att rättstjänaren kastar dig i fängelse.
Jag säger dig: Du skall icke slippa ut därifrån, förrän du har betalt ända till den yttersta skärven.»
Vid samma tid kommo några och berättade för honom om de galiléer vilkas blod Pilatus hade blandat med deras offer.
Då svarade han och sade till dem: »Menen I att dessa galiléer voro större syndare än alla andra galiléer, eftersom de fingo lida sådant?
Nej, säger jag eder; men om I icke gören bättring, skolen I alla sammalunda förgås.
Eller de aderton som dödades, när tornet i Siloam föll på dem, menen I att de voro mer brottsliga än alla andra människor som bo i Jerusalem?
Nej, säger jag eder; men om I icke gören bättring, skolen I alla sammalunda förgås.»
Och han framställde denna liknelse: »En man hade ett fikonträd planterat i sin vingård; och han kom och sökte frukt därpå, men fann ingen.
Då sade han till vingårdsmannen: 'Se, nu i tre år har jag kommit och sökt frukt på detta fikonträd, utan att finna någon.
Hugg bort det.
Varför skall det därjämte få utsuga jorden?'
Men vingårdsmannen svarade och sade till honom: 'Herre, låt det stå kvar också detta år, för att jag under tiden må gräva omkring det och göda det;
kanhända skall det så till nästa å bära frukt.
Varom icke, så må du då hugga bort det.'»
När han en gång på sabbaten undervisade i en synagoga,
var där en kvinna som i aderton år hade varit besatt av en sjukdomsande, och hon var så hopkrumpen, att hon alls icke kunde räta upp sin kropp.
Då nu Jesus fick se henne, kallade han henne till sig och sade till henne »Kvinna, du är fri ifrån din sjuk dom»,
och han lade därvid händerna på henne.
Och strax rätade hon upp sig och prisade Gud.
Men det förtröt synagogföreståndaren att Jesus på sabbaten botade sjuka; och han tog till orda och sade till folket: »Sex dagar finnas, på vilka man bör arbeta.
På dem mån I alltså komma och låta bota eder, men icke på sabbatsdagen.
Då svarade Herren honom och sade: »I skrymtare, löser icke var och en av eder på sabbaten sin oxe eller åsna från krubban och leder den bort för att vattna den?
Och denna kvinna, en Abrahams dotter, som Satan har hållit bunden nu i aderton år, skulle då icke hon på sabbatsdagen få lösas från sin boja?»
När han sade detta, blygdes alla hans motståndare; och allt folket gladde sig över alla de härliga gärningar som gjordes av honom.
Så sade han då: »Vad är Guds rike likt, ja, vad skall jag likna det vid?
Det är likt ett senapskorn som en man tager och lägger ned i sin trädgård, och det växer och bliver ett träd, och himmelens fåglar bygga sina nästen på dess grenar.»
Ytterligare sade han: »Vad skall jag likna Guds rike vid?
Det är likt en surdeg som en kvinna tager och blandar in i tre skäppor mjöl, till dess alltsammans bliver syrat.»
Och han vandrade från stad till stad och från by till by och undervisade folket, under det att han fortsatte sin färd till Jerusalem.
Och någon frågade honom: »Herre, är det allenast få som bliva frälsta?»
Då svarade han dem:
»Kämpen för att komma in genom den trånga dörren; ty många, säger jag eder, skola försöka att komma in och skola dock icke förmå det.
Om husbonden har stått upp och tillslutit dörren, och I sedan kommen och ställen eder därutanför och klappen på dörren och sägen: 'Herre, låt upp för oss', så skall han svara och säga till eder: 'Jag vet icke varifrån I ären.'
Och I skolen då säga: 'Vi hava ju ätit och druckit med dig, och du har undervisat på våra gator.'
Men han skall svara: 'Jag säger eder: Jag vet icke varifrån I ären; gån bort ifrån mig, alla I ogärningsmän.'
Där skall då bliva gråt och tandagnisslan, när I fån se Abraham, Isak och Jakob och alla profeterna vara i Guds rike, men finnen eder själva utkastade.
Ja, människor skola komma från öster och väster, från norr och söder och bliva bordsgäster i Guds rike.
Och se, då skola somliga som äro de sista bliva de första, och somliga som äro de första bliva de sista.
I samma stund kommo några fariséer fram och sade till honom: »Begiv dig åstad bort härifrån; ty Herodes vill dräpa dig.»
Då svarade han dem: »Gån och sägen den räven, att jag i dag och i morgon driver ut onda andar och botar sjuka, och att jag först på tredje dagen är färdig.
Men jag måste vandra i dag och i morgon och i övermorgon, ty det är icke i sin ordning att en profet förgöres annorstädes än i Jerusalem. --
Jerusalem, Jerusalem, du som dräper profeterna och stenar dem som äro sända till dig!
Huru ofta har jag icke velat församla dina barn, likasom hönan församlar sina kycklingar under sina vingar!
Men haven icke velat.
Se, edert hus skall komma att stå övergivet.
Men jag säger eder: I skolen icke se mig, förrän den tid kommen, då I sägen: 'Välsignad vare han som kommer, i Herrens namn.'
När han på en sabbat hade kommit in till en av de förnämligaste fariséerna för att intaga en måltid, hände sig, medan man där vaktade på honom,
att en vattusiktig man kom dit och stod framför honom.
Då tog Jesus till orda och sade till de lagkloke och fariséerna: »Är det lovligt att bota sjuka på sabbaten, eller är det icke lovligt?»
Men de tego.
Då tog han mannen vid handen och gjorde honom frisk och lät honom gå.
Sedan sade han till dem: »Om någon av eder har en åsna eller en oxe som faller i en brunn, går han icke då strax och drager upp den, jämväl på sabbatsdagen?»
Och de förmådde icke svara något härpå.
Då han nu märkte huru gästerna utvalde åt sig de främsta platserna, framställde han för dem en liknelse; han sade till dem:
»När du av någon har blivit bjuden till bröllop, så tag icke den främsta platsen vid bordet.
Ty kanhända finnes bland gästerna någon som är mer ansedd än du,
och då kommer till äventyrs den som har bjudit både dig och honom och säger till dig: 'Giv plats åt denne'; och så måste du med skam intaga den nedersta platsen.
Nej, när du har blivit bjuden, så gå och tag den nedersta platsen vid bordet.
Ty det kan då hända att den som har bjudit dig säger till dig, när han kommer: 'Min vän, stig högre upp.'
Då vederfares dig heder inför alla de andra bordsgästerna.
Ty var och en som upphöjer sig, han skall bliva förödmjukad, och den som ödmjukar sig, han skall bliva upphöjd.»
Han sade ock till den som hade bjudit honom: »När du gör ett gästabud, på middagen eller på aftonen, så inbjud icke dina vänner eller dina bröder eller dina fränder, ej heller rika grannar, så att de bjuda dig igen och du därigenom får vedergällning.
Nej, när du gör gästabud, så bjud fattiga, krymplingar, halta, blinda.
Salig är du då; ty eftersom de icke förmå vedergälla dig, skall du få din vedergällning vid de rättfärdigas uppståndelse.»
Då nu en av de andra vid bordet hörde detta, sade denne till honom: »Salig är den som får bliva bordsgäst i Guds rike!»
Då sade han till honom: »En man tillredde ett stort gästabud och bjöd många.
Och när gästabudet skulle hållas, sände han ut sin tjänare och lät säga till dem som voro bjudna: 'Kommen, ty nu är allt redo.'
Men de begynte alla strax ursäkta sig.
Den förste sade till honom: 'Jag har köpt ett jordagods, och jag måste gå ut och bese det.
Jag beder dig, tag emot min ursäkt.'
En annan sade: 'Jag har köpt fem par oxar, och jag skall nu gå åstad och försöka dem.
Jag beder dig, tag emot min ursäkt.'
Åter en annan sade: 'Jag har tagit mig hustru, och därför kan jag icke komma.'
Och tjänaren kom igen och omtalade detta för sin herre.
Då blev husbonden vred och sade till sin tjänare: 'Gå strax ut på gator och gränder i staden, och för hitin fattiga och krymplingar och blinda och halta.'
Sedan sade tjänaren: 'Herre, vad du befallde har blivit gjort, men har är ännu rum.'
Då sade herren till tjänaren: 'Gå ut på vägar och stigar, och nödga människorna att komma hitin, så att mitt hus bliver fullt.
Ty jag säger eder att ingen av de män som voro bjudna skall smaka sin måltid.'»
Och mycket folk gick med honom; och han vände sig om och sade till dem:
»Om någon kommer till mig, och han därvid ej hatar sin fader och sin moder, och sin hustru och sina barn, och sina bröder och systrar, därtill ock sitt eget liv, så kan han icke vara min lärjunge.
Den som icke bär sitt kors och efterföljer mig, han kan icke vara min lärjunge.
Ty om någon bland eder vill bygga ett torn, sätter han sig icke då först ned och beräknar kostnaden och mer till, om han äger vad som behöves för att bygga det färdigt?
Eljest, om han lade grunden, men icke förmådde fullborda verket skulle ju alla som finge se det begynna att begabba honom
och säga: 'Den mannen begynte bygga, men förmådde icke fullborda sitt verk.'
Eller om en konung vill draga ut i krig för att drabba samman med en annan konung, sätter han sig icke då först ned och tänker efter, om han förmår att med tio tusen möta den som kommer emot honom med tjugu tusen?
Om så icke är, måste han ju, medan den andre ännu är långt borta, skicka sändebud och underhandla om fred.
Likaså kan ingen av eder vara min lärjunge, om han icke försakar allt vad han äger. --
Så är väl saltet en god sak, men om till och med saltet mister sin sälta, varmed skall man då återställa dess kraft?
Varken för jorden eller för gödselhögen är det tjänligt; man kastar ut det.
Den som har öron till att höra, han höre.»
Och till honom kom allt vad publikaner och syndare hette för att höra honom.
Men fariséerna och de skriftlärde knorrade och sade: »Denne tager emot syndare och äter med dem.»
Då framställde han för dem denna liknelse; han sade:
»Om ibland eder finnes en man som har hundra får, och han förlorar ett av dem, lämnar han icke då de nittionio i öknen och går och söker efter det förlorade, till dess han finner det?
Och när han har funnit det, lägger han det på sina axlar med glädje.
Och när han kommer hem, kallar han tillhopa sina vänner och grannar och säger till dem: 'Glädjens med mig, ty jag har funnit mitt får, som var förlorat.'
Jag säger eder att likaså bliver mer glädje i himmelen över en enda syndare som gör bättring, än över nittionio rättfärdiga som ingen bättring behöva.
Eller om en kvinna har tio silverpenningar, och hon tappar bort en av dem, tänder hon icke då upp ljus och sopar huset och söker noga, till dess hon finner den?
Och när hon har funnit den, kallar hon tillhopa sina väninnor och grannkvinnor och säger: 'Glädjens med mig, ty jag har funnit den penning som jag hade tappat bort.'
Likaså, säger jag eder, bliver glädje hos Guds änglar över en enda syndare som gör bättring.
Ytterligare sade han: »En man hade två söner.
Och den yngre av dem sade till fadern: 'Fader, giv mig den del av förmögenheten, som faller på min lott.'
Då skiftade han sina ägodelar mellan dem.
Och icke lång tid därefter lade den yngre sonen allt sitt tillhopa och for långt bort till ett främmande land.
Där levde han i utsvävningar och förfor så sin förmögenhet.
Men sedan han hade slösat bort allt, kom en svär hungersnöd över det landet, och han begynte lida nöd.
Då gick han bort och gav sig under en man där i landet, och denne sände honom ut på sina marker för att vakta svin.
Och han åstundade att få fylla sin buk med de fröskidor som svinen åto; men ingen gav honom något.
Då kom han till besinning och sade: 'Huru många legodrängar hos min fader hava icke bröd i överflöd, medan jag har förgås av hunger!
Jag vill stå upp och gå till min fader och säga till honom: Fader, jag har syndat mot himmelen och inför dig;
jag är icke mer värd att kallas din son.
Låt mig bliva såsom en av dina legodrängar.'
Så stod han upp och gick till sin fader.
Och medan han ännu var långt borta, fick hans fader se honom och ömkade sig över honom och skyndade emot honom och föll honom om halsen och kysste honom innerligt.
Men sonen sade till honom: 'Fader, jag har syndat mot himmelen och inför dig; jag är icke mer värd att kallas din son.'
Då sade fadern till sina tjänare 'Skynden eder att taga fram den yppersta klädnaden och kläden honom i den, och sätten en ring på hans hand och skor på hans fötter.
Och hämten den gödda kalven och slakten den, så vilja vi äta och gör oss glada.
Ty denne min son var död, men har fått liv igen; han var förlorad men är återfunnen.'
Och de begynte göra sig glada.
Men hans äldre son var ute på marken.
När denne nu vände tillbaka och hade kommit nära huset fick han höra spel och dans.
Då kallade han till sig en av tjänarna och frågade vad detta kunde betyda.
Denne svarade honom: 'Din broder har kommit hem; och då nu din fader har fått honom välbehållen tillbaka, har han låtit slakta den gödda kalven.'
Då blev han vred och ville icke gå in.
Hans fader gick då ut och talade vanligt med honom.
Men han svarade och sade till sin fader: 'Se, i så många år har jag nu tjänat dig, och aldrig har jag överträtt något ditt bud; och lik väl har du åt mig aldrig givit ens en killing, för att jag skulle kunna göra mig glad med mina vänner.
Men när denne din son, som har förtärt dina ägodelar tillsammans med skökor, nu har kommit tillbaka, så har du för honom låtit slakta den gödda kalven.'
Då sade han till honom: 'Min son, du är alltid hos mig, och all mitt är ditt.
Men nu måste vi fröjda oss och vara glada; ty denne din broder var död, men har fått liv igen, han var förlorad, men är återfunnen.'»
Han sade också till sina lärjungar: »En rik man hade en förvaltare som hos honom blev angiven för förskingring av hans ägodelar.
Då kallade han honom till sig och sade till honom: 'Vad är det jag hör om dig?
Gör räkenskap för din förvaltning; ty du kan icke längre få vara förvaltare.'
Men förvaltaren sade vid sig själv: 'Vad skall jag göra, då min herre nu tager ifrån mig förvaltningen?
Gräva orkar jag icke; att tigga blyges jag för.
Dock, nu vet jag vad jag skall göra, för att man må upptaga mig i sina hus, när jag bliver avsatt ifrån förvaltningen.'
Och han kallade till sig sin herres gäldenärer, var och en särskilt.
Och han frågade den förste: 'Huru mycket är du skyldig min herre?'
Han svarade: 'Hundra fat olja.'
Då sade han till honom: 'Tag här ditt skuldebrev, och sätt dig nu strax ned och skriv femtio.'
Sedan frågade han en annan: 'och du, huru mycket är du skyldig?'
Denne svarade: 'hundra tunnor vete.'
Då sade han till honom: 'Tag här ditt skuldebrev och skriv åttio.'
Och husbonden prisade den orättrådige förvaltaren för det att han hade handlat klokt.
Ty denna tidsålders barn skicka sig klokare mot sitt släkte än ljusets barn.
Och jag säger eder: Skaffen eder vänner medelst den orättrådige Mamons goda, för att de, när detta har tagit slut, må taga emot eder i de eviga hyddorna.
Den som är trogen i det minsta, han är ock trogen i vad mer är, och den som är orättrådig i det minsta, han är ock orättrådig i vad mer är.
Haven I nu icke varit trogna, när det gällde den orättrådige Mamons goda, vem vill då betro eder det sannskyldiga goda?
Och haven I icke varit trogna, när det gällde vad som tillhörde en annan, vem vill då giva eder det som hör eder till?
Ingen som tjänar kan tjäna två herrar; ty antingen kommer han då att hata den ene och älska den andre, eller kommer han att hålla sig till den förre och förakta den senare.
I kunnen icke tjäna både Gud och Mamon.»
Allt detta hörde nu fariséerna, som voro penningkära, och de drevo då gäck med honom.
Men han sade till dem: »I hören till dem som göra sig rättfärdiga inför människorna.
Men Gud känner edra hjärtan; ty det som bland människor är högt är en styggelse inför Gud.
Lagen och profeterna hava haft sin tid intill Johannes.
Sedan dess förkunnas evangelium om Guds rike, och var man vill storma ditin.
Men snarare kunna himmel och jord förgås, än en enda prick av lagen kan falla bort.
Var och en som skiljer sig från sin hustru och tager sig en annan hustru, han begår äktenskapsbrott.
Och den som tager till hustru en kvinna som är skild från sin man, han begår äktenskapsbrott.
Det var en rik man som klädde sig i purpur och fint linne och levde var dag i glädje och prakt.
Men en fattig man, vid namn Lasarus, låg vid hans port, full av sår,
och åstundade att få stilla sin hunger med vad som kunde falla ifrån den rike mannens bord.
Ja, det gick så långt att hundarna kommo och slickade hans sår.
Så hände sig att den fattige dog och blev förd av änglarna till Abrahams sköte.
Också den rike dog och blev begraven.
När han nu låg i dödsriket och plågades, lyfte han upp sina ögon och fick se Abraham långt borta och Lasarus i hans sköte.
Då ropade han och sade: 'Fader Abraham, förbarma dig över mig, och sänd Lasarus att doppa det yttersta av sitt finger i vatten och svalka min tunga, ty jag pinas svårt i dessa lågor.'
Men Abraham svarade: 'Min son kom ihåg att du, medan du levde, fick ut ditt goda och Lasarus däremot vad ont var; nu åter får han här hugnad, under det att du pinas.
Och till allt detta kommer, att ett stort svalg är satt mellan oss och eder, för att de som vilja begiva sig över härifrån till eder icke skola kunna det, och för att ej heller någon därifrån skall kunna komma över till oss.»
Då sade han: 'Så beder jag dig då, fader, att du sänder honom till min faders hus,
där jag har fem bröder, och låter honom varna dem, så att icke också de komma till detta pinorum.'
Men Abraham sade: 'De hava Moses och profeterna; dem må de lyssna till.'
Han svarade: 'Nej, fader Abraham; men om någon kommer till dem från de döda, så skola de göra bättring.'
Då sade han till honom: 'Lyssna de icke till Moses och profeterna, så skola de icke heller låta övertyga sig, om någon uppstår från de döda.'»
Och han sade till sina lärjungar: »Det är icke annat möjligt än att förförelser måste komma, men ve den genom vilken de komma!
För honom vore det bättre att en kvarnsten hängdes om hans hals och han kastades i havet, än att han skulle förföra en av dessa små.
Tagen eder till vara!
Om din broder försyndat sig, så tillrättavisa honom; och om han då ångrar sig, så förlåt honom.
Ja, om han sju gånger om dagen försyndar sig mot dig och sju gånger kommer tillbaka till dig och säger: 'Jag ångrar mig' så skall du förlåta honom.»
Och apostlarna sade till Herren: »Föröka vår tro.»
Då sade Herren: »Om I haden tro, vore den ock blott såsom ett senapskorn, så skullen I kunna säga till detta mullbärsfikonträd: 'Ryck dig upp med rötterna, och plantera dig i havet', och det skulle lyda eder.
Om någon bland eder har en tjänare som kör plogen eller vaktar boskap, icke säger han väl till tjänaren, när denne kommer hem från marken: 'Gå du nu strax till bords'?
Säger han icke fastmer till honom: 'Red till min måltid, och fäst så upp din klädnad och betjäna mig, medan jag äter och dricker; sedan må du själv äta och dricka'?
Icke tackar han väl tjänaren för att denne gjorde det som blev honom befallt?
Sammalunda, när I haven gjort allt som har blivit eder befallt, då skolen I säga: 'Vi äro blott ringa tjänare: vi hava endast gjort vad vi voro pliktiga att göra.'»
Då han nu var stadd på sin färd till Jerusalem, tog han vägen mellan Samarien och Galileen.
Och när han kom in i en by, möttes han av tio spetälska män.
Dessa stannade på avstånd
och ropade och sade: »Jesus, Mästare, förbarma dig över oss.»
När han fick se dem, sade han till dem: »Gån och visen eder för prästerna.»
Och medan de voro på väg dit, blevo de rena.
Och en av dem vände tillbaka, när han såg att han hade blivit botad, och prisade Gud med hög röst
och föll ned på mitt ansikte för Jesu fötter och tackade honom.
Och denne var en samarit.
Då svarade Jesus och sade: »Blevo icke alla tio gjorda rena?
Var äro de nio?
Fanns då ibland dem ingen som vände tillbaka för att prisa Gud, utom denne främling?»
Och han sade till honom: »Stå upp och gå dina färde.
Din tro har frälst dig.»
Och då han blev tillfrågad av fariséerna när Guds rike skulle komma, svarade han dem och sade: »Guds rike kommer icke på sådant sätt att det kan förnimmas med ögonen,
ej heller skall man kunna säga: 'Se här är det', eller: 'Där är det.'
Ty se, Guds rike är invärtes i eder.»
Och han sade till lärjungarna: »Den tid skall komma, då I gärna skullen vilja se en av Människosonens dagar, men I skolen icke få det.
Väl skall man då säga till eder: 'Se där är han', eller: 'Se här är han'; men gån icke dit, och löpen icke därefter.
Ty såsom ljungelden, när den ljungar fram, lyser från himmelens ena ända till den andra, så skall det vara med Människosonen på hand dag.
Men först måste han lida mycket och bliva förkastad av detta släkte.
Och såsom det skedde på Noas tid, så skall det ock ske i Människosonens dagar:
människorna åto och drucko, män togo sig hustrur, och hustrur gåvos åt män, ända till den dag då Noa gick in i arken; då kom floden och förgjorde dem allasammans.
Likaledes, såsom det skedde på Lots tid: människorna åto och drucko, köpte och sålde, planterade och byggde,
men på den dag då Lot gick ut från Sodom regnade eld och svavel ned från himmelen och förgjorde dem allasammans,
alldeles på samma sätt skall det ske den dag då Människosonen uppenbaras.
Den som den dagen är på taket och har sitt bohag inne i huset, han må icke stiga ned för att hämta det; ej heller må den som är ute på marken vända tillbaka.
Kommen ihåg Lots hustru.
Den som står efter att vinna sitt liv, han skall mista det; men den som mister det, han skall rädda det.
Jag säger eder: Den natten skola två ligga i samma säng; den ene skall bliva upptagen, den andre skall lämnas kvar.
Två kvinnor skola mala tillhopa; den ena skall bliva upptagen, den andra skall lämnas kvar.»
Då frågade de honom: »Var då, Herre?»
Han svarade dem: »Där den döda kroppen är, dit skola ock rovfåglarna församla sig.»
Och han framställde för dem en liknelse, för att lära dem att de alltid borde bedja, utan att förtröttas.
Han sade: »I en stad fanns en domare som icke fruktade Gud och ej heller hade försyn för någon människa.
I samma stad fanns ock en änka som åter och åter kom till honom och sade: 'Skaffa mig rätt av min motpart.'
Till en tid ville han icke.
Men omsider sade han vid sig själv: 'Det må nu vara, att jag icke fruktar Gud och ej heller har försyn för någon människa;
likväl, eftersom denna änka är mig så besvärlig, vill jag ändå skaffa henne rätt, för att hon icke med sina ideliga besök skall alldeles pina ut mig.'»
Och Herren tillade: »Hören vad den orättfärdige domaren här säger.
Skulle då Gud icke skaffa rätt åt sina utvalda, som ropa till honom dag och natt, och skulle han icke hava tålamod med dem?
Jag säger eder: Han skall snart skaffa dem rätt.
Men skall väl Människosonen, när han kommer, finna tro här på jorden?»
Ytterligare framställde han denna liknelse för somliga som förtröstade på sig själva och menade sig vara rättfärdiga, under det att de föraktade andra:
»Två män gingo upp i helgedomen för att bedja; den ene var en farisé och den andre en publikan.
Fariséen trädde fram och bad så för sig själv: 'Jag tackar dig, Gud, för att jag icke är såsom andra människor, rövare, orättrådiga, äktenskapsbrytare, ej heller såsom denne publikan.
Jag fastar två gånger i veckan; jag giver tionde av allt vad jag förvärvar.'
Men publikanen stod långt borta och ville icke ens lyfta sina ögon upp mot himmelen, utan slog sig för sitt bröst och sade: 'Gud, misskunda dig över mig syndare.' --
Jag säger eder: Denne gick hem igen rättfärdig mer an den andre.
Ty var och en som upphöjer sig, han skall bliva förödmjukad, men den som ödmjukar sig, han skall bliva upphöjd.»
Man bar fram till honom också späda barn, för att han skulle röra vid dem; men när hans lärjungar sågo detta, visade de bort dem.
Då kallade Jesus barnen till sig, i det han sade: »Låten barnen komma till mig, och förmenen dem det icke; ty Guds rike hör sådana till.
Sannerligen säger jag eder: Den som icke tager emot Guds rike såsom ett barn, han kommer aldrig ditin.»
Och en överhetsperson frågade honom och sade: »Gode Mästare, vad skall jag göra för att få evigt liv till arvedel?»
Jesus sade till honom: »Varför kallar du mig god?
Ingen är god utom Gud allena.
Buden känner du: 'Du skall icke begå äktenskapsbrott', 'Du skall icke dräpa', 'Du skall icke stjäla', 'Du skall icke bära falskt vittnesbörd', 'Hedra din fader och din moder.'»
Då svarade han: »Allt detta har jag hållit från min ungdom.»
När Jesus hörde detta, sade han till honom: »Ett återstår dig ännu: sälj allt vad du äger och dela ut åt de fattiga; då skall du få en skatt i himmelen.
Och kom sedan och följ mig.»
Men när han hörde detta, blev han djupt bedrövad, ty han var mycket rik.
Då nu Jesus såg huru det var med honom, sade han: »Huru svårt är det icke för dem som hava penningar att komma in i Guds rike!
Ja, det är lättare för en kamel att komma in genom ett nålsöga, än för den som är rik att komma in i Guds rike.»
Då sade de som hörde detta: »Vem kan då bliva frälst?»
Men han svarade: »Vad som är omöjligt för människor, det är möjligt för Gud.»
Då sade Petrus: »Se, vi hava övergivit allt som var vårt och hava följt dig.»
Han svarade dem: »Sannerligen säger jag eder: Ingen som för Guds rikes skull har övergivit hus, eller hustru, eller bröder, eller föräldrar eller barn,
ingen sådan finnes, som icke skall mångfaldigt igen redan här i tiden, och i den tillkommande tidsåldern evigt liv.»
Och han tog till sig de tolv och sade till dem: »Se, vi gå nu upp till Jerusalem, och allt skall fullbordas, som genom profeterna är skrivet om Människosonen.
Ty han skall bliva överlämnad åt hedningarna och bliva begabbad och skymfad och bespottad,
och de skola gissla honom och döda honom; men på tredje dagen skall han uppstå igen.»
Och de förstodo intet härav; ja, detta som han talade var dem så fördolt, att de icke fattade vad som sades.
Då han nu nalkades Jeriko, hände sig att en blind man satt vid vägen och tiggde.
När denne hörde en hop människor gå där fram, frågade han vad det var.
Och man omtalade för honom att det var Jesus från Nasaret som kom på vägen.
Då ropade han och sade: »Jesus, Davids son, förbarma dig över mig.»
Och de som gingo framför tillsade honom strängeligen att han skulle tiga; men han ropade ännu mycket mer: »Davids son, förbarma dig över mig.»
Då stannade Jesus och bjöd att mannen skulle ledas fram till honom.
Och när han hade kommit fram, frågade han honom:
»Vad vill du att jag skall göra dig?»
Han svarade: »Herre, låt mig få min syn.»
Jesus sade till honom: »Hav din syn; din tro har hjälpt dig.»
Och strax fick han sin syn och följde honom och prisade Gud.
Och allt folket som såg detta lovade Gud.
Och han kom in i Jeriko och gick fram genom staden.
Där fanns en man, vid namn Sackeus, som var förman för publikanerna och en rik man.
Denne ville gärna veta vem som var Jesus och ville se honom, men han kunde det icke för folkets skull, ty han var liten till växten.
Då skyndade han i förväg och steg upp i ett mullbärsfikonträd för att få se honom, ty han skulle komma den vägen fram.
När Jesus nu kom till det stället, såg han upp och sade till honom: »Sackeus, skynda dig ned, ty i dag måste jag gästa i ditt hus.»
Och han skyndade sig ned och tog emot honom med glädje.
Men alla som sågo det knorrade och sade: »Han har gått in för att gästa hos en syndare.»
Men Sackeus trädde fram och sade till Herren: »Herre, hälften av mina ägodelar giver jag nu åt de fattiga; och om jag har utkrävt för mycket av någon, så giver jag fyradubbelt igen.
Och Jesus sade om honom: »I dag har frälsning vederfarits detta hus, eftersom också han är en Abrahams son.
Ty Människosonen har kommit för att uppsöka och frälsa det som var förlorat.»
Medan de hörde härpå, framställde han ytterligare en liknelse, eftersom han var nära Jerusalem och de nu menade att Guds rike strax skulle uppenbaras.
Han sade alltså: »En man av förnämlig släkt tänkte fara bort till ett avlägset land för att utverka åt sig konungslig värdighet; sedan skulle han komma tillbaka.
Och han kallade till sig tio sin tjänare och gav dem tio pund och sade till dem: 'Förvalten dessa, till dess jag kommer tillbaka.'
Men hans landsmän hatade honom och sände, efter hans avfärd, åstad en beskickning och läto säga: 'Vi vilja icke att denne skall bliva konung över oss.»
När han sedan kom tillbaka, efter att hava utverkat åt sig den konungsliga värdigheten, lät han kalla till sig de tjänare åt vilka han hade givit penningarna, ty han ville veta vad var och en genom sin förvaltning hade förvärvat.
Då kom den förste fram och sade: 'Herre, ditt pund har givit i vinst tio pund.'
Han svarade honom: 'Rätt så, du gode tjänare!
Eftersom du har varit trogen i en mycket ringa sak, skall du få makt och myndighet över tio städer.'
Därefter kom den andre i ordningen och sade: 'Herre, ditt pund har avkastat fem pund.'
Då sade han jämväl till denne: 'Så vare ock du satt över fem städer.'
Och den siste kom fram och sade: 'Herre, se här är ditt pund; jag har haft det förvarat i en duk.
Ty jag fruktade för dig, eftersom du är en sträng man; du vill taga upp vad du icke har lagt ned, och skörda vad du icke har sått.'
Han sade till honom: 'Efter dina egna ord vill jag döma dig, du onde tjänare.
Du visste alltså att jag är en sträng man, som vill taga upp vad jag icke har lagt ned, och skörda vad jag icke har sått?
Varför satte du då icke in mina penningar i en bank?
Då hade jag, när jag kom hem, fått uppbära dem med ränta.'
Och han sade till dem som stodo vid hans sida: 'Tagen ifrån honom hans pund, och given det åt den som har de tio punden.'
De sade till honom: 'Herre, han har ju redan tio pund.'
Han svarade: 'Jag säger eder: Var och en som har, åt honom skall varda givet; men den som icke har, från honom skall tagas också det han har.
Men dessa mina ovänner, som icke ville hava mig till konung över sig, fören dem hit huggen ned dem här inför mig.»
Sedan Jesus hade sagt detta, gick han framför de andra upp mot Jerusalem.
När han då nalkades Betfage och Betania, vid det berg som kallas Oljeberget, sände han åstad två av lärjungarna
och sade: »Gån in i byn som ligger här mitt framför.
Och när I kommen ditin, skolen I finna en åsnefåle stå där bunden, som ingen människa någonsin har suttit på, lösen den och fören den hit.
Och om någon frågar eder varför I lösen den skolen I svara så: 'Herren behöver den.'»
Och de som hade blivit utsända gingo åstad och funno det så som han hade sagt dem.
Och när de löste fålen, frågade ägaren dem: »Varför lösen I fålen?»
De svarade: »Herren behöver den.»
Och de förde fålen till Jesus och lade sina mantlar på den och läto Jesus sätta sig därovanpå.
Och där han färdades fram bredde de ut sina mantlar under honom på vägen.
Och då han var nära foten av Oljeberget, begynte hela lärjungaskaran i sin glädje att med hög röst lova Gud för alla de kraftgärningar som de hade sett;
och de sade: »Välsignad vare han som kommer, konungen, i Herrens namn.
Frid vare i himmelen och ära i höjden!»
Och några fariséer som voro med i folkhopen sade till honom: »Mästare, förbjud dina lärjungar att ropa så.»
Men han svarade och sade: »Jag säger eder: Om dessa tiga, skola stenarna ropa.»
Då han nu kom närmare och fick se staden, begynte han gråta över den
och sade: »O att du i dag hade insett, också du, vad din frid tillhör!
Men nu är det fördolt för dina ögon.
Ty den tid skall komma över dig, då dina fiender skola omgiva dig med belägringsvall och innesluta dig och tränga dig på alla sidor.
Och de skola slå ned dig till jorden, tillika med dina barn, som äro i dig, och skola icke lämna kvar i dig sten på sten, därför att du icke aktade på den tid då du var sökt.»
Och han gick in i helgedomen och begynte driva ut dem som sålde därinne;
och han sade till dem: »Det är skrivet: 'Och mitt hus skall vara ett bönehus.'
Men I haven gjort det till en rövarkula.»
Och han undervisade var dag i helgedomen.
Och översteprästerna och de skriftlärde och folkets förnämste män sökte efter tillfälle att förgöra honom;
men de kunde icke finna någon utväg därtill, ty allt folket höll sig till honom och hörde honom.
Och en dag, då han undervisade folket i helgedomen och förkunnade evangelium, trädde översteprästerna och de skriftlärde, tillika med de äldste, fram
och talade till honom och sade: »Säg oss, med vad myndighet gör du detta?
Och vem är det som har rivit dig sådan myndighet?»
Han svarade och sade till dem: »Också jag vill ställa en fråga till eder; svaren mig på den.
Johannes' döpelse, var den från himmelen eller från människor?»
Då överlade de med varandra och sade: »Om vi svara: 'Från himmelen' så frågar han: 'Varför trodden I honom då icke?'
Men om vi svara: 'Från människor', då kommer allt folket att stena oss, ty de äro förvissade om att Johannes var en profet.»
De svarade alltså att de icke visste varifrån den var.
Då sade Jesus till dem: »Så säger icke heller jag eder med vad myndighet jag gör detta.»
Och han framställde för folket denna liknelse: »En man planterade en vingård och lejde ut den åt vingårdsmän och för utrikes för lång tid.
När sedan rätta tiden var inne, sände han en tjänare till vingårdsmännen, för att de åt denne skulle lämna någon del av vingårdens frukt.
Men vingårdsmännen misshandlade honom och läto honom gå tomhänt bort.
Ytterligare sände han en annan tjänare.
Också honom misshandlade och skymfade de och läto honom gå tomhänt bort.
Ytterligare sände han en tredje.
Men också denne slogo de blodig och drevo bort honom.
Då sade vingårdens herre: 'Vad skall jag göra?
Jo, jag vill sända min älskade son; för honom skola de väl ändå hava försyn.'
Men när vingårdsmannen fingo se honom, överlade de med varandra och sade: 'Denne är arvingen; låt oss dräpa honom, för att arvet må bliva vårt.'
Och de förde honom ut ur vingården och dräpte honom. »Vad skall nu vingårdens herre göra med dem?
Jo, han skall komma och förgöra de vingårdsmännen och lämna vingården åt andra.»
När de hörde detta, sade de: »Bort det!»
Då såg han på dem och sade: »Vad betyder då detta skriftens ord: 'Den sten som byggningsmännen förkastade, den har blivit en hörnsten'?
Var och en som faller på den stenen, han skall bliva krossad; men den som stenen faller på, honom skall den söndersmula.»
Och de skriftlärde och översteprästerna hade gärna velat i samma stund gripa honom, men de fruktade för folket.
Ty de förstodo att det var om dem som han hade talat i denna liknelse.
Och de vaktade på honom och sände ut några som försåtligen skulle låtsa sig vara rättsinniga män, för att dessa skulle fånga honom genom något hans ord, så att de skulle kunna överlämna honom åt överheten, i landshövdingens våld.
Dessa frågade honom och sade: »Mästare, vi veta att du talar och undervisar rätt och icke har anseende till personen, utan lär om Guds väg vad sant är.
Är det lovligt för oss att giva kejsaren skatt, eller är det icke lovligt?»
Men han märkte deras illfundighet och sade till dem:
»Låten mig se en penning.
Vems bild och överskrift bär den?»
De svarade: »Kejsarens.»
Då sade han till dem: »Given alltså kejsaren vad kejsaren tillhör, och Gud vad Gud tillhör.»
Och de förmådde icke fånga honom genom något hans ord inför folket, utan förundrade sig över hans svar och tego.
Därefter trädde några sadducéer fram och ville påstå att det icke gives någon uppståndelse.
Dessa frågade honom
och sade: »Mästare, Moses har givit oss den föreskriften, att om någon har en broder som är gift, men dör barnlös, så skall han taga sin broders hustru till akta och skaffa avkomma åt sin broder.
Nu voro här sju bröder.
Den förste tog sig en hustru, men dog barnlös.
Då tog den andre i ordningen henne
och därefter den tredje; sammalunda alla sju.
Men de dogo alla, utan att någon av dem lämnade barn efter sig.
Slutligen dog ock hustrun.
Vilken av dem skall då vid uppståndelsen få kvinnan till hustru?
De hade ju alla sju tagit henne till hustru.»
Jesus svarade dem: »Med den nuvarande tidsålderns barn är det så, att män taga sig hustrur, och hustrur givas åt män;
men de som bliva aktade värdiga att få del i den nya tidsåldern och i uppståndelsen från de döda, med dem är det så, att varken män tag sig hustrur, eller hustrur givas män.
De kunna ju ej heller mer dö ty de äro lika änglarna och äro, Guds söner, eftersom de hava blivit delaktiga av uppståndelsen.
Men att de döda uppstå, det har ock Moses, på det ställe där det talas om törnbusken, givit till känna, när han kallar Herren 'Abrahams Gud och Isaks Gud och Jakobs Gud';
Och han är en Gud icke för döda, utan för levande, ty för honom leva alla.»
Då svarade några av de skriftlärde och sade: »Mästare, du har talat rätt.»
De dristade sig nämligen icke att vidare ställa någon fråga på honom.
Men han sade till dem: »Huru kan man säga att Messias är Davids son?
David själv säger ju i Psalmernas bok: Herren sade till min herre: Sätt dig på min högra sida,
till dess jag har lagt dina fiender dig till en fotapall.'
David kallar honom alltså 'herre'; huru kan han då vara hans son?»
Och han sade till sina lärjungar, så att allt folket hörde det:
»Tagen eder till vara för de skriftlärde, som gärna gå omkring i fotsida kläder och gärna vilja bliva hälsade på torgen och gärna sitta främst i synagogorna och på de främsta platserna vid gästabuden --
detta under det att de utsuga änkors hus, medan de för syns skull hålla långa baner.
Del skola få en dess hårdare dom.»
Och när han såg upp, fick han se huru de rika lade ned sina gåvor i offerkistorna.
Därvid fick han ock se huru en fattig änka lade ned två skärvar.
Då sade han: »Sannerligen säger jag eder: Denna fattiga änka lade dit mer än alla de andra.
Ty det var av sitt överflöd som alla dessa lade ned något bland gåvorna, men hon lade dit av sitt armod allt vad hon hade i sin ägo.»
Och då några talade om helgedomen, huru den var uppförd av härliga stenar och prydd med helgedomsskänker, sade han:
»Dagar skola komma, då av allt detta som I nu sen icke skall lämnas sten på sten, utan allt skall bliva nedbrutet.»
Då frågade de honom och sade: »Mästare, när skall detta ske?
Och vad bliver tecknet till att tiden är inne, då detta kommer att ske?»
Han svarade: »Sen till, att I icke bliven förvillade.
Ty många skola komma under mitt namn och säga: 'Det är jag' och: 'Tiden är nära'.
Men följen dem icke.
Och när I fån höra krigslarm och upprorslarm, så bliven icke förfärade; ty sådant måste först komma, men därmed är icke strax änden inne.»
Därefter sade han till dem: »Folk skall resa sig upp mot folk och rike mot rike;
och det skall bliva stora jordbävningar, så ock hungersnöd och farsoter på den ena orten efter den andra, och skräcksyner skola visa sig och stora tecken på himmelen.
Men före allt detta skall man gripa eder, man skall förfölja eder och draga eder inför synagogorna och sätta eder i fängelse och föra eder fram inför konungar och landshövdingar, för mitt namns skull.
Så skolen I få tillfälle att frambära vittnesbörd.
Märken därför noga att I icke förut mån göra eder bekymmer för huru I skolen försvara eder.
Ty jag skall giva eder sådana ord och sådan vishet, att ingen av edra vedersakare skall kunna stå emot eller säga något emot.
I skolen bliva förrådda till och med av föräldrar och bröder och fränder och vänner; och somliga av eder skall man döda.
Och I skolen bliva hatade av alla för mitt namns skull.
Men icke ett hår på edra huvuden skall gå förlorat.
Genom att vara ståndaktiga skolen I vinna edra själar.
Men när I fån se Jerusalem omringas av krigshärar, då skolen I veta att dess ödeläggelse är nära.
Då må de som äro i Judeen fly bort till bergen, och de som äro inne i staden må draga ut därifrån och de som äro ute på landsbygden må icke gå ditin.
Ty detta är en hämndens tid, då allt som är skrivet skall uppfyllas.
Ve dem som äro havande, eller som giva di på den tiden!
Ty stor nöd skall då komma i landet, och en vredesdom över detta folk.
Och de skola falla för svärdsegg och bliva bortförda i fångenskap till allahanda hednafolk; och Jerusalem skall bliva förtrampat av hedningarna, till dess att hedningarnas tider äro fullbordade.
Och tecken skola ske i solen och månen och i stjärnorna, och på jorden skall ångest komma över folken, och de skola stå rådlösa vid havets och vågornas dån,
då nu människor uppgiva andan av förskräckelse och ängslan för det som skall övergå världen; ty himmelens makter skola bäva.
Och då skall man få se 'Människosonen komma i en sky', med stor makt och härlighet.
Men när detta begynner ske, då mån I resa eder upp och upplyfta edra huvuden, ty då nalkas eder förlossning.»
Och han framställde för dem en liknelse: »Sen på fikonträdet och på alla andra träd.
När I fån se att de skjuta knopp, då veten I av eder själva att sommaren redan är nära.
Likaså, när I sen detta ske, då kunnen I ock veta att Guds rike är nära.
Sannerligen säger jag eder: Detta släkte skall icke förgås, förrän allt detta sker.
Himmel och jord skola förgås, men mina ord skola aldrig förgås.
Men tagen eder till vara för att låta edra hjärtan förtyngas av omåttlighet och dryckenskap och timliga omsorger, så att den dagen kommer på eder oförtänkt;
ty såsom en snara skall den komma över hela jordens alla inbyggare.
Men vaken alltjämt, och bedjen att I mån kunna undfly allt detta som skall komma, och kunna bestå inför Människosonen.»
Och han undervisade om dagarna i helgedomen, men om aftnarna gick han ut till det berg som kallas Oljeberget och stannade där över natten.
Och allt folket kom bittida om morgonen till honom i helgedomen för att höra honom.
Det osyrade brödets högtid, som ock kallas påsk, var nu nära.
Och översteprästerna och de skriftlärde sökte efter tillfälle att röja honom ur vägen.
De fruktade nämligen för folket.
Men Satan for in i Judas, som kallades Iskariot, och som var en av de tolv.
Denne gick bort och talade med översteprästerna och befälhavarna för tempelvakten om huru han skulle överlämna honom åt dem.
Då blevo de glada och förklarade sig villiga att giva honom en summa penningar.
Och han gick in på deras anbud och sökte sedan efter lägligt tillfälle att förråda honom åt dem, utan att någon folkskockning uppstod.
Så kom nu den dag i det osyrad brödets högtid, då man skulle slakta påskalammet.
Då sände han åstad Petrus och Johannes och sade: »Gån åstad och reden till åt oss, så att vi kunna äta påskalammet.»
De frågade honom: Var vill du att vi skola reda till det?»
Han svarade dem: När I kommen in i staden, skolen I möta en man som bär en kruka vatten.
Följen honom till det hus där han går in.
Och sägen till husbonden i det huset: 'Mästaren frågar dig: Var finnes härbärget där jag skall äta påskalammet med mina lärjungar?'
Då skall han visa eder en stor sal i övre våningen, ordnad för måltid; reden till där.»
Och de gingo åstad och funno det så som han hade sagt dem; och de redde till påskalammet.
Och när stunden var inne, lade han sig till bords, och apostlarna med honom.
Och han sade till dem: »Jag har högeligen åstundat att äta detta påskalamm med eder, förrän mitt lidande begynner;
ty jag säger eder att jag icke mer skall fira denna högtid, förrän den kommer till fullbordan i Guds rike.»
Och han lät giva sig en kalk och tackade Gud och sade: »Tagen detta och delen eder emellan;
ty jag säger eder att jag härefter icke, förrän Guds rike kommer, skall dricka av det som kommer från vinträd.»
Sedan tog han ett bröd och tackade Gud och bröt det och gav åt dem och sade: »Detta är min lekamen, som varder utgiven för eder.
Gören detta till min åminnelse.»
Sammalunda tog han ock kalken, efter måltiden, och sade: »Denna kalk är det nya förbundet, i mitt blod, som varder utgjutet för eder.
Men se, den som förråder mig, hans hand är med mig på bordet.
Ty Människosonen skall gå bort, såsom förut är bestämt; men ve den människa genom vilken han bliver förrådd!»
Och de begynte tala med varandra om vilken av dem det väl kunde vara som skulle göra detta.
En tvist uppstod ock mellan dem om vilken av dem som skulle räknas för den störste.
Då sade han till dem: »Konungarna uppträda mot sina folk såsom härskare, och de som hava myndighet över folken låta kalla sig 'nådige herrar'.
Men så är det icke med eder; utan den som är störst bland eder, han vare såsom den yngste, och den som är den förnämste, han vare såsom en tjänare.
Ty vilken är större: den som ligger till bords eller den som tjänar?
Är det icke den som ligger till bords?
Och likväl är jag här ibland eder såsom en tjänare. --
Men I ären de som hava förblivit hos mig i mina prövningar;
och såsom min Fader har överlåtit konungslig makt åt mig, så överlåter jag likadan makt åt eder,
så att I skolen få äta och dricka vid mitt bord i mitt rike och sitta på troner såsom domare över Israels tolv släkter.
Simon, Simon!
Se, Satan har begärt att få eder i sitt våld, för att kunna sålla eder såsom vete;
men jag har bett för dig, att din tro icke må bliva om intet.
Och när du en gång har omvänt dig, så styrk dina bröder.»
Då sade han till honom: »Herre, jag är redo att med dig både gå i fängelse och gå i döden.»
Men han svarade: »Jag säger dig, Petrus: I dag skall icke hanen gala, förrän du tre gånger har förnekat mig och sagt att du icke känner mig.»
Ytterligare sade han till dem: »När jag sände eder åstad utan penningpung, utan ränsel, utan skor, icke fattades eder då något?»
De svarade: »Intet.»
Då sade han till dem: »Nu åter må den som har en penningpung taga den med sig, och den som har en ränsel, han göre sammalunda; och den som icke har något svärd, han sälje sin mantel och köpe sig ett sådant.
Ty jag säger eder att på mig måste fullbordas detta skriftens ord: 'Han blev räknad bland ogärningsmän'.
Ja, det som är förutsagt om mig, det går nu i fullbordan»
Då sade de: »Herre, se här äro två svärd.»
Han svarade dem: »Det är nog.»
Och han gick ut och begav sig till Oljeberget, såsom hans sed var; och hans lärjungar följde honom.
Men när han hade kommit till platsen, sade han till dem: »Bedjen att I icke mån komma i frestelse.»
Sedan gick han bort ifrån dem, vid pass ett stenkast, och föll ned på sina knän och bad
och sade: »Fader, om det är din vilja, så tag denna kalk ifrån mig.
Dock, ske icke min vilja, utan din.»
Då visade sig för honom en ängel från himmelen, som styrkte honom.
Men han hade kommit i svår ångest och bad allt ivrigare, och hans svett blev såsom blodsdroppar, som föllo ned på jorden.
När han sedan stod upp från bönen och kom tillbaka till lärjungarna, fann han dem insomnade av bedrövelse.
Då sade han till dem: »Varför soven I?
Stån upp, och bedjen att I icke mån komma i frestelse.»
Och se, medan han ännu talade, kom en folkskara; och en av de tolv, den som hette Judas, gick framför dem.
Och han trädde fram till Jesus för att kyssa honom.
Men Jesus sade till honom: »Judas, förråder du Människosonen med en kyss?»
Då nu de som voro med Jesus sågo vad som var på färde, frågade de: »Herre, skola vi hugga till med svärd?»
Och en av dem högg till översteprästens tjänare och högg så av honom högra örat.
Då svarade Jesus och sade: »Låten det gå så långt.»
Och han rörde vid hans öra och helade honom.
Sedan sade Jesus till dem som hade kommit emot honom, till översteprästerna och befälhavarna för tempelvakten och de äldste: »Såsom mot en rövare haven I gått ut med svärd och stavar.
Fastän jag var dag har varit med eder i helgedomen, haven I icke sträckt ut edra händer emot mig men detta är eder stund, och nu råder mörkrets makt.»
Så grepo de honom och förde honom åstad in i översteprästens hus.
Och Petrus följde efter på avstånd.
Och de tände upp en eld mitt på gården och satte sig där tillsammans, och Petrus satte sig ibland dem.
Men en tjänstekvinna, som fick se honom, där han satt vid elden fäste ögonen på honom och sade: »Också denne var med honom.
Men han nekade och sade: »Kvinna, jag känner honom icke.»
Kort därefter fick en annan, en av mannen, se honom och sade: »Också du är en av dem.»
Men Petrus svarade: »Nej, det är jag icke.»
Vid pass en timme därefter kom en annan som bedyrade och sade: »Förvisso var också denne med honom; han är ju ock en galilé.»
Då svarade Petrus: »Jag förstår icke vad du menar.»
Och i detsamma, medan han ännu talade, gol hanen.
Då vände Herren sig om och såg på Petrus; och Petrus kom då ihåg Herrens ord, huru han hade sagt till honom: »Förrän hanen i dag har galit, skall du tre gånger förneka mig.»
Och han gick ut och grät bitterligen.
Och de män som höllo Jesus fången begabbade honom och misshandlade honom.
De höljde över honom och frågade honom och sade: »Profetera: vem var det som slog dig?»
Många andra smädliga ord talade de ock mot honom.
Men när det blev dag, församlade sig folkets äldste, överstepräster och skriftlärde, och läto föra honom inför sitt Stora råd
och sade: »Är du Messias, så säg oss det.»
Men han svarade dem: »Om jag säger eder det, så tron I det icke.
Och om jag frågar, så svaren I icke.
Men härefter skall Människosonen sitta på den gudomliga Maktens högra sida.»
Då sade de alla: »Så är du då Guds Son?»
Han svarade dem: »I sägen det själva, att jag är det.»
Då sade de: »Vad behöva vi mer något vittnesbörd?
Vi hava ju själva nu hört det av hans egen mun.»
Och de stodo upp, hela hopen, och förde honom till Pilatus.
Där begynte de anklaga honom och sade: »Vi hava funnit att denne man förleder vårt folk och vill förhindra att man giver kejsaren skatt, och att han säger sig vara Messias, en konung.»
Då frågade Pilatus honom och sade: Är du judarnas konung?»
Han svarade honom och sade: »Du säger det själv.»
Men Pilatus sade till översteprästerna och till folket: »Jag finner intet brottsligt hos denne man.»
Då blevo de ännu ivrigare och sade: »Han uppviglar med sin lära folket i hela Judeen, allt ifrån Galileen och ända hit.»
När Pilatus hörde detta, frågade han om mannen var från Galileen.
Och då han fick veta att han var från det land som lydde under Herodes' välde, sände han honom bort till Herodes, som under dessa dalar också var i Jerusalem.
När Herodes fick se Jesus, blev han mycket glad, ty han hade sedan lång tid velat se honom; han hade nämligen hört talas om honom, och han hoppades nu att få se honom göra något tecken.
Men fastän han ställde ganska många frågor på Jesus, svarade denne honom intet.
Och översteprästerna och de skriftlärde stodo där och anklagade honom häftigt.
Men Herodes och hans krigsfolk bemötte honom med förakt och begabbade honom; och sedan de hade satt på honom en lysande klädnad, sände de honom tillbaka till Pilatus.
Och Herodes och Pilatus blevo den dagen vänner med varandra; Förut hade nämligen dem emellan rått ovänskap.
Sedan kallade Pilatus tillhopa översteprästerna och rådsherrarna och folket
och sade till dem: »I haven fört till mig denne man och sagt att han förleder folket; och jag har nu i eder närvaro anställt rannsakning med honom, men icke funnit honom skyldig till något av det som I anklagen honom för.
Och ej heller Herodes har funnit honom skyldig; han har ju sänt honom tillbaka till oss.
I sen alltså att denne icke har gjort något som förtjänar döden.
Därför vill jag giva honom lös, medan jag har tuktat honom.»
Då skriade hela hopen och sade: »Hav bort denne, och giv oss Barabbas lös.»
(Denne man hade blivit kastad i fängelse på grund av ett upplopp, som hade ägt rum i staden, och för ett dråps skull.)
Åter talade Pilatus till dem, ty han önskade att kunna giva Jesus lös.
Men de ropade emot honom: »Korsfäst, korsfäst honom!»
Då talade han till dem för tredje gången och frågade: »Vad ont har denne då gjort?
Jag har icke funnit honom skyldig till något som förtjänar döden Därför vill jag giva honom lös, sedan jag har tuktat honom.»
Men de lågo över honom med höga rop och begärde att han skulle låta korsfästa honom; och deras rop blevo honom övermäktiga.
Då dömde Pilatus att så skulle ske, som de begärde.
Och han lösgav den man de begärde, den som hade blivit kastad i fängelse för upplopp och dråp; men Jesus utlämnade han, för att med honom skulle ske efter deras vilja.
När de sedan förde bort honom, fingo de fatt en man, Simon från Cyrene, som kom utifrån marken; på honom lade de korset, för att han skulle bära det efter Jesus.
Men en stor hop folk följde med honom, bland dem också kvinnor som jämrade sig och gräto över honom.
Då vände Jesus sig om till dem och sade: »I Jerusalems döttrar, gråten icke över mig, utan gråten över eder själva och över edra barn.
Ty se, den tid skall komma, då man skall säga: 'Saliga äro de ofruktsamma, de moderliv som icke hava fött barn, och de bröst som icke hava givit di.'
Då skall man begynna säga till: bergen: 'Fallen över oss', och till höjderna: 'Skylen oss.'
Ty om han gör så med det friska trädet, vad skall icke då ske med det torra!»
Jämväl två andra, två ogärningsmän, fördes ut för att avlivas tillika med honom.
Och när de hade kommit till den plats som kallades »Huvudskallen» korsfäste de honom där, så ock ogärningsmännen, den ene på högra sidan och den andre på vänstra.
Men Jesus sade. »Fader, förlåt dem; ty de veta icke vad de göra.
Och de delade hans kläder mellan sig och kastade lott om dem. --
Men folket stod och såg därpå.
Och jämväl rådsherrarna drevo gäck med honom och sade: »Andra har han hjälpt; nu må han hjälpa sig själv, om han är Guds Smorde, den utvalde.»
Också krigsmännen gingo fram och begabbade honom och räckte honom ättikvin
och sade: »Är du judarnas konung, så hjälp dig själv.»
Men över honom hade man ock satt upp en överskrift: »Denne är judarnas konung.»
Och en av de ogärningsmän som voro där upphängda smädade honom och sade: »Du är ju Messias; hjälp då dig själv och oss.»
Då tillrättavisade honom den andre och svarade och sade: »Fruktar icke heller du Gud, du som är under samma dom?
Oss vederfares detta med all rätt, ty vi lida vad våra gärningar äro värda, men denne man har intet ont gjort.»
Sedan sade han: »Jesus, tänk på mig, när du kommer i ditt rike.»
Han svarade honom: »Sannerligen säger jag dig: I dag skall du vara med mig i paradiset.»
Det var nu omkring sjätte timmen; då kom över hela landet ett mörker, som varade ända till nionde timmen,
i det att solen miste sitt sken.
Och förlåten i templet rämnade mitt itu.
Och Jesus ropade med hög röst och sade: »Fader, i dina händer befaller jag min ande.»
Och när han hade sagt detta, gav han upp andan.
Men när hövitsmannen såg vad som skedde, prisade han Gud och sade: »Så var då denne verkligen en rättfärdig man!»
Och när allt folket, de som hade kommit tillsammans för att se härpå, sågo vad som skedde, slogo de sig för bröstet och vände hem igen.
Men alla hans vänner stodo på avstånd och sågo detta, bland dem också några kvinnor, de som hade följt med honom från Galileen.
Nu var där en rådsherre, vi namn Josef, en god och rättfärdig man,
som icke hade samtyckt till deras rådslag och gärning.
Han var från Arimatea, en stad i Judeen; och han väntade på Guds rike.
Denne gick till Pilatus och utbad sig att få Jesu kropp.
Och han tog ned den och svepte den i en linneduk.
Sedan lade han den i en grav som var uthuggen i klippan, och där ännu ingen hade varit lagd.
Det var då tillredelsedag, och sabbatsdagen begynte ingå.
Och de kvinnor, som med honom hade kommit från Galileen, följde efter och sågo graven och sågo huru hans kropp lades ned däri.
Sedan vände de hem igen och redde till välluktande kryddor och smörjelse; men på sabbaten voro de stilla, efter lagens bud.
Men på första veckodagen kommo de, tidigt i själva dagbräckningen, till graven med de välluktande kryddor som de hade tillrett.
Och de funno stenen vara bortvältrad från graven.
Då gingo de ditin, men funno icke Herren Jesu kropp.
När de nu icke visste vad de skulle tänka härom, se, då stodo två man framför dem i skinande kläder.
Och de blevo förskräckta och böjde sina ansikten ned mot jorden.
Då sade mannen till dem »Varför söken I den levande bland de döda?
Han är icke har, han är uppstånden.
Kommen ihåg vad han talade till eder, medan han ännu var i Galileen, huru han sade:
'Människosonen måste bliva överlämnad i syndiga människors händer och bliva korsfäst; men på tredje dagen skall han uppstå igen.'»
Då kommo de ihåg hans ord.
Och de vände tillbaka från graven och omtalade allt detta för de elva och för alla de andra. --
Kvinnorna voro Maria från Magdala och Johanna och den Maria som var Jakobs moder.
Och jämväl de andra kvinnorna instämde med dem och sade detsamma till apostlarna.
Deras ord syntes dock för dessa vara löst tal, och de trodde dem icke.
Men Petrus stod upp och skyndade till graven; och när han lutade sig ditin såg han där allenast linnebindlarna.
Sedan gick han hem till sitt, uppfylld av förundran över det som hade skett.
Men två av dem voro samma dag stadda på vandring till en by som hette Emmaus, och som låg sextio stadiers väg från Jerusalem.
Och de samtalade med varandra om allt detta som hade skett.
Medan de nu samtalade och överlade med varandra, nalkades Jesus själv och gick med dem.
Men deras ögon voro tillslutna, så att de icke kände igen honom.
Och han sade till dem: »Vad är det I talen om med varandra, medan I gån här?»
Då stannade de och sågo bedrövade ut.
Och den ene, som hette Kleopas, svarade och sade till honom: »Du är väl en främling i Jerusalem, den ende som icke har hört vad där har skett i dessa dagar?»
Han frågade dem: »Vad då?»
De svarade honom: »Det som har skett med Jesus från Nasaret, vilken var en profet, mäktig i gärningar och ord inför Gud och allt folket:
huru nämligen våra överstepräster och rådsherrar hava utlämnat honom till att dömas till döden och hava korsfäst honom.
Men vi hoppades att han var den som skulle förlossa Israel.
Och likväl, till allt detta kommer att det redan är tredje dagen sedan detta skedde.
Men nu hava därjämte några av våra kvinnor gjort oss häpna; ty sedan de bittida på morgonen hade varit vid graven
och icke funnit hans kropp, kommo de igen och sade att de till och med hade sett en änglasyn, och änglarna hade sagt att han levde.
Och när några av dem som voro. med oss gingo bort till graven, funno de det vara så som kvinnorna hade sagt, men honom själv sågo de icke.»
Då sade han till dem: »O, huru oförståndiga ären I icke och tröghjärtade till att tro på allt vad profeterna hava talat!
Måste icke Messias lida detta, för I att så ingå i sin härlighet?»
Och han begynte att genomgå Moses och alla profeterna och uttydde för dem vad som i alla skrifterna var sagt om honom.
När de nu nalkades byn dit de voro på väg, ställde han sig som om han ville gå vidare.
Men de nödgade honom och sade: »Bliv kvar hos oss, ty det lider mot aftonen, och dagen nalkas redan sitt slut.»
Då gick han ditin och stannade kvar hos dem.
Och när han nu låg till bords med dem, tog han brödet och välsignade och bröt det och räckte åt dem.
Därvid öppnades deras ögon, så att de kände igen honom.
Men då försvann han ur deras åsyn.
Och de sade till varandra: »Voro icke våra hjärtan brinnande i oss, när han talade med oss på vägen och uttydde skrifterna för oss?»
Och i samma stund stodo de upp och vände tillbaka till Jerusalem; och de funno där de elva församlade, så ock de andra som hade slutit sig till dem.
Och dessa sade: »Herren är verkligen uppstånden, och han har visat sig för Simon.»
Då förtäljde de själva vad som hade skett på vägen, och huru han hade blivit igenkänd av dem, när han bröt brödet.
Medan de nu talade härom, stod han själv mitt ibland dem och sade till dem: »Frid vare med eder.
Då blevo de förfärade och uppfylldes av fruktan och trodde att det var en ande de sågo.
Men han sade till dem: »Varför ären I så förskräckta, och varför uppstiga tvivel i edra hjärtan?
Sen här mina händer och mina fötter, och sen att det är jag själv; ja, tagen på mig och sen.
En ande har ju icke kött och ben, såsom I sen mig hava.»
Och när han hade sagt detta, visade han dem sina händer och sina fötter.
Men då de ännu icke trodde, för glädjes skull, utan allenast förundrade sig, sade han till dem: »Haven I här något att äta?»
Då räckte de honom ett stycke stekt fisk och något av en honungskaka;
och han tog det och åt därav i deras åsyn.
Och han sade till dem: »Det är såsom jag sade till eder, medan jag ännu var bland eder, att allt måste fullbordas, som är skrivet om mig i Moses' lag och hos profeterna och i psalmerna.»
Därefter öppnade han deras sinnen, så att de förstodo skrifterna.
Och han sade till dem: »Det är så skrivet, att Messias skulle lida och på tredje dagen uppstå från de döda,
och att bättring till syndernas förlåtelse i hans namn skulle predikas bland alla folk, och först i Jerusalem.
I kunnen vittna härom.
Och se, jag vill sända till eder vad min Fader har utlovat.
Men I skolen stanna kvar här i staden, till dess I från höjden bliven beklädda med kraft.»
Sedan förde han dem ut till Betania; och där lyfte han upp sina händer och välsignade dem.
Och medan han välsignade dem, försvann han ifrån dem och blev upptagen till himmelen.
Då tillbådo de honom och vände sedan tillbaka till Jerusalem, uppfyllda av stor glädje.
Och de voro sedan alltid i helgedomen och lovade Gud.
I begynnelsen var Ordet, och Ordet var hos Gud, och Ordet var Gud.
Detta var i begynnelsen hos Gud.
Genom det har allt blivit till, och utan det har intet blivit till, som är till.
I det var liv, och livet var människornas ljus.
Och ljuset lyser i mörkret, och mörkret har icke fått makt därmed.
En man uppträdde, sänd av Gud; hans namn var Johannes.
Han kom såsom ett vittne, för att vittna om ljuset, på det att alla skulle komma till tro genom honom.
Icke var han ljuset, men han skulle vittna om ljuset.
Det sanna ljuset, det som lyser över alla människor, skulle nu komma i världen.
I världen var han, och genom honom hade världen blivit till, men världen ville icke veta av honom.
Han kom till sitt eget, och hans egna togo icke emot honom.
Men åt alla dem som togo emot honom gav han makt att bliva Guds barn, åt dem som tro på hans namn;
och de hava blivit födda, icke av blod, ej heller av köttslig vilja, ej heller av någon mans vilja, utan av Gud.
Och Ordet vart kött och tog sin boning ibland oss, och vi sågo hans härlighet, vi sågo likasom en enfödd Sons härlighet från sin Fader, och han var full av nåd och sanning.
Johannes vittnar om honom, han ropar och säger: »Det var om denne jag sade: 'Den som kommer efter mig, han är före mig; ty han var förr än jag.'»
Av hans fullhet hava vi ju alla fått, ja, nåd utöver nåd;
ty genom Moses blev lagen given, men nåden och sanningen hava kommit genom Jesus Kristus.
Ingen har någonsin sett Gud; den enfödde Sonen, som är i Faderns sköte, han har kungjort vad Gud är.
Och detta är vad Johannes vittnade, när judarna hade sänt till honom präster och leviter från Jerusalem för att fråga honom vem han var.
Han svarade öppet och förnekade icke; han sade öppet: »Jag är icke Messias.»
Åter frågade de honom: »Vad är du då?
Är du Elias?»
Han svarade: »Det är jag icke.» -- »Är du Profeten?»
Han svarade: »Nej.»
Då sade de till honom: »Vem är du då?
Säg oss det, så att vi kunna giva dem svar, som hava sänt oss.
Vad säger du om dig själv?»
Han svarade: »Jag är rösten av en som ropar i öknen: 'Jämnen vägen för Herren', såsom profeten Esaias sade.»
Och männen voro utsända ifrån fariséerna.
Och de frågade honom och sade till honom: »Varför döper du då, om du icke är Messias, ej heller Elias, ej heller Profeten?»
Johannes svarade dem och sade: »Jag döper i vatten; men mitt ibland eder står en som I icke kännen:
han som kommer efter mig, vilkens skorem jag icke är värdig att upplösa.»
Detta skedde i Betania, på andra sidan Jordan, där Johannes döpte.
Dagen därefter såg han Jesus nalkas; då sade han: »Se, Guds Lamm, som borttager världens synd!
Om denne var det som jag sade: 'Efter mig kommer en man som är före mig; ty han var förr än jag.'
Och jag kände honom icke; men för att han skall bliva uppenbar för Israel, därför är jag kommen och döper i vatten.»
Och Johannes vittnade och sade: »Jag såg Anden såsom en duva sänka sig ned från himmelen; och han förblev över honom.
Och jag kände honom icke; men den som sände mig till att döpa i vatten, han sade till mig: 'Den över vilken du får se Anden sänka sig ned och förbliva, han är den som döper i helig ande.'
Och jag har sett det, och jag har vittnat att denne är Guds Son.»
Dagen därefter stod Johannes åter där med två av sina lärjungar.
När då Jesus kom gående, såg Johannes på honom och sade: »Se, Guds Lamm!»
Och de två lärjungarna hörde hans ord och följde Jesus.
Då vände sig Jesus om, och när han såg att de följde honom, frågade han dem: »Vad viljen I?»
De svarade honom: »Rabbi» (det betyder mästare) »var bor du?»
Han sade till dem: »Kommen och sen.»
Då gingo de med honom och sågo var han bodde; och de stannade den dagen hos honom. -- Detta skedde vid den tionde timmen.
En av de två som hade hört var Johannes sade, och som hade följt Jesus, var Andreas, Simon Petrus' broder.
Denne träffade först sin broder Simon och sade till honom: »Vi hava funnit Messias» (det betyder detsamma som Kristus).
Och han förde honom till Jesus.
Då såg Jesus på honom och sade: »Du är Simon, Johannes' son; du skall heta Cefas» (det betyder detsamma som Petrus).
Dagen därefter ville Jesus gå därifrån till Galileen, och han träffade då Filippus.
Och Jesus sade till honom: »Följ mig.»
Och Filippus var från Betsaida, Andreas' och Petrus' stad.
Filippus träffade Natanael och sade till honom: »Den som Moses har skrivit om i lagen och som profeterna hava skrivit om, honom hava vi funnit, Jesus, Josefs son, från Nasaret.»
Natanael sade till honom: »Kan något gott komma från Nasaret?»
Filippus svarade honom: »Kom och se.»
När nu Jesus såg Natanael nalkas, sade han om honom: »Se, denne är en rätt israelit, i vilken icke finnes något svek.»
Natanael frågade honom: »Huru kunna du känna mig?»
Jesus svarade och sade till honom: »Förrän Filippus kallade dig, såg jag dig, där du var under fikonträdet.»
Natanael svarade honom: »Rabbi, du är Guds Son, du är Israels konung.»
Jesus svarade och sade till honom: »Eftersom jag sade dig att jag såg dig under fikonträdet, tror du?
Större ting än vad detta är skall du få se.»
Därefter sade han till honom: »Sannerligen, sannerligen säger jag eder: I skolen få se himmelen öppen och Guds änglar fara upp och fara ned över Människosonen.»
På tredje dagen var ett bröllop i Kana i Galileen, och Jesu moder var där.
Också Jesus och hans lärjungar blevo bjudna till bröllopet.
Och vinet begynte taga slut.
Då sade Jesu moder till honom: »De hava intet vin.»
Jesus svarade henne: »Låt mig vara, moder; min stund är ännu icke kommen.»
Hans moder sade då till tjänarna: »Vadhelst han säger till eder, det skolen I göra.»
Nu stodo där sex stenkrukor, sådana som judarna hade för sina reningar; de rymde två eller tre bat-mått var.
Jesus sade till dem: »Fyllen krukorna med vatten.»
Och de fyllde dem ända till brädden.
Sedan sade han till dem: »Ösen nu upp och bären till övertjänaren.»
Och de gjorde så.
Och övertjänaren smakade på vattnet, som nu hade blivit vin; och han visste icke varifrån det hade kommit, vilket däremot tjänarna visste, de som hade öst upp vattnet.
Då kallade övertjänaren på brudgummen.
och sade till honom: »Man brukar eljest alltid sätta fram det goda vinet, och sedan, när gästerna hava fått för mycket, det som är sämre.
Du har gömt det goda vinet ända tills nu.»
Detta var det första tecknet som Jesus gjorde.
Han gjorde det i Kana i Galileen och uppenbarade så sin härlighet; och hans lärjungar trodde på honom.
Därefter begav han sig ned till Kapernaum med sin moder och sina bröder och sina lärjungar; och där stannade de några få dagar.
Judarnas påsk var nu nära, och Jesus begav sig då upp till Jerusalem.
Och när han fick i helgedomen se huru där sutto män som sålde fäkreatur och får och duvor, och huru växlare sutto där.
Då gjorde han sig ett gissel av tåg och drev dem alla ut ur helgedomen, med får och fäkreatur, och slog ut växlarnas penningar och stötte omkull deras bord.
Och till duvomånglarna sade han: »Tagen bort detta härifrån; gören icke min Faders hus till ett marknadshus.»
Hans lärjungar kommo då ihåg att det var skrivet: »Nitälskan för ditt hus skall förtära mig.»
Då togo judarna till orda och sade till honom: »Vad för tecken låter du oss se, eftersom du gör på detta sätt?»
Jesus svarade och sade till dem: »Bryten ned detta tempel, så skall jag inom tre dagar låta det uppstå igen.»
Då sade judarna: »I fyrtiosex år har man byggt på detta tempel, och du skulle låta det uppstå igen inom tre dagar?»
Men det var om sin kropps tempel han talade.
Sedan, när han hade uppstått från de döda, kommo hans lärjungar ihåg att han hade sagt detta; och de trodde då skriften och det ord som Jesus hade sagt.
Medan han nu var i Jerusalem, under påsken, vid högtiden, kommo många till tro på hans namn, när de sågo de tecken som han gjorde.
Men själv betrodde sig Jesus icke åt dem, eftersom han kände alla
och icke behövde någon annans vittnesbörd om människorna; ty av sig själv visste han vad i människan var.
Men bland fariséerna var en man som hette Nikodemus, en av judarnas rådsherrar.
Denne kom till Jesus om natten och sade till honom: »Rabbi, vi veta att det är från Gud du har kommit såsom lärare; ty ingen kan göra sådana tecken som du gör, om icke Gud är med honom.»
Jesus svarade och sade till honom: »Sannerligen, sannerligen säger jag dig: Om en människa icke bliver född på nytt, så kan hon icke få se Guds rike.»
Nikodemus sade till honom: »Huru kan en människa födas, när hon är gammal?
Icke kan hon väl åter gå in i sin moders liv och födas?»
Jesus svarade: »Sannerligen, sannerligen säger jag dig: Om en människa icke bliver född av vatten och ande, så kan hon icke komma in i Guds rike.
Det som är fött av kött, det är kött; och det som är fött av Anden, det är ande.
Förundra dig icke över att jag sade dig att I måsten födas på nytt.
Vinden blåser vart den vill, och du hör dess sus, men du vet icke varifrån den kommer, eller vart den far; så är det med var och en som är född av Anden.»
Nikodemus svarade och sade till honom: »Huru kan detta ske?»
Jesus svarade och sade till honom: »Är du Israels lärare och förstår icke detta?
Sannerligen, sannerligen säger jag dig: Vad vi veta, det tala vi, och vad vi hava sett, det vittna vi om, men vårt vittnesbörd tagen I icke emot.
Tron i icke, när jag talar till eder om jordiska ting, huru skolen I då kunna tro, när jag talar till eder om himmelska ting?
Och likväl har ingen stigit upp till himmelen, utom den som steg ned från himmelen, Människosonen, som var i himmelen.
Och såsom Moses upphöjde ormen i öknen, så måste Människosonen bliva upphöjd,
så att var och en som tror skall i honom hava evigt liv.
Ty så älskade Gud världen, att han utgav sin enfödde Son, på det att var och en som tror på honom skall icke förgås, utan hava evigt liv.
Ty icke sände Gud sin Son i världen för att döma världen, utan för att världen skulle bliva frälst genom honom.
Den som tror på honom, han bliver icke dömd, men den som icke tror, han är redan dömd, eftersom han icke tror på Guds enfödde Sons namn.
Och detta är domen, att när ljuset hade kommit i världen, människorna dock älskade mörkret mer än ljuset, eftersom deras gärningar voro onda,
Ty var och en som gör vad ont är, han hatar ljuset och kommer icke till ljuset, på det att hans gärningar icke skola bliva blottade.
Men den som gör sanningen, han kommer till ljuset, för att det skall bliva uppenbart att hans gärningar äro gjorda i Gud.»
Därefter begav sig Jesus med sina lärjungar till den judiska landsbygden, och där vistades han med dem och döpte.
Men också Johannes döpte, i Enon, nära Salim, ty där fanns mycket vatten; och folket kom dit och lät döpa sig.
Johannes hade nämligen ännu icke blivit kastad i fängelse.
Då uppstod mellan Johannes' lärjungar och en jude en tvist om reningen.
Och de kommo till Johannes och sade till honom: »Rabbi, se, den som var hos dig på andra sidan Jordan, den som du har vittnat om, han döper, och alla komma till honom.»
Johannes svarade och sade: »En människa kan intet taga, om det icke bliver henne givet från himmelen.»
I kunnen själva giva mig det vittnesbördet att jag sade: 'Icke är jag Messias; jag är allenast sänd framför honom.'
Brudgum är den som har bruden; men brudgummens vän, som står där och hör honom, han gläder sig storligen åt brudgummens röst.
Den glädjen är mig nu given i fullt mått.
Det är såsom sig bör att han växer till, och att jag förminskas. --
Den som kommer ovanifrån, han är över alla; den som är från jorden, han är av jorden, och av jorden talar han.
Ja, den som kommer från himmelen, han är över alla,
och vad han har sett och hört, det vittnar han om; och likväl tager ingen emot hans vittnesbörd.
Men om någon tager emot hans vittnesbörd, så bekräftar han därmed att Gud är sannfärdig.
Ty den som Gud har sänt, han talar Guds ord; Gud giver nämligen icke Anden efter mått.
Fadern älskar Sonen, och allt har han givit i hans hand.
Den som tror på Sonen, han har evigt liv; men den som icke hörsammar Sonen, han skall icke få se livet, utan Guds vrede förbliver över honom.»
Men Herren fick nu veta att fariséerna hade hört hurusom Jesus vann flera lärjungar och döpte flera än Johannes;
dock var det icke Jesus själv som döpte, utan hans lärjungar.
Då lämnade han Judeen och begav sig åter till Galileen.
Därvid måste han taga vägen genom Samarien.
Så kom han till en stad i Samarien som hette Sykar, nära det jordstycke som Jakob gav åt sin son Josef.
Och där var Jakobs brunn.
Eftersom nu Jesus var trött av vandringen, satte han sig strax ned vid brunnen.
Det var vid den sjätte timmen.
Då kom en samaritisk kvinna för att hämta vatten.
Jesus sade till henne: »Giv mig att dricka.»
Hans lärjungar hade nämligen gått in i staden för att köpa mat.
Då sade den samaritiska kvinnan till honom: »Huru kan du, som är jude, bedja mig, som är en samaritisk kvinna, om något att dricka?»
Judarna hava nämligen ingen umgängelse med samariterna.
Jesus svarade och sade till henne: »Förstode du Guds gåva, och vem den är som säger till dig: 'Giv mig att dricka', så skulle i stället du hava bett honom, och han skulle då hava givit dig levande vatten.»
Kvinnan sade till honom: »Herre, du har ju intet att hämta upp vatten med, och brunnen är djup.
Varifrån får du då det friska vattnet?»
Icke är du väl förmer än vår fader Jakob, som gav oss brunnen och själv med sina barn och sin boskap drack ur den?»
Jesus svarade och sade till henne: »Var och en som dricker av detta vatten, han bliver törstig igen;
men den som dricker av det vatten som jag giver honom, han skall aldrig någonsin törsta, utan det vatten jag giver honom skall bliva i honom en källa vars vatten springer upp med evigt liv.»
Kvinnan sade till honom: »Herre, giv mig det vattnet, så att jag icke mer behöver törsta och komma hit för att hämta vatten.»
Han sade till henne: »Gå och hämta din man, och kom sedan tillbaka.»
Kvinnan svarade och sade: »Jag har ingen man.»
Jesus sade till henne: »Du har rätt i vad du säger, att du icke har någon man.»
Ty fem män har du haft, och den du nu har är icke din man; däri sade du sant.
Då sade kvinnan till honom: »Herre, jag ser att du är en profet.
Våra fäder hava tillbett på detta berg, men I sägen att i Jerusalem den plats finnes, där man bör tillbedja.»
Jesus sade till henne: »Tro mig, kvinna: den tid kommer, då det varken är på detta berg eller i Jerusalem som I skolen tillbedja Fadern.
I tillbedjen vad I icke kännen, vi tillbedja vad vi känna -- ty frälsningen kommer från judarna --
men den tid skall komma, ja, den är redan inne, då sanna tillbedjare skola tillbedja Fadern i ande och sanning; ty sådana tillbedjare vill Fadern hava.
Gud är ande, och de som tillbedja måste tillbedja i ande och sanning.»
Kvinnan sade till honom: »Jag vet att Messias skall komma, han som ock kallas Kristus; när han kommer, skall han förkunna oss allt.»
Jesus svarade henne: »Jag, som talar med dig, är den du nu nämnde.»
I detsamma kommo hans lärjungar; och de förundrade sig över att han talade med en kvinna.
Dock frågade ingen vad han ville henne, eller varför han talade med henne.
Men kvinnan lät sin kruka stå och gick in i staden och sade till folket:
»Kommen och sen en man som har sagt mig allt vad jag har gjort.
Månne icke han är Messias?»
Då gingo de ut ur staden och kommo till honom.
Under tiden bådo lärjungarna honom och sade: »Rabbi, tag och ät.»
Men han svarade dem: »Jag har mat att äta som I icke veten om.»
Då sade lärjungarna till varandra: »Kan väl någon hava burit mat till honom?»
Jesus sade till dem: »Min mat är att göra dens vilja, som har sänt mig, och att fullborda hans verk.»
I sägen ju att det ännu är fyra månader innan skördetiden kommer.
Men se, jag säger eder: Lyften upp edra ögon, och sen på fälten, huru de hava vitnat till skörd.
Redan nu får den som skördar uppbära sin lön och samla in frukt till evigt liv; så kunna den som sår och den som skördar tillsammans glädja sig.
Ty här sannas det ordet, att en är den som sår och en annan den som skördar.
Jag har sänt eder att skörda, där I icke haven arbetat.
Andra hava arbetat, och I haven fått gå in i deras arbete.»
Och många samariter från den staden kommo till tro på honom för kvinnans ords skull, då hon vittnade att han hade sagt henne allt vad hon hade gjort.
När sedan samariterna kommo till honom, både de honom att stanna kvar hos dem.
Så stannade han där i två dagar.
Och långt flera kommo då till tro för hans egna ords skull.
Och de sade till kvinnan: »Nu är det icke mer för dina ords skull som vi tro, ty vi hava nu själva hört honom, och vi veta nu att han i sanning är världens Frälsare.»
Men efter de två dagarna gick han därifrån till Galileen.
Ty Jesus vittnade själv att en profet icke är aktad i sitt eget fädernesland.
När han nu kom till Galileen, togo galiléerna vänligt emot honom, eftersom de hade sett allt vad han hade gjort i Jerusalem vid högtiden.
Också de hade nämligen varit där vid högtiden.
Så kom han åter till Kana i Galileen, där han hade gjort vattnet till vin.
I Kapernaum fanns då en man i konungens tjänst, vilkens son låg sjuk.
När han nu hörde att Jesus hade kommit från Judeen till Galileen, begav han sig åstad till honom och bad att han skulle komma ned och bota hans son; ty denne låg för döden.
Då sade Jesus till honom: »Om I icke sen tecken och under, så tron I icke.»
Mannen sade till honom: »Herre, kom ned, förrän mitt barn dör.»
Jesus svarade honom: »Gå, din son får leva.»
Då trodde mannen det ord som Jesus sade till honom, och gick.
Och medan han ännu var på vägen hem, mötte honom hans tjänare och sade: »Din son kommer att leva.»
Då frågade han dem vid vilken timme det hade blivit bättre med honom.
De svarade honom: »I går vid den sjunde timmen lämnade febern honom.»
Då märkte fadern att det hade skett just den timme då Jesus sade till honom: »Din son får leva.»
Och han kom till tro, så ock hela hans hus.
Detta var nu åter ett tecken, det andra i ordningen som Jesus gjorde, sedan han hade kommit från Judeen till Galileen.
Därefter inföll en av judarnas högtider, och Jesus for upp till Jerusalem.
Vid Fårporten i Jerusalem ligger en damm, på hebreiska kallad Betesda, och invid den finnas fem pelargångar.
I dessa lågo många sjuka, blinda, halta, förtvinade.
262820
Där fanns nu en man som hade varit sjuk i trettioåtta år.
Då Jesus fick se denne, där han låg, och fick veta att han redan lång tid hade varit sjuk, sade han till honom: »Vill du bliva frisk?»
Den sjuke svarade honom: »Herre, jag har ingen som hjälper mig ned i dammen, när vattnet har kommit i rörelse; och så stiger en annan ditned före mig, medan jag ännu är på väg.»
Jesus sade till honom: »Stå upp, tag din säng och gå.»
Och strax blev mannen frisk och tog sin säng och gick.
Men det var sabbat den dagen.
Därför sade judarna till mannen som hade blivit botad: »Det är sabbat; det är icke lovligt för dig att bära sängen.»
Men han svarade dem: »Den som gjorde mig frisk, han sade till mig: 'Tag din säng och gå.'»
Då frågade de honom: »Vem var den mannen som sade till dig att du skulle taga sin säng och gå?»
Men mannen som hade blivit botad visste icke vem det var; ty Jesus hade dragit sig undan, eftersom mycket folk var där på platsen. --
Sedan träffade Jesus honom i helgedomen och sade till honom: »Se, du har blivit frisk; synda icke härefter, på det att icke något värre må vederfaras dig.»
Mannen gick då bort och omtalade för judarna, att det var Jesus som hade gjort honom frisk.
Därför förföljde nu judarna Jesus, eftersom han gjorde sådant på sabbaten.
Men han svarade dem: »Min Fader verkar ännu alltjämt; så verkar ock jag.»
Och därför stodo judarna ännu mer efter att döda honom, eftersom han icke allenast ville göra sabbaten om intet, utan ock kallade Gud sin Fader och gjorde sig själv lik Gud.
Då talade Jesus åter och sade till dem: »Sannerligen, sannerligen säger jag eder: Sonen kan icke göra något av sig själv, utan han gör allenast vad han ser Fadern göra; ty vad han gör, det gör likaledes ock Sonen.
Ty Fadern älskar Sonen och låter honom se allt vad han själv gör; och större gärningar, än dessa äro, skall han låta honom se, så att I skolen förundra eder.
Ty såsom Fadern uppväcker döda och gör dem levande, så gör ock Sonen levande vilka han vill.
Icke heller dömer Fadern någon, utan all dom har han överlåtit åt Sonen,
för att alla skola ära Sonen såsom de ära Faderns.
Den som icke ärar Sonen, han ärar icke heller Fadern, som har sänt honom.
Sannerligen, sannerligen säger jag eder: Den som hör mina ord och tror honom som har sänt mig, han har evigt liv och kommer icke under någon dom, utan har övergått från döden till livet.
Sannerligen säger jag eder: Den stund kommer, jag, den är redan inne, så de döda skola höra Guds Sons röst, och de som höra den skola bliva levande.
Ty såsom Fadern har liv i sig själv, så har han ock givit åt Sonen att hava liv i sig själv.
Och han har givit honom makt att hålla dom, eftersom han är Människoson.
Förundren eder icke över detta.
Ty den stund kommer, då alla som äro i gravarna skola höra hans röst
och gå ut ur dem: de som hava gjort vad gott är skola uppstå till liv, och de som hava gjort vad ont är skola uppstå till dom.
Jag kan icke göra något av mig själv.
Såsom jag hör, så dömer jag; och min dom är rättvis, ty jag söker icke min vilja, utan dens vilja, som har sänt mig.
Om jag själv vittnar om mig, så gäller icke mitt vittnesbörd.
Men det är en annan som vittnar om mig, och jag vet att hans vittnesbörd om mig är sant.
I haven sänt bud till Johannes, och han har vittnat för sanningen,
Dock, det är icke av någon människa som jag tager emot vittnesbörd om mig; men jag säger detta, för att I skolen bliva frälsta.
Han var den brinnande, skinande lampan, och för en liten stund villen I fröjdas i dess ljus.
Men jag har ett vittnesbörd om mig, som är förmer än Johannes' vittnesbörd: de gärningar som Fadern har givit mig att fullborda, just de gärningar som jag gör, de vittna om mig, att Fadern har sänt mig.
Ja, Fadern, som har sänt mig, han har själv vittnat om mig.
Hans röst haven I aldrig någonsin hört, ej heller haven I sett hans gestalt,
och hans ord haven I icke låtit förbliva i eder.
Ty den han har sänt, honom tron I icke.
I rannsaken skrifterna, därför att I menen eder i dem hava evigt liv; och det är dessa som vittna om mig.
Men I viljen icke komma till mig för att få liv.
Jag tager icke emot pris av människor;
men jag känner eder och vet att I icke haven Guds kärlek i eder.
Jag har kommit i min Faders namn, och I tagen icke emot mig; kommer en annan i sitt eget namn, honom skolen I nog mottaga.
Huru skullen I kunna tro, I som tagen emot pris av varandra och icke söken det pris som kommer från honom som allena är Gud?
Menen icke att det är jag som skall anklaga eder hos Fadern.
Den som anklagar eder är Moses, han till vilken I sätten edert hopp.
Trodden I Moses, så skullen I ju tro mig, ty om mig har han skrivit.
Men tron I icke hans skrifter, huru skolen I då kunna tro mina ord?»
Därefter for Jesus över Galileiska sjön, »Tiberias' sjö».
Och mycket folk följde efter honom, därför att de sågo de tecken som han gjorde med de sjuka.
Men Jesus gick upp på berget och satte sig där med sina lärjungar.
Och påsken, judarnas högtid, var nära.
Då nu Jesus lyfte upp sina ögon och såg att mycket folk kom till honom, sade han till Filippus: »Varifrån skola vi köpa bröd, så att dessa få äta?»
Men detta sade han för att sätta honom på prov, ty själv visste han vad han skulle göra.
Filippus svarade honom: »Bröd för två hundra silverpenningar vore icke nog för att var och en skulle få ett litet stycke.»
Då sade till honom en annan av hans lärjungar, Andreas, Simon Petrus' broder:
»Här är en gosse som har fem kornbröd och två fiskar; men vad förslår det för så många?»
Jesus sade: »Låten folket lägga sig här.»
Och på det stället var mycket gräs.
Då lägrade sig männen där, och deras antal var vid pass fem tusen.
Därefter tog Jesus bröden och tackade Gud och delade ut åt dem som hade lagt sig ned där, likaledes ock av fiskarna, så mycket de ville hava.
Och när de voro mätta, sade han till sina lärjungar: »Samlen tillhopa de överblivna styckena, så att intet förfares.»
Då samlade de dem tillhopa och fyllde tolv korgar med stycken, som av de fem kornbröden hade blivit över efter dem som hade ätit.
Då nu människorna hade det tecken som han hade gjort, sade de: »Denne är förvisso Profeten som skulle komma i världen.»
När då Jesus märkte att de tänkte komma och med våld föra honom med sig och göra honom till konung, drog han sig åter undan till berget, helt allena.
Men när det blev afton, gingo hans lärjungar ned till sjön
och stego i en båt för att fara över sjön till Kapernaum.
Det hade då redan blivit mörkt, och Jesus hade ännu icke kommit till dem;
och sjön gick hög, ty det blåste hårt.
När de så hade rott vid pass tjugufem eller trettio stadier, fingo de se Jesus komma gående på sjön och nalkas båten.
Då blevo de förskräckta.
Men han sade till dem: »Det är jag; varen icke förskräckta.»
De ville då taga honom upp i båten; och strax var båten framme vid landet dit de foro.
Dagen därefter hände sig detta.
Folket som stod kvar på andra sidan sjön hade lagt märke till att där icke fanns mer än en enda båt, och att Jesus icke hade stigit i den båten med sina lärjungar, utan att lärjungarna hade farit bort allena.
Andra båtar hade likväl kommit från Tiberias och lagt till nära det ställe där folket bespisades efter det att Herren hade uttalat tacksägelsen.
När alltså folket nu såg att Jesus icke var där, ej heller hans lärjungar, stego de själva i båtarna och foro till Kapernaum för att söka efter Jesus.
Och då de funno honom där på andra sidan sjön, frågade de honom: »Rabbi, när kom du hit?»
Jesus svarade dem och sade: »Sannerligen, sannerligen säger jag eder: I söken mig icke därför att I haven sett tecken, utan därför att I fingen äta av bröden och bleven mätta.
Verken icke för att få den mat som förgås, utan för att få den mat som förbliver och har med sig evigt liv, den som Människosonen skall giva eder; ty honom har Fadern, Gud själv, låtit undfå sitt insegel.»
Då sade de till honom: »Vad skola vi göra för att utföra Guds gärningar?»
Jesus svarade och sade till dem: »Detta är Guds gärning, att I tron på den han har sänt.»
De sade till honom: »Vad för tecken gör du då?
Låt oss se något tecken, så att vi kunna tro dig.
Vilken gärning utför du?
Våra fäder fingo äta manna i öknen, såsom det är skrivet: 'Han gav dem bröd från himmelen att äta.'»
Då svarade Jesus dem: »Sannerligen, sannerligen säger jag eder: Det är icke Moses som har givit eder brödet från himmelen, men det är min Fader som giver eder det rätta brödet från himmelen.
Ty Guds bröd är det bröd som kommer ned från himmelen och giver världen liv.»
Då sade de till honom: »Herre, giv oss alltid det brödet.»
Jesus svarade: »Jag är livets bröd.
Den som kommer till mig, han skall aldrig hungra, och den som tror på mig, han skall aldrig törsta.
Men det är såsom jag har sagt eder: fastän I haven sett mig, tron I dock icke.
Allt vad min Fader giver mig, det kommer till mig; och den som kommer till mig, honom skall jag sannerligen icke kasta ut.
Ty jag har kommit ned från himmelen, icke för att göra min vilja, utan för att göra dens vilja, som har sänt mig.
Och detta är dens vilja, som har sänt mig, att jag icke skall låta någon enda gå förlorad av dem som han har givit mig, utan att jag skall låta dem uppstå på den yttersta dagen.
Ja, detta är min Faders vilja, att var och en som ser Sonen och tror på honom, han skall hava evigt liv, och att jag skall låta honom uppstå på den yttersta dagen.»
Då knorrade judarna över honom, därför att han hade sagt: »Jag är det bröd som har kommit ned från himmelen.»
Och de sade: »Är denne icke Jesus, Josefs son, vilkens fader och moder vi känna?
Huru kan han då säga: 'Jag har kommit ned från himmelen'?»
Jesus svarade och sade till dem: »Knorren icke eder emellan.
Ingen kan komma till mig, om icke Fadern, som har sänt mig, drager honom; och jag skall låta honom uppstå på den yttersta dagen.
Det är skrivet hos profeterna: 'De skola alla hava fått lärdom av Gud.'
Var och en som har lyssnat till Fadern och lärt av honom, han kommer till mig.
Icke som om någon skulle hava sett Fadern, utom den som är från Gud; han har sett Fadern.
Sannerligen, sannerligen säger jag eder: Den som tror, han har evigt liv.
Jag är livets bröd.
Edra fäder åto manna i öknen, och de dogo.
Men med det bröd som kommer ned från himmelen är det så, att om någon äter därav, så skall han icke dö.
Jag är det levande brödet som har kommit ned från himmelen.
Om någon äter av det brödet, så skall han leva till evig tid.
Och det bröd som jag skall giva är mitt kött; och jag giver det, för att världen skall leva.»
Då tvistade judarna med varandra och sade: »Huru skulle denne kunna giva oss sitt kött att äta?»
Jesus sade då till dem: »Sannerligen, sannerligen säger jag eder: Om I icke äten Människosonens kött och dricken hans blod, så haven I icke liv i eder.
Den som äter mitt kött och dricker mitt blod, han har evigt liv, och jag skall låta honom uppstå på den yttersta dagen.
Ty mitt kött är sannskyldig mat, och mitt blod är sannskyldig dryck.
Den som äter mitt kött och dricker mitt blod, han förbliver i mig, och jag förbliver i honom.
Såsom Fadern, han som är den levande, har sänt mig, och såsom jag lever genom Fadern, så skall ock den som äter mig leva genom mig.
Så är det med det bröd som har kommit ned från himmelen.
Det är icke såsom det fäderna fingo äta, vilka sedan dogo; den som äter detta bröd, han skall leva till evig tid.»
Detta sade han, när han undervisade i synagogan i Kapernaum.
Många av hans lärjungar, som hörde detta, sade då: »Detta är ett hårt tal; vem står ut med att höra på honom?»
Men Jesus visste inom sig att hans lärjungar knorrade över detta; och han sade till dem: »Är detta för eder en stötesten?
Vad skolen I då säga, om I fån se Människosonen uppstiga dit där han förut var? --
Det är anden som gör levande; köttet är till intet gagneligt.
De ord som jag har talat till eder äro ande och äro liv.
Men bland eder finnas några som icke tro.»
Jesus visste nämligen från begynnelsen vilka de voro som icke trodde, så ock vilken den var som skulle förråda honom.
Och han tillade: »Fördenskull har jag sagt eder att ingen kan komma till mig, om det icke bliver honom givet av Fadern.»
För detta tals skull drogo sig många av hans lärjungar tillbaka, så att de icke längre vandrade med honom.
Då sade Jesus till de tolv: »Icke viljen väl också I gå bort?»
Simon Petrus svarade honom: »Herre, till vem skulle vi gå?
Du har det eviga livets ord,
och vi tro och förstå att du är Guds helige.»
Jesus svarade dem: »Har icke jag själv utvalt eder, I tolv?
Och likväl är en av eder en djävul.»
Detta sade han om Judas, Simon Iskariots son; ty det var denne som skulle förråda honom, och han var en av de tolv.
Därefter vandrade Jesus omkring i Galileen, ty i Judeen ville han icke vandra omkring, då nu judarna stodo efter att döda honom.
Men judarnas lövhyddohögtid var nu nära.
Då sade hans bröder till honom: »Begiv dig härifrån och gå till Judeen, så att också dina lärjungar få se de gärningar som du gör.
Ty ingen som vill vara känd bland människor utför sitt verk i hemlighet.
Då du nu gör sådana gärningar, så träd öppet fram för världen.»
Det var nämligen så, att icke ens hans bröder trodde på honom.
Då sade Jesus till dem: »Min tid är ännu icke kommen, men för eder är tiden alltid läglig.
Världen kan icke hata eder, men mig hatar hon, eftersom jag vittnar om henne, att hennes gärningar äro onda.
Gån I upp till högtiden; jag är icke stadd på väg upp till denna högtid, ty min tid är ännu icke fullbordad.»
Detta sade han till dem och stannade så kvar i Galileen.
Men när hans bröder hade gått upp till högtiden, då gick också han ditupp, dock icke öppet, utan likasom i hemlighet.
Och judarna sökte efter honom under högtiden och sade: »Var är han?»
Och bland folket talades i tysthet mycket om honom.
Somliga sade: »Han är en rättsinnig man», men andra sade: »Nej, han förvillar folket.»
Dock talade ingen öppet om honom, av fruktan för judarna.
Men när redan halva högtiden var förliden, gick Jesus upp i helgedomen och undervisade.
Då förundrade sig judarna och sade: »Varifrån har denne sin lärdom, han som icke har fått undervisning?»
Jesus svarade dem och sade: »Min lära är icke min, utan hans som har sänt mig.
Om någon vill göra hans vilja, så skall han förstå om denna lära är från Gud, eller om jag talar av mig själv.
Den som talar av sig själv, han söker sin egen ära; men den som söker dens ära, som har sänt honom, han är sannfärdig, och orättfärdighet finnes icke i honom. --
Har icke Moses givit eder lagen?
Och likväl fullgör ingen av eder lagen.
Varför stån I efter att döda mig?»
Folket svarade: »Du är besatt av en ond ande.
Vem står efter att döda dig?»
Jesus svarade och sade till dem: »En gärning allenast gjorde jag, och alla förundren I eder över den.
Moses har givit eder omskärelsen -- icke som om den vore ifrån Moses, ty den är ifrån fäderna -- och så omskären I människor också på en sabbat.
Om nu en människa undfår omskärelsen på en sabbat, för att Moses' lag icke skall göras om intet, huru kunnen I då vredgas på mig, därför att jag på en sabbat gjorde en människa hel och frisk?
Dömen icke efter skenet, utan dömen en rätt dom.»
Då sade några av folket i Jerusalem: »Är det icke denne som de stå efter att döda?
Och ändå får han tala fritt, utan att de säga något till honom.
Hava då rådsherrarna verkligen blivit förvissade om att denne är Messias?
Dock, denne känna vi, och vi veta varifrån han är; men när Messias kommer, känner ingen varifrån han är.»
Då sade Jesus med hög röst, där han undervisade i helgedomen: »Javäl, I kännen mig, och I veten varifrån jag är.
Likväl har jag icke kommit av mig själv, men han som har sänt mig är en som verkligen har myndighet att sända, han som I icke kännen.
Men jag känner honom, ty från honom är jag kommen, och han har sänt mig.»
Då ville de gripa honom; dock kom ingen med sin hand vid honom, ty hans stund var ännu icke kommen.
Men många av folket trodde på honom, och de sade: »Icke skall väl Messias, när han kommer, göra flera tecken än denne har gjort?»
Sådant fingo fariséerna höra folket i tysthet tala om honom.
Då sände översteprästerna och fariséerna ut rättstjänare för att gripa honom.
Men Jesus sade: »Ännu en liten tid är jag hos eder; sedan går jag bort till honom som har sänt mig.
I skolen då söka efter mig, men I skolen icke finna mig, och där jag är, dit kunnen I icke komma.»
Då sade judarna till varandra: »Vart tänker denne gå, eftersom vi icke skola kunna finna honom?
Månne han tänker gå till dem som bo kringspridda bland grekerna?
Tänker han då undervisa grekerna?
Vad betyder det ord som han sade: 'I skolen söka efter mig, men I skolen icke finna mig, och där jag är, dit kunnen I icke komma'?»
På den sista dagen i högtiden, som ock var den förnämsta, stod Jesus där och ropade och sade: »Om någon törstar, så komme han till mig och dricke.
Den som tror på mig, av hans innersta skola strömmar av levande vatten flyta fram, såsom skriften säger.»
Detta sade han om Anden, vilken de som trodde på honom skulle undfå; ty ande var då ännu icke given, eftersom Jesus ännu icke hade blivit förhärligad.
Några av folket, som hörde dessa ord, sade då: »Denne är förvisso Profeten.»
Andra sade: »Han är Messias.»
Andra åter sade: »Icke kommer väl Messias från Galileen?
Säger icke skriften att Messias skall komma av Davids säd och från den lilla staden Betlehem, där David bodde?
Så uppstodo för hans skull stridiga meningar bland folket,
och somliga av dem ville gripa honom; dock kom ingen med sin hand vid honom.
När sedan rättstjänarna kommo tillbaka till översteprästerna och fariséerna, frågade dessa dem: »Varför haven I icke fört honom hit?»
Tjänarna svarade: »Aldrig har någon människa talat, som den mannen talar.»
Då svarade fariséerna dem: »Haven nu också I blivit förvillade?
Har då någon av rådsherrarna trott på honom?
Eller någon av fariséerna?
Nej; men detta folk, som icke känner lagen, det är förbannat.
Då sade Nikodemus till dem, han som förut hade besökt honom, och som själv var en av dem:
»Icke dömer väl vår lag någon, utan att man först har förhört honom och utrönt vad han förehar?»
De svarade och sade till honom: »Kanske också du är från Galileen?
Rannsaka, så skall du finna att ingen profet kommer från Galileen.»
h de gingo hem, var och en till sitt.
Och Jesus gick ut till Oljeberget.
Men i dagbräckningen kom han åter till helgedomen.
Då förde översteprästerna och fariséerna dit en kvinna som hade blivit beträdd med äktenskapsbrott; och när de hade lett henne fram,
sade de till honom: »Mästare, denna kvinna har på bar gärning blivit beträdd med äktenskapsbrott.
Nu bjuder Moses i lagen att sådana skola stenas.
Vad säger då du?»
Detta sade de för att snärja honom, på det att de skulle få något att anklaga honom för.
Då böjde Jesus sig ned och skrev med fingret på jorden.
Men när de stodo fast vid sin fråga, reste han sig upp och sade till dem: »Den av eder som är utan synd, han kaste första stenen på henne.»
Sedan böjde han sig åter ned och skrev på jorden.
När de hörde detta, gingo de ut, den ene efter den andre, först de äldsta, och Jesus blev lämnad allena med kvinnan, som stod där kvar.
Då såg Jesus upp och sade till kvinnan: »Var äro de andra?
Har ingen dömt dig?»
Hon svarade: »Herre, ingen.»
Då sade han till henne: »Icke heller jag dömer dig.
Gå, och synda icke härefter.»]
Åter talade Jesus till dem och sade: »Jag är världens ljus; den som följer mig, han skall förvisso icke vandra i mörkret, utan skall hava livets ljus.»
Då sade fariséerna till honom: »Du vittnar om dig själv; ditt vittnesbörd gäller icke.»
Jesus svarade och sade till dem: »Om jag än vittnar om mig själv, så gäller dock mitt vittnesbörd, ty jag vet varifrån jag har kommit, och vart jag går; men I veten icke varifrån jag kommer, eller vart jag går.
I dömen efter köttet; jag dömer ingen.
Och om jag än dömer, så är min dom en rätt dom, ty jag är därvid icke ensam, utan med mig är han som har sänt mig.
I eder lag är ju ock skrivet att vad två människor vittna, det gäller såsom sant.
Här är nu jag som vittnar om mig; om mig vittnar också Fadern, som har sänt mig.
Då sade de till honom: »Var är då din Fader?»
Jesus svarade: »I kännen varken mig eller min Fader.
Om I känden mig, så känden I ock min Fader.»
Det var på det ställe där offerkistorna stodo som han talade dessa ord, medan han undervisade i helgedomen; men ingen bar hand på honom, ty hans stund var ännu icke kommen.
Åter sade han till dem: »Jag går bort, och I skolen då söka efter mig; men I skolen dö i eder synd.
Dig jag går, dit kunnen I icke komma.»
Då sade judarna: »Icke vill han väl dräpa sig själv, eftersom han säger: 'Dit jag går, dit kunnen I icke komma'?»
Men han svarade dem: »I ären härnedifrån, jag är ovanifrån; I ären av denna världen, jag är icke av denna världen.
Därför sade jag till eder att I skullen dö i edra synder; ty om I icke tron att jag är den jag är, så skolen I dö i edra synder.»
Då frågade de honom: »Vem är du då?»
Jesus svarade dem: »Det som jag redan från begynnelsen har uttalat för eder.
Mycket har jag ännu att tala och att döma i fråga om eder.
Men han som har sänt mig är sannfärdig, och vad jag har hört av honom, det talar jag ut inför världen.»
Men de förstodo icke att det var om Fadern som han talade till dem.
Då sade Jesus: »När I haven upphöjt Människosonen, då skolen I första att jag är den jag är, och att jag icke gör något av mig själv, utan talar detta såsom Fadern har lärt mig.
Och han som har sänt mig är med mig; han har icke lämnat mig allena, eftersom jag alltid gör vad honom behagar.»
När han talade detta, kommo många till tro på honom.
Då sade Jesus till de judar som hade satt tro till honom: »Om I förbliven i mitt ord, så ären I i sanning mina lärjungar;
Och I skolen då förstå sanningen, och sanningen skall göra eder fria.»
De svarade honom: »Vi äro Abrahams säd och hava aldrig varit trälar under någon.
Huru kan du då säga: 'I skolen bliva fria'?»
Jesus svarade dem: »Sannerligen, sannerligen säger jag eder: Var och en som gör synd, han är syndens träl.
Men trälen får icke förbliva i huset för alltid; sonen får förbliva där för alltid.
Om nu Sonen gör eder fria, så bliven i verkligen fria.
Jag vet att I ären Abrahams säd; men I stån efter att döda mig, eftersom mitt ord icke får någon ingång i eder.
Jag talar vad jag har sett hos min Fader; så gören ock I vad I haven hört av eder fader.»
De svarade och sade till honom: »Vår fader är ju Abraham.»
Jesus svarade till dem: »Ären I Abrahams barn, så gören ock Abrahams gärningar.
Men nu stån I efter att döda mig, en man som har sagt eder sanningen, såsom jag har hört den av Gud.
Så handlade icke Abraham.
Nej, I gören eder faders gärningar.»
De sade till honom: »Vi äro icke födda i äktenskapsbrott.
Vi hava Gud till fader och ingen annan.»
Jesus svarade dem: »Vore Gud eder fader, så älskaden I ju mig, ty från Gud har jag utgått, och från honom är jag kommen.
Ja, jag har icke kommit av mig själv, utan det är han som har sänt mig.
Varför fatten I då icke vad jag talar?
Jo, därför att I icke 'stån ut med' att höra på mitt ord.
I haven djävulen till eder fader, och vad eder fader har begär till, det viljen i göra.
Han har varit en mandråpare från begynnelsen, och i sanningen står han icke, ty sanning finnes icke i honom.
När han talar lögn, då talar han av sitt eget, ty han är en lögnare, ja, lögnens fader.
Men mig tron I icke, just därför att jag talar sanning.
Vilken av eder kan överbevisa mig om någon synd?
Om jag alltså talar sanning, varför tron I mig då icke?
Den som är av Gud, han lyssnar till Guds ord; och det är därför att I icke ären av Gud som I icke lyssnen därtill.
Judarna svarade och sade till honom: »Hava vi icke rätt, då vi säga att du är en samarit och är besatt av en ond ande?»
Jesus svarade: »Jag är icke besatt av någon ond ande; fastmer hedrar jag min Fader.
I åter skymfen mig.
Men jag söker icke min egen ära; en finnes dock som söker den och som dömer.
Sannerligen, sannerligen säger jag eder: Den som håller mitt ord, han skall aldrig någonsin se döden.»
Judarna sade till honom: »Nu förstå vi att du är besatt av en ond ande.
Abraham har dött, så ock profeterna, och likväl säger du: 'Den som håller mitt ord, han skall aldrig någonsin smaka döden.'
Icke är väl du förmer än vår Fader Abraham?
Och han har ju dött.
Profeterna hava också dött.
Till vem gör du då dig själv?»
Jesus svarade: »Om jag själv ville skaffa mig ära, så vore min ära intet; men det är min Fader som förlänar mig ära, han som I säger vara eder Gud.
Dock, I haven icke lärt känna honom, men jag känner honom; och om jag sade att jag icke kände honom, så bleve jag en lögnare likasom I; men jag känner honom och håller hans ord.
Abraham, eder fader, fröjdade sig över att han skulle få se min dag.
Han fick se den och blev glad.»
Då sade judarna till honom: »Femtio år gammal är du icke ännu, och Abraham har du sett!»
Jesus sade till dem: »Sannerligen, sannerligen säger jag eder: Förrän Abraham blev till, är jag.»
Då togo de upp stenar för att kasta på honom.
Men Jesus gömde sig undan och gick sedan ut ur helgedomen.
När han nu gick vägen fram, fick han se en man som var född blind.
Då frågade hans lärjungar honom och sade: »Rabbi, vilken har syndat, denne eller hans föräldrar, så att han har blivit född blind?»
Jesus svarade: »Det är varken denne som har syndat eller hans föräldrar, utan så har skett, för att Guds gärningar skulle uppenbaras på honom.
Medan dagen varar, måste vi göra dens gärningar, som har sänt mig; natten kommer, då ingen kan verka.
Så länge jag är i världen, är jag världens ljus.»
När han hade sagt detta, spottade han på jorden och gjorde en deg av spotten och lade degen på mannens ögon
och sade till honom: »Gå bort och två dig i dammen Siloam» (det betyder utsänd).
Mannen gick då dit och tvådde sig; och när han kom igen, kunde han se.
Då sade grannarna och andra som förut hade sett honom såsom tiggare: »Är detta icke den man som att och tiggde?»
Somliga svarade: »Det är han.»
Andra sade: »Nej, men han är lik honom.»
Själv sade han: »Jag är den mannen.»
Och de frågade honom: »Huru blevo då dina ögon öppnade?»
Han svarade: »Den man som heter Jesus gjorde en deg och smorde därmed mina ögon och sade till mig: 'Gå bort till Siloam och två dig.'
Jag gick då dit och tvådde mig, och så fick jag min syn.»
De frågade honom: »Var är den mannen?»
Han svarade: »Det vet jag icke.»
Då förde de honom, mannen som förut hade varit blind, bort till fariséerna.
Och det var sabbat den dag då Jesus gjorde degen och öppnade hans ögon.
När nu jämväl fariséerna i sin ordning frågade honom huru han hade fått sin syn, svarade han dem: »Han lade en deg på mina ögon, och jag fick två mig, och nu kan jag se.»
Då sade några av fariséerna: »Den mannen är icke från Gud, eftersom han icke håller sabbaten.»
Andra sade: »Huru skulle någon som är en syndare kunna göra sådana tecken?»
Så funnos bland dem stridiga meningar.
Då frågade de åter den blinde: »Vad säger du själv om honom, då det ju var dina ögon han öppnade?»
Han svarade: »En profet är han.»
Men judarna trodde icke att han hade varit blind och fått sin syn, förrän de hade kallat till sig mannen föräldrar, hans som hade fått sin syn.
Dem frågade de och sade: »Är detta eder son, den som I sägen vara född blind?
Huru kommer det då till, att han nu kan se?»
Då svarade han föräldrar och sade: »Att denne är vår son, och att han föddes blind, det veta vi.
Men huru han nu kan se, det veta vi icke, ej heller veta vi vem som har öppnat hans ögon.
Frågen honom själv; han är gammal nog, han må själv tala för sig.»
Detta sade hans föräldrar, därför att de fruktade judarna; ty judarna hade redan kommit överens om att den som bekände Jesus vara Messias, han skulle utstötas ur synagogan.
Därför var det som hans föräldrar sade: »Han är gammal nog; frågen honom själv.»
Då kallade de för andra gången till sig mannen som hade varit blind och sade till honom: »Säg nu sanningen, Gud till pris.
Vi veta att denne man är en syndare.»
Han svarade: »Om han är en syndare vet jag icke; ett vet jag: att jag, som var blind, nu kan se.»
Då frågade de honom: »Vad gjorde han med dig?
På vad sätt öppnade han dina ögon?»
Han svarade dem: »Jag har ju redan sagt eder det, men I hörden icke på mig.
Varför viljen I då åter höra det?
Kanske viljen också I bliva hans lärjungar?»
Då bannade de honom och sade: »Du är själv hans lärjunge; vi äro Moses' lärjungar.
Till Moses har Gud talat, det veta vi; men varifrån denne är, det veta vi icke.»
Mannen svarade och sade till dem: »Ja, däri ligger det förunderliga, att I icke veten varifrån han är, och ändå har han öppnat mina ögon.
Vi veta ju att Gud icke hör syndare, men också att om någon är gudfruktig och gör hans vilja, då hör han honom.
Aldrig förut har man hört att någon har öppnat ögonen på en som föddes blind.
Vore denne icke från Gud, så kunde han intet göra.»
De svarade och sade till honom: »Du är hel och hållen född i synd, och du vill undervisa oss!»
Och så drevo de ut honom.
Jesus fick sedan höra att de hade drivit ut honom, och när han så träffade honom, sade han: »Tror du på Människosonen?»
Han svarade och sade: »Herre, vem är han då?
Säg mig det, så att jag kan tro på honom.»
Jesus sade till honom: »Du har sett honom; det är han som talar med dig.»
Då sade han: »Herre, jag tror.»
Och han föll ned för honom.
Och Jesus sade: »Till en dom har jag kommit hit i världen, för att de som icke se skola varda seende, och för att de som se skola varda blinda.»
När några fariséer som voro i hans närhet hörde detta, sade de till honom: »Äro då kanske också vi blinda?»
Jesus svarade dem: »Voren I blinda, så haden I icke synd.
Men nu sägen I: 'Vi se', därför står eder synd kvar.»
»Sannerligen, sannerligen säger jag eder: Den som icke går in i fårahuset genom dörren, utan stiger in någon annan väg, han är en tjuv och en rövare.
Men den som går in genom dörren, han är fårens herde.
För honom öppnar dörrvaktaren, och fåren lyssna till hans röst, och han kallar sina får vid namn och för dem ut.
Och när han har släppt ut alla sina får, går han framför dem, och fåren följa honom, ty de känna hans röst.
Men en främmande följa de alls icke, utan fly bort ifrån honom, ty de känna icke de främmandes röst.»
Så talade Jesus till dem i förtäckta ord; men de förstodo icke vad det var som han talade till dem.
Åter sade Jesus till dem: »Sannerligen, sannerligen säger jag eder: Jag är dörren in till fåren.
Alla de som hava kommit före mig äro tjuvar och rövare, men fåren hava icke lyssnat till dem.
Jag är dörren; den som går in genom mig, han skall bliva frälst, och han skall få gå ut och in och skall finna bete.
Tjuven kommer allenast för att stjäla och slakta och förgöra.
Jag har kommit, för att de skola hava liv och hava över nog.
Jag är den gode herden.
En god herde giver sitt liv för fåren.
Men den som är lejd och icke är herden själv, när han, den som fåren icke tillhöra, ser ulven komma, då övergiver han fåren och flyr, och ulven rövar bort dem och förskingrar dem.
Han är ju lejd och frågar icke efter fåren.
Jag är den gode herden, och jag känner mina får, och mina får känna mig,
såsom Fadern känner mig, och såsom jag känner Fadern; och jag giver mitt liv för fåren.
Jag har ock andra får, som icke höra till detta fårahus; också dem måste jag draga till mig, och de skola lyssna till min röst.
Så skall det bliva en hjord och en herde.
Därför älskar Fadern mig, att jag giver mitt liv -- för att sedan taga igen det.
Ingen tager det ifrån mig, utan jag giver det av fri vilja.
Jag har makt att giva det, och jag har makt att taga igen det.
Det budet har jag fått av min Fader.»
För dessa ords skull uppstodo åter stridiga meningar bland judarna.
Många av dem sade: »Han är besatt av en ond ande och är från sina sinnen.
Varför hören I på honom?»
Andra åter sade: »Sådana ord talar icke den som är besatt.
Icke kan väl en ond ande öppna blindas ögon?»
Därefter inföll tempelinvigningens högtid i Jerusalem.
Det var nu vinter,
och Jesus gick fram och åter i Salomos pelargång i helgedomen.
Då samlade sig judarna omkring honom och sade till honom: »Huru länge vill du hålla oss i ovisshet?
Om du är Messias, så säg oss det öppet.»
Jesus svarade dem: »Jag har sagt eder det, men I tron mig icke.
De gärningar som jag gör i min Faders namn, de vittna om mig.
Men I tron mig icke, ty I ären icke av mina får.
Mina får lyssna till min röst, och jag känner dem, och de följa mig.
Och jag giver dem evigt liv, och de skola aldrig någonsin förgås, och ingen skall rycka dem ur min hand.
Min Fader, som har givit mig dem, är större än alla, och ingen kan rycka dem ur min Faders hand.
Jag och Fadern äro ett.»
Då togo judarna åter upp stenar för att stena honom.
Men Jesus sade till dem: »Många goda gärningar, som komma från min Fader, har jag låtit eder se.
För vilken av dessa gärningar är det som I viljen stena mig?»
Judarna svarade honom: »Det är icke för någon god gärnings skull som vi vilja stena dig, utan därför att du hädar och gör dig själv till Gud, du som är en människa.»
Jesus svarade dem: »Det är ju så skrivet i eder lag: 'Jag har sagt att I ären gudar'.
Om han nu har kallat för gudar dem som Guds ord kom till -- och skriften kan ju icke bliva om intet --
huru kunnen då I, på den grund att jag har sagt mig vara Guds Son, anklaga mig för hädelse, mig som Fadern har helgat och sänt i världen?
Gör jag icke min Faders gärningar, så tron mig icke.
Men gör jag dem, så tron gärningarna, om I än icke tron mig; då skolen I fatta och förstå att Fadern är i mig, och att jag är i Fadern.»
Då ville de åter gripa honom, men han gick sin väg, undan deras händer.
Sedan begav han sig åter bort till det ställe på andra sidan Jordan, där Johannes först hade döpt, och stannade kvar där.
Och många kommo till honom.
Och de sade: »Väl gjorde Johannes intet tecken, men allt vad Johannes sade om denne var sant.»
Och många kommo där till tro på honom.
Och en man vid namn Lasarus låg sjuk; han var från Betania, den by där Maria och hennes syster Marta bodde.
Det var den Maria som smorde Herren med smörjelse och torkade hans fötter med sitt hår.
Och nu låg hennes broder Lasarus sjuk.
Då sände systrarna bud till Jesus och läto säga: »Herre, se, han som du har så kär ligger sjuk.»
När Jesus hörde detta, sade han: »Den sjukdomen är icke till döds, utan till Guds förhärligande, så att Guds Son genom den bliver förhärligad.»
Och Jesus hade Marta och hennes syster och Lasarus kära.
När han nu hörde att denne låg sjuk, stannade han först två dagar där han var;
men därefter sade han till lärjungarna: »Låt oss gå tillbaka till Judeen.»
Lärjungarna sade till honom: »Rabbi, nyligen ville judarna stena dig, och åter går du dit?»
Jesus svarade: »Dagen har ju tolv timmar; den som vandrar om dagen, han stöter sig icke, ty han ser då denna världens ljus.
Men den som vandrar om natten, han stöter sig, ty han har då intet som lyser honom.»
Sedan han hade talat detta, sade han ytterligare till dem: »Lasarus, vår vän, har somnat in; men jag går för att väcka upp honom ur sömnen.»
Då sade hans lärjungar till honom: »Herre, sover han, så bliver han frisk igen.»
Men Jesus hade talat om hans död; de åter menade att han talade om vanlig sömn.
Då sade Jesus öppet till dem: »Lasarus är död.
Och för eder skull, för att I skolen tro, gläder jag mig över att jag icke var där.
Men låt oss nu gå till honom.»
Då sade Tomas, som kallades Didymus, till de andra lärjungarna: »Låt oss gå med, för att vi må dö med honom.»
När så Jesus kom dit, fann han att den döde redan hade legat fyra dagar i graven.
Nu låg Betania nära Jerusalem, vid pass femton stadier därifrån,
och många judar hade kommit till Marta och Maria för att trösta dem i sorgen över deras broder.
Då nu Maria fick höra att Jesus kom, gick hon honom till mötes; men Maria satt kvar hemma.
Och Marta sade till Jesus: »Herre, hade du varit här, så vore min broder icke död.
Men jag vet ändå att allt vad du beder Gud om, det skall Gud giva dig.»
Jesus sade till henne: »Din broder skall stå upp igen.»
Marta svarade honom: »Jag vet att han skall stå upp, vid uppståndelsen på den yttersta dagen.»
Jesus svarade till henne: »Jag är uppståndelsen och livet.
Den som tror på mig, han skall leva, om han än dör;
och var och en som lever och tror på mig, han skall aldrig någonsin dö.
Tror du detta?»
Hon svarade honom: »Ja, Herre, jag tror att du är Messias, Guds Son, han som skulle komma i världen.»
När hon hade sagt detta, gick hon bort och kallade på Maria, sin syster, och sade hemligen till henne: »Mästaren är här och kallar dig till sig.»
När hon hörde detta, stod hon strax upp och gick åstad till honom.
Men Jesus hade ännu icke kommit in i byn, utan var kvar på det ställe där Marta hade mött honom.
Då nu de judar, som voro inne i huset hos Maria för att trösta henne, sågo att hon så hastigt stod upp och gick ut, följde de henne, i tanke att hon gick till graven för att gråta där.
När så Maria kom till det ställe där Jesus var och fick se honom, föll hon ned för hans fötter och sade till honom: »Herre, hade du varit där, så vore min broder icke död.»
Då nu Jesus såg henne gråta och såg jämväl att de judar, som hade kommit med henne, gräto, upptändes han i sin ande och blev upprörd
och frågade: »Var haven I lagt honom?»
De svarade honom: »Herre, kom och se.»
Och Jesus grät.
Då sade judarna: »Se huru kär han hade honom!»
Men somliga av dem sade:
»Kunde icke han, som öppnade den blindes ögon, ock hava så gjort att denne icke hade dött?»
Då upptändes Jesus åter i sitt innersta och gick bort till graven.
Den var urholkad i berget, och en sten låg framför ingången.
Jesus sade: »Tagen bort stenen.»
Då sade den dödes syster Marta till honom: »Herre, han luktar redan, ty han har varit död i fyra dygn.»
Jesus svarade henne: »Sade jag dig icke, att om du trodde, skulle du få se Guds härlighet?»
Då togo de bort stenen.
Och Jesus lyfte upp sina ögon och sade: »Fader, jag tackar dig för att du har hört mig.
Jag visste ju förut att du alltid hör mig; men för folkets skull, som står här omkring, säger jag detta, för att de skola tro att det är du som har sänt mig.»
När han hade sagt detta, ropade han med hög röst: »Lasarus, kom ut.»
Och han som hade varit död kom ut, med händer och fötter inlindade i bindlar och med ansiktet inhöljt i en duk.
Jesus sade till dem: »Lösen honom, och låten honom gå.»
Många judar, som hade kommit till Maria och hade sett vad Jesus hade gjort, trodde då på honom.
Men några av dem gingo bort till fariséerna och omtalade för dem vad Jesus hade gjort.
Då sammankallade översteprästerna och fariséerna en rådsförsamling och sade: »Vad skola vi taga oss till?
Denne man gör ju många tecken.
Om vi skola låta honom så fortfara, skola alla tro på honom, och romarna komma då att taga ifrån oss både land och folk.»
Men en av dem, Kaifas, som var överstepräst för det året, sade till dem: »I förstån intet,
och I besinnen icke huru mycket bättre det är för eder att en man dör för folket, än att hela folket förgås.»
Detta sade han icke av sig själv, utan genom profetisk ingivelse, eftersom han var överstepräst för det året; ty Jesus skulle dö för folket.
Ja, icke allenast »för folket»; han skulle dö också för att samla och förena Guds förskingrade barn.
Från den dagen var deras beslut fattat att döda honom.
Så vandrade då Jesus icke längre öppet bland judarna, utan drog sig undan till en stad som hette Efraim, på landsbygden, i närheten av öknen; där stannade han kvar med sina lärjungar.
Men judarnas påsk var nära, och många begåvo sig då, före påsken, från landsbygden upp till Jerusalem för att helga sig.
Och de sökte efter Jesus och sade till varandra, där de stodo i helgedom: »Vad menen I?
Skall han då alls icke komma till högtiden?»
Och översteprästerna och fariséerna hade utfärdat påbud om att den som finge veta var han fanns skulle giva det till känna, för att de måtte kunna gripa honom.
Sex dagar före påsk kom nu Jesus till Betania, där Lasarus bodde, han som av Jesus hade blivit uppväckt från de döda.
Där gjorde man då för honom ett gästabud, och Marta betjänade dem, men Lasarus var en av dem som lågo till bords jämte honom.
Då tog Maria ett skålpund smörjelse av dyrbar äkta nardus och smorde därmed Jesu fötter; sedan torkade hon hans fötter med sitt hår.
Och huset uppfylldes med vällukt av smörjelsen.
Men Judas Iskariot, en av hans lärjungar, den som skulle förråda honom, sade då:
»Varför sålde man icke hellre denna smörjelse för tre hundra silverpenningar och gav dessa åt de fattiga?»
Detta sade han, icke därför, att han frågade efter de fattiga, utan därför, att han var en tjuv och plägade taga vad som lades i penningpungen, vilken han hade om hand.
Men Jesus sade: »Låt henne vara; må hon få fullgöra detta för min begravningsdag.
De fattiga haven I ju alltid ibland eder, men mig haven I icke alltid.»
Nu hade det blivit känt för den stora hopen av judarna att Jesus var där, och de kommo dit, icke allenast för hans skull, utan ock för att se Lasarus, som han hade uppväckt från de döda.
Då beslöto översteprästerna att döda också Lasarus.
Ty för hans skull gingo många judar bort och trodde på Jesus.
När dagen därefter det myckna folk som hade kommit till högtiden fick höra att Jesus var på väg till Jerusalem,
togo de palmkvistar och gingo ut för att möta honom och ropade: »Hosianna!
Välsignad vare han som kommer, i Herrens namn, han som är Israels konung.»
Och Jesus fick sig en åsnefåle och satte sig upp på den, såsom det är skrivet:
»Frukta icke, du dotter Sion.
Se, din konung kommer, sittande på en åsninnas fåle.»
Detta förstodo hans lärjungar icke då strax, men när Jesus hade blivit förhärligad, då kommo de ihåg att detta var skrivet om honom, och att man hade gjort detta med honom.
Så gav nu folket honom sitt vittnesbörd, de som hade varit med honom, när han kallade Lasarus ut ur graven och uppväckte honom från de döda.
Därför kom också det övriga folket emot honom, eftersom de hörde att han hade gjort det tecknet.
Då sade fariséerna till varandra: »I sen att I alls intet kunnen uträtta; hela världen löper ju efter honom.»
Nu voro där ock några greker, av dem som plägade fara upp för att tillbedja under högtiden.
Dessa kommo till Filippus, som var från Betsaida i Galileen, och bådo honom och sade: »Herre, vi skulle vilja se Jesus.»
Filippus gick och sade detta till Andreas; Andreas och Filippus gingo och sade det till Jesus.
Jesus svarade dem och sade: »Stunden är kommen att Människosonen skall förhärligas.
Sannerligen, sannerligen säger jag eder: Om icke vetekornet faller i jorden och dör, så förbliver det ett ensamt korn; men om det dör, så bär det mycken frukt.
Den som älskar sitt liv, han mister det, men den som hatar sitt liv i denna världen, han skall behålla det och skall hava evigt liv.
Om någon vill tjäna mig, så följe han mig; och där jag är, där skall också min tjänare få vara.
Om någon tjänar mig, så skall min Fader ära honom.
Nu är min själ i ångest; vad skall jag väl säga?
Fader, fräls mig undan denna stund.
Dock, just därför har jag kommit till denna stund.
Fader, förhärliga ditt namn.»
Då kom en röst från himmelen: »Jag har redan förhärligat det, och jag skall ytterligare förhärliga det.»
Folket, som stod där och hörde detta, sade då: »Det var ett tordön.»
Andra sade: »Det var en ängel som talade med honom.»
Då svarade Jesus och sade: »Denna röst kom icke för min skull, utan för eder skull.»
Nu går en dom över denna världen, nu skall denna världens furste utkastas.
Och när jag har blivit upphöjd från jorden, skall jag draga alla till mig.»
Med dessa ord gav han till känna på vad sätt han skulle dö.
Då svarade folket honom: »Vi hava hört av lagen att Messias skall stanna kvar för alltid.
Huru kan du då säga att Människosonen måste bliva upphöjd?
Vad är väl detta för en Människoson?»
Jesus sade till dem: »Ännu en liten tid är ljuset ibland eder.
Vandren medan I haven ljuset, på det att mörkret icke må få makt med eder; den som vandrar i mörkret, han vet ju icke var han går.
Tron på ljuset, medan I haven ljuset, så att I bliven ljusets barn.»
Detta talade Jesus och gick sedan bort och dolde sig för dem.
Men fastän han hade gjort så många tecken inför dem, trodde de icke på honom.
Ty det ordet skulle fullbordas, som profeten Esaias säger: »Herre, vem trodde, vad som predikades för oss, och för vem var Herrens arm uppenbar?»
Alltså kunde de icke tro; Esaias säger ju ytterligare:
»Han har förblindat deras ögon och förstockat deras hjärtan, så att de icke kunna se med sina ögon eller förstå med sina hjärtan och omvända sig och bliva helade av mig.»
Detta kunde Esaias säga, eftersom han hade sett hans härlighet, när han talade med honom. --
Dock funnos jämväl bland rådsherrarna många som trodde på honom; men för fariséernas skulle ville de icke bekänna det, för att de icke skulle bliva utstötta ur synagogan.
Ty de skattade högre att bliva ärade av människor än att bliva ärade av Gud.
Men Jesus sade med hög röst: »Den som tror på mig, han tror icke på mig, utan på honom som har sänt mig.
Och den som ser mig, han ser honom som har sänt mig.
Såsom ett ljus har jag kommit i världen, för att ingen av dem som tro på mig skall förbliva i mörkret.
Om någon hör mina ord, men icke håller dem, så dömer icke jag honom; ty jag har icke kommit för att döma världen, utan för att frälsa världen.
Den som förkastar mig och icke tager emot mina ord, han har dock en domare över sig; det ord som jag har talat, det skall döma honom på den yttersta dagen.
Ty jag har icke talat av mig själv, utan Fadern, som har sänt mig, han har bjudit mig vad jag skall säga, och vad jag skall tala.
Och jag vet att hans bud är evigt liv; därför, vad jag talar, det talar jag såsom Fadern har sagt mig.»
Före påskhögtiden hände sig detta.
Jesus visste att stunden var kommen för honom att gå bort ifrån denna världen till Fadern; och såsom han allt hittills hade älskat sina egna här i världen, så gav han dem nu ett yttersta bevis på sin kärlek.
De höllo nu aftonmåltid, och djävulen hade redan ingivit Judas Iskariot, Simons son, i hjärtat att förråda Jesus.
Och Jesus visste att Fadern hade givit allt i hans händer, och att han hade gått ut från Gud och skulle gå till Gud.
Men han stod upp från måltiden och lade av sig överklädnaden och tog en linneduk och band den om sig.
Sedan slog han vatten i ett bäcken och begynte två lärjungarnas fötter och torkade dem med linneduken som han hade bundit om sig.
Så kom han till Simon Petrus.
Denne sade då till honom: »Herre, skulle du två mina fötter?»
Jesus svarade och sade till honom: »Vad jag gör förstår du icke nu, men framdeles skall du fatta det.»
Petrus sade till honom: »Aldrig någonsin skall du två mina fötter!»
Jesus svarade honom: »Om jag icke tvår dig, så har du ingen del med mig.»
Då sade Simon Petrus till honom: »Herre, icke allenast mina fötter, utan ock händer och huvud!»
Jesus svarade honom: »Den som är helt tvagen, han behöver allenast två fötterna; han är ju i övrigt hel och hållen ren.
Så ären ock I rena -- dock icke alla.»
Han visste nämligen vem det var som skulle förråda honom; därför sade han att de icke alla voro rena.
Sedan han nu hade tvagit deras fötter och tagit på sig överklädnaden och åter lagt sig ned vid bordet, sade han till dem: »Förstån I vad jag har gjort med eder?
I kallen mig 'Mästare' och 'Herre', och I säger rätt, ty jag är så.
Har nu jag, eder Herre och Mästare, tvagit edra fötter, så ären ock I pliktiga att två varandras fötter.
Jag har ju givit eder ett föredöme, för att I skolen göra såsom jag har gjort mot eder.
Sannerligen, sannerligen säger jag eder: Tjänaren är icke förmer än sin herre, ej heller sändebudet förmer än den som har sänt honom.
Då I veten detta, saliga ären I, om I ock gören det.
Jag talar icke om eder alla; jag vet vilka jag har utvalt.
Men detta skriftens ord skulle ju fullbordas: 'Den som åt mitt bröd, han lyfte mot mig sin häl.'
Redan nu, förrän det sker, säger jag eder det, för att I, när det har skett, skolen tro att jag är den jag är.
Sannerligen, sannerligen säger jag eder: Den som tager emot den jag sänder, han tager emot mig; och den som tager emot mig, han tager emot honom som har sänt mig.»
När Jesus hade sagt detta, blev han upprörd i sin ande och betygade och sade: »Sannerligen, sannerligen säger jag eder: En av eder skall förråda mig.»
Då sågo lärjungarna på varandra och undrade vilken han talade om.
Nu var där bland lärjungarna en som låg till bords invid Jesu bröst, den lärjunge som Jesus älskade.
Åt denne gav då Simon Petrus ett tecken och sade till honom: »Säg vilken det är som han talar om.»
Han lutade sig då mot Jesu bröst och frågade honom: »Herre, vilken är det?»
Då svarade Jesus: »Det är den åt vilken jag räcker brödstycket som jag nu doppar.»
Därvid doppade han brödstycket och räckte det åt Judas, Simon Iskariots son.
Då, när denne hade tagit emot brödstycket, for Satan in i honom.
Och Jesus sade till honom: »Gör snart vad du gör.»
Men ingen av dem som lågo där till bords förstod varför han sade detta till honom.
Ty eftersom Judas hade penningpungen om hand, menade några att Jesus hade velat säga till honom: »Köp vad vi behöva till högtiden», eller ock att han hade tillsagt honom att giva något åt de fattiga.
Då han nu hade tagit emot brödstycket, gick han strax ut; och det var natt.
Och när han hade gått ut, sade Jesus: »Nu är Människosonen förhärligad, och Gud är förhärligad i honom.
Är nu Gud förhärligad i honom, så skall ock Gud förhärliga honom i sig själv, och han skall snart förhärliga honom.
Kära barn, allenast en liten tid är jag ännu hos eder; I skolen sedan söka efter mig, men det som jag sade till judarna: 'Dit jag går, dit kunnen I icke komma', detsamma säger jag nu ock till eder.
Ett nytt bud giver jag eder, att I skolen älska varandra; ja, såsom jag har älskat eder, så skolen ock I älska varandra.
Om I haven kärlek inbördes, så skola alla därav förstå att I ären mina lärjungar.»
Då frågade Simon Petrus honom: »Herre, vart går du?»
Jesus svarade: »Dit jag går, dit kan du icke nu följa mig; men framdeles skall du följa mig.»
Petrus sade till honom: »Herre, varför kan jag icke följa dig nu?
Mitt liv vill jag giva för dig.»
Jesus svarade: »Ditt liv vill du giva för mig?
Sannerligen, sannerligen säger jag dig: Hanen skall icke gala, förrän du tre gånger har förnekat mig.»
»Edra hjärtan vare icke oroliga.
Tron på Gud; tron ock på mig.
I min Faders hus äro många boningar; om så icke voro, skulle jag nu säga eder att jag går bort för att bereda eder rum.
Och om jag än går bort för att bereda eder rum, så skall jag dock komma igen och taga eder till mig; ty jag vill att där jag är, där skolen I ock vara.
Och vägen som leder dit jag går, den veten I.»
Tomas sade till honom: »Herre, vi veta icke vart du går; huru kunna vi då veta vägen?»
Jesus svarade honom: »Jag är vägen och sanningen och livet; ingen kommer till Fadern utom genom mig.
Haden I känt mig, så haden I ock känt min Fader; nu kännen I honom och haven sett honom.»
Filippus sade till honom: »Herre, låt oss se Fadern, så hava vi nog.»
Jesus svarade honom: »Så lång tid har jag varit hos eder, och du har icke lärt känna mig, Filippus?
Den som har sett mig, han har sett Fadern.
Huru kan du då säga: 'Låt oss se Fadern'?
Tror du icke att jag är i Fadern, och att Fadern är i mig?
De ord jag talar till eder talar jag icke av mig själv.
Och gärningarna, dem gör Fadern, som bor i mig; de äro hans verk.
Tron mig; jag är i Fadern, och Fadern i mig.
Varom icke, så tron för själva gärningarnas skull.
Sannerligen, sannerligen säger jag eder: Den som tror på mig, han skall ock själv göra de gärningar som jag gör; och ännu större än dessa skall han göra.
Ty jag går till Fadern,
och vadhelst I bedjen om i mitt namn, det skall jag göra, på det att Fadern må bliva förhärligad i Sonen.
Ja, om I bedjen om något i mitt namn, så skall jag göra det.
Älsken I mig, så hållen I mina bud,
och jag skall bedja Fadern, och han skall giva eder en annan Hjälpare, som för alltid skall vara hos eder:
sanningens Ande, som världen icke kan taga emot, ty hon ser honom icke och känner honom icke.
Men I kännen honom, ty han bor hos eder och skall vara i eder.
Jag skall icke lämna eder faderlösa; jag skall komma till eder.
Ännu en liten tid, och världen ser mig icke mer, men I sen mig.
Ty jag lever; I skolen ock leva.
På den dagen skolen I förstå att jag är i min Fader, och att I ären i mig, och att jag är i eder.
Den som har mina bud och håller dem, han är den som älskar mig; och den som älskar mig, han skall bliva älskad av min Fader, och jag skall älska honom och jag skall uppenbara mig för honom.»
Judas -- icke han som kallades Iskariot -- sade då till honom: »Herre, varav kommer det att du tänker uppenbara dig för oss, men icke för världen?»
Jesus svarade och sade till honom: »Om någon älskar mig, så håller han mitt ord; och min Fader skall älska honom, och vi skola komma till honom och taga vår boning hos honom.
Den som icke älskar mig, han håller icke mina ord; och likväl är det ord som I hören icke mitt, utan Faderns, som har sänt mig.
Detta har jag talat till eder, medan jag ännu är kvar hos eder.
Men Hjälparen, den helige Ande, som Fadern skall sända i mitt namn, han skall lära eder allt och påminna eder om allt vad jag har sagt eder.
Frid lämnar jag efter mig åt eder, min frid giver jag eder; icke giver jag eder den såsom världen giver.
Edra hjärtan vare icke oroliga eller försagda.
I hörden att jag sade till eder: 'Jag går bort, men jag kommer åter till eder.'
Om I älskaden mig, så skullen I ju glädjas över att jag går bort till Fadern, ty Fadern är större än jag.
Och nu har jag sagt eder det, förrän det sker, på det att I mån tro, när det har skett.
Härefter talar jag icke mycket med eder, ty denna världens furste kommer.
I mig finnes intet som hör honom till;
men detta sker, för att världen skall förstå att jag älskar Fadern och gör såsom Fadern har bjudit mig.
Stån upp, låt oss gå härifrån.»
»Jag är det sanna vinträdet, och min Fader är vingårdsmannen.
Var gren i mig, som icke bär frukt, den tager han bort; och var och en som bär frukt, den rensar han, för att den skall bära mer frukt.
I ären redan nu rena, i kraft av det ord som jag har talat till eder.
Förbliven i mig, så förbliver ock jag i eder.
Såsom grenen icke kan bära frukt av sig själv, utan allenast om den förbliver i vinträdet, så kunnen I det ej heller, om I icke förbliven i mig.
Jag är vinträdet, I ären grenarna.
Om någon förbliver i mig, och jag i honom, så bär han mycken frukt; ty mig förutan kunnen I intet göra.
Om någon icke förbliver i mig, så kastas han ut såsom en avbruten gren och förtorkas; och man samlar tillhopa sådana grenar och kastar dem i elden, och de brännas upp.
Om I förbliven i mig, och mina ord förbliva i eder, så mån I bedja om vadhelst I viljen, och det skall vederfaras eder.
Därigenom bliver min Fader förhärligad, att i bären mycken frukt och bliven mina lärjungar.
Såsom Fadern har älskat mig, så har ock jag älskat eder; förbliven i min kärlek.
Om I hållen mina bud, så förbliven I i min kärlek, likasom jag har hållit min Faders bud och förbliver i hans kärlek.
Detta har jag talat till eder, för att min glädje skall bo i eder, och för att eder glädje skall bliva fullkomlig.
Detta är mitt bud, att I skolen älska varandra, såsom jag har älskat eder.
Ingen har större kärlek, än att han giver sitt liv för sina vänner.
I ären mina vänner, om I gören vad jag bjuder eder.
Jag kallar eder nu icke längre tjänare, ty tjänaren får icke veta vad hans herre gör; vänner kallar jag eder, ty allt vad jag har hört av min Fader har jag kungjort för eder.
I haven icke utvalt mig, utan jag har utvalt eder; och jag har bestämt om eder att I skolen gå åstad och bära frukt, sådan frukt som bliver beståndande, på det att Fadern må giva eder vadhelst I bedjen honom om i mitt namn.
Ja, det bjuder jag eder, att I skolen älska varandra.
Om världen hatar eder, så betänken att hon har hatat mig förr än eder.
Voren I av världen, så älskade ju världen vad henne tillhörde; men eftersom I icke ären av världen, utan av mig haven blivit utvalda och tagna ut ur världen, därför hatar världen eder.
Kommen ihåg det ord som jag sade till eder: 'Tjänaren är icke förmer än sin herre.'
Hava de förföljt mig, så skola de ock förfölja eder; hava de hållit mitt ord, så skola de ock hålla edert.
Men allt detta skola de göra mot eder för mitt namns skull, eftersom de icke känna honom som har sänt mig.
Hade jag icke kommit och talat till dem, så skulle de icke hava haft synd; men nu hava de ingen ursäkt för sin synd.
Den som hatar mig, han hatar ock min Fader.
Hade jag icke bland dem gjort sådana gärningar, som ingen annan har gjort, så skulle de icke hava haft synd; men nu hava de sett dem, och hava likväl hatat både mig och min Fader.
Men det ordet skulle ju fullbordas, som är skrivet i deras lag: 'De hava hatat mig utan sak.'
Dock, när Hjälparen kommer, som jag skall sända eder ifrån Fadern, sanningens Ande, som utgår ifrån Fadern, då skall han vittna om mig.
Också I kunnen vittna, eftersom I haven varit med mig från begynnelsen.»
»Detta har jag talat till eder, för att I icke skolen komma på fall.
Man skall utstöta eder ur synagogorna; ja, den tid kommer, då vemhelst som dräper eder skall mena sig därmed förrätta offertjänst åt Gud.
Och så skola de göra, därför att de icke hava lärt känna Fadern, ej heller mig.
Men detta har jag talat till eder, för att I, när den tiden är inne, skolen komma ihåg att jag har sagt eder det.
Jag sade eder det icke från begynnelsen, ty jag var ju hos eder.
Och nu går jag bort till honom som har sänt mig; och ingen av eder frågar mig vart jag går.
Men edra hjärtan äro uppfyllda av bedrövelse, därför att jag har sagt eder detta.
Dock säger jag eder sanningen: Det är nyttigt för eder att jag går bort, ty om jag icke ginge bort, så komme icke Hjälparen till eder; men då jag nu går bort, skall jag sända honom till eder.
Och när han kommer, skall han låta världen få veta sanningen i fråga om synd och rättfärdighet och dom:
i fråga om synd, ty de tro icke på mig;
i fråga om rättfärdighet, ty jag går till Fadern, och I sen mig icke mer;
i fråga om dom, ty denna världens furste är nu dömd.
Jag hade ännu mycket att säga eder, men I kunnen icke nu bära det.
Men när han kommer, som är sanningens Ande, då skall han leda eder fram till hela sanningen.
Ty han skall icke tala av sig själv, utan vad han hör, allt det skall han tala; och han skall förkunna för eder vad komma skall.
Han skall förhärliga mig, ty av mitt skall han taga och skall förkunna det för eder.
Allt vad Fadern har, det är mitt; därför sade jag att han skall taga av mitt och förkunna det för eder.
En liten tid, och I sen mig icke mer; och åter en liten tid, och I fån se mig.»
Då sade några av hans lärjungar till varandra: »Vad är detta som han säger till oss: 'En liten tid, och I sen mig icke; och åter en liten tid, och I fån se mig', så ock: 'Jag går till Fadern'?»
De sade alltså: »Vad är detta som han säger: 'En liten tid'?
Vi förstå icke vad han talar.»
Då märkte Jesus att de ville fråga honom, och han sade till dem: »I talen med varandra om detta som jag sade: 'En liten tid, och I sen mig icke; och åter en liten tid, och I fån se mig.'
Sannerligen, sannerligen säger jag eder: I skolen bliva bedrövade, men eder bedrövelse skall vändas i glädje.
När en kvinna föder barn, har hon bedrövelse, ty hennes stund är kommen; men när hon har fött barnet, kommer hon icke mer ihåg sin vedermöda, ty hon gläder sig över att en människa är född till världen.
Så haven ock I nu bedrövelse; men jag skall se eder åter, och då skola edra hjärtan glädja sig, och ingen skall taga eder glädje ifrån eder.
Och på den dagen skolen I icke fråga mig om något.
Sannerligen, sannerligen säger jag eder: Vad I bedjen Fadern om, det skall han giva eder i mitt namn.
Hittills haven I icke bett om något i mitt namn; bedjen, och I skolen få, för att eder glädje skall bliva fullkomlig.
Detta har jag talat till eder i förtäckta ord; den tid kommer, då jag icke mer skall tala till eder i förtäckta ord, utan öppet förkunna för eder om Fadern.
På den dagen skolen I bedja i mitt namn.
Och jag säger eder icke att jag skall bedja Fadern för eder,
ty Fadern själv älskar eder, eftersom I haven älskat mig och haven trott att jag är utgången från Gud.
Ja, jag har gått ut ifrån Fadern och har kommit i världen; åter lämnar jag världen och går till Fadern.»
Då sade hans lärjungar: »Se, nu talar du öppet och brukar inga förtäckta ord.
Nu veta vi att du vet allt, och att det icke är behövligt för dig att man frågar dig; därför tro vi att du är utgången från Gud.»
Jesus svarade dem: »Nu tron I?
Se, den stund kommer, ja, den är redan kommen, så I skolen förskingras, var och en åt sitt håll, och lämna mig allena.
Dock, jag är icke allena, ty Fadern är med mig.
Detta har jag talat till eder, för att I skolen hava frid i mig.
I världen liden i betryck; men varen vid gott mod, jag har övervunnit världen.»
Sedan Jesus hade talat detta, lyfte han upp sina ögon mot himmelen och sade: »Fader, stunden är kommen; förhärliga din Son, på det att din Son må förhärliga dig,
eftersom du har givit honom makt över allt kött, för att han skall giva evigt liv åt alla dem som du har givit åt honom.
Och detta är evigt liv, att de känna dig, den enda sanne Guden, och den du har sänt, Jesus Kristus.
Jag har förhärligat dig på jorden, genom att fullborda det verk som du har givit mig att utföra.
Och nu, Fader, förhärliga du mig hos dig själv, med den härlighet som jag hade hos dig, förrän världen var till.
Jag har uppenbarat ditt namn för de människor som du har tagit ut ur världen och givit åt mig.
De voro dina, och du har givit dem åt mig, och de hava hållit ditt ord.
Nu hava de förstått att allt vad du har givit åt mig, det kommer från dig.
Ty de ord som du har givit åt mig har jag givit åt dem: och de hava tagit emot dem och hava i sanning förstått att jag är utgången från dig, och de tro att du har sänt mig.
Jag beder för dem; det är icke för världen jag beder, utan för dem som du har givit åt mig, ty de äro dina
-- såsom allt mitt är ditt, och ditt är mitt -- och jag är förhärligad i dem.
Jag är nu icke längre kvar i världen, men de äro kvar i världen, när jag går till dig.
Helige Fader, bevara dem i ditt namn -- det som du har förtrott åt mig -- för att de må vara ett, likasom vi äro ett.
Medan jag var hos dem, bevarade jag dem i ditt namn, det som du har förtrott åt mig; jag vakade över dem, och ingen av dem gick i fördärvet, ingen utom fördärvets man, ty skriften skulle ju fullbordas.
Nu går jag till tid; dock talar jag detta, medan jag ännu är här i världen, för att de skola hava min glädje fullkomlig i sig.
Jag har givit dem ditt ord; och världen har hatat dem, eftersom de icke äro av världen, likasom icke heller jag är av världen.
Jag beder icke att du skall taga dem bort ur världen, utan att du skall bevara dem från det onda.
De äro icke av världen, likasom icke heller jag är av världen.
Helga dem i sanningen; ditt ord är sanning.
Såsom du har sänt mig i världen, så har ock jag sänt dem i världen.
Och jag helgar mig till ett offer för dem, på det att ock de må vara i sanning helgade.
Men icke för dessa allenast beder jag, utan ock för dem som genom deras ord komma till tro på mig;
jag beder att de alla må vara ett, och att, såsom du, Fader, är i mig, och jag i dig, också de må vara i oss, för att världen skall tro att du har sänt mig.
Och den härlighet som du har givit mig, den har jag givit åt dem, för att de skola vara ett, såsom vi äro ett
-- jag i dem, och du i mig -- ja, för att de skola vara fullkomligt förenade till ett, så att världen kan förstå att du har sänt mig, och att du har älskat dem, såsom du har älskat mig.
Fader, jag vill att där jag är, där skola ock de som du har givit mig vara med mig, så att de få se min härlighet, som du har givit mig; ty du har älskat mig före världens begynnelse.
Rättfärdige Fader, världen har icke lärt känna dig, men jag känner dig, och dessa hava förstått att du har sänt mig.
Och jag har kungjort för dem ditt namn och skall kungöra det, på det att den kärlek, som du har älskat mig med, må vara i dem, och jag i dem.»
När Jesus hade sagt detta, begav han sig med sina lärjungar därifrån och gick över bäcken Kidron till andra sidan.
Där var en örtagård, och i den gick han in med sina lärjungar.
Men också Judas, han som förrådde honom, kände till det stället, ty där hade Jesus och hans lärjungar ofta kommit tillsammans.
Och Judas tog nu med sig den romerska vakten, så ock några av översteprästernas och fariséernas tjänare, och kom dit med bloss och lyktor och vapen.
Och Jesus, som visste allt vad som skulle övergå honom, gick fram och sade till dem: »Vem söken I?»
De svarade honom: »Jesus från Nasaret.»
Jesus sade till dem: »Det är jag.»
Och Judas, förrädaren, stod också där ibland dem.
När Jesus nu sade till dem: »Det är jag», veko de tillbaka och föllo till marken.
Åter frågade han dem då: »Vem söken I?»
De svarade: »Jesus från Nasaret.»
Jesus sade: »Jag har sagt eder att det är jag; om det alltså är mig I söken, så låten dessa gå.»
Ty det ordet skulle fullbordas, som han hade sagt: »Av dem som du har givit mig har jag icke förlorat någon.»
Och Simon Petrus, som hade ett svärd, drog ut det och högg till översteprästens tjänare och högg så av honom högra örat; och tjänarens namn var Malkus.
Då sade Jesus till Petrus: »Stick ditt svärd i skidan.
Skulle jag icke dricka den kalk som min Fader har givit mig?»
Den romerska vakten med sin överste och de judiska rättstjänarna grepo då Jesus och bundo honom
och förde honom bort, först till Hannas; denne var nämligen svärfader till Kaifas, som var överstepräst det året.
Och det var Kaifas som under rådplägningen hade sagt till judarna, att det vore bäst om en man finge dö för folket.
Och Simon Petrus jämte en annan lärjunge följde efter Jesus.
Den lärjungen var bekant med översteprästen och gick med Jesus in på översteprästens gård;
men Petrus stod utanför vid porten.
Den andre lärjungen, den som var bekant med översteprästen, gick då ut och talade med portvakterskan och fick så föra Petrus ditin.
Tjänstekvinnan som vaktade porten sade därvid till Petrus: »Är icke också du en av den mannens lärjungar?»
Han svarade: »Nej, det är jag icke.»
Men tjänarna och rättsbetjänterna hade gjort upp en koleld, ty det var kallt, och de stodo där och värmde sig; bland dem stod också Petrus och värmde sig.
Översteprästen frågade nu Jesus om hans lärjungar och om hans lära.
Jesus svarade honom: »Jag har öppet talat för världen, jag har alltid undervisat i synagogan eller i helgedomen, på ställen där alla judar komma tillsammans; hemligen har jag intet talat.
Varför frågar du då mig?
Dem som hava hört mig må du fråga om vad jag har talat till dem.
De veta ju vad jag har sagt.»
När Jesus sade detta, gav honom en av rättstjänarna, som stod där bredvid, ett slag på kinden och sade: »Skall du så svara översteprästen?»
Jesus svarade honom: »Har jag talat orätt, så bevisa att det var orätt; men har jag talat rätt, varför slår du mig då?»
Och Hannas sände honom bunden till översteprästen Kaifas.
Men Simon Petrus stod och värmde sig.
Då sade de till honom: »Är icke också du en av hans lärjungar?»
Han nekade och sade: »Det är jag icke.»
Då sade en av översteprästens tjänare, en frände till den som Petrus hade huggit örat av: »Såg jag icke själv att du var med honom i örtagården?»
Då nekade Petrus åter.
Och i detsamma gol hanen.
Sedan förde de Jesus från Kaifas till pretoriet; och det var nu morgon.
Men själva gingo de icke in i pretoriet, för att de icke skulle bliva orenade, utan skulle kunna äta påskalammet.
Då gick Pilatus ut till dem och sade: »Vad haven I för anklagelse att frambära mot denne man?»
De svarade och sade till honom: »Vore han icke en illgärningsman, så hade vi icke överlämnat honom åt dig.»
Då sade Pilatus till dem: »Tagen I honom, och dömen honom efter eder lag.»
Judarna svarade honom: »För oss är det icke lovligt att avliva någon.»
Ty Jesu ord skulle fullbordas, det som han hade sagt för att giva till känna på vad sätt han skulle dö.
Pilatus gick åter in i pretoriet och kallade Jesus till sig och sade till honom: »Är du judarnas konung?»
Jesus svarade: »Säger du detta av dig själv, eller hava andra sagt dig det om mig?»
Pilatus svarade: »Jag är väl icke en jude!
Ditt eget folk och översteprästerna hava överlämnat dig åt mig.
Vad har du gjort?»
Jesus svarade: »Mitt rike är icke av denna världen.
Om mitt rike vore av denna världen, så hade väl mina tjänare kämpat för att jag icke skulle bliva överlämnad åt judarna.
Men nu är mitt rike icke av denna världen.»
Så sade Pilatus till honom: »Så är du dock en konung?»
Jesus svarade: »Du säger det själv, att jag är en konung.
Ja, därtill är jag född, och därtill har jag kommit i världen, att jag skall vittna för sanningen.
Var och en som är av sanningen, han hör min röst.»
Pilatus sade till honom: »Vad är sanning?»
När han hade sagt detta, gick han åter ut till judarna och sade till dem: »Jag finner honom icke skyldig till något brott.
Nu är det en sedvänja hos eder, att jag vid påsken skall giva eder en fånge lös.
Viljen I då att jag skall giva eder 'judarnas konung' lös?»
Då skriade de åter och sade: »Icke honom, utan Barabbas.»
Men Barabbas var en rövare.
Så tog då Pilatus Jesus och lät gissla honom.
Och krigsmännen vredo samman en krona av törnen och satte den på hans huvud och klädde på honom en purpurfärgad mantel.
Sedan trädde de fram till honom och sade: »Hell dig, du judarnas konung!» och slogo honom på kinden.
Åter gick Pilatus ut och sade till folket: »Se, jag vill föra honom ut till eder, på det att I mån förstå att jag icke finner honom skyldig till något brott.»
Och Jesus kom då ut, klädd i törnekronan och den purpurfärgade manteln.
Och han sade till dem: »Se mannen!»
Då nu översteprästerna och rättstjänarna fingo se honom, skriade de: »Korsfäst!
Korsfäst!»
Pilatus sade till dem: »Tagen I honom, och korsfästen honom; jag finner honom icke skyldig till något brott.»
Judarna svarade honom: »Vi hava själva en lag, och efter den lagen måste han dö, ty han har gjort sig till Guds Son.»
När Pilatus hörde dem tala så, blev hans fruktan ännu större.
Och han gick åter in i pretoriet och frågade Jesus: »Varifrån är du?»
Men Jesus gav honom intet svar.
Då sade Pilatus till honom: »Svarar du mig icke?
Vet du då icke att jag har makt att giva dig lös och makt att korsfästa dig?»
Jesus svarade honom: »Du hade alls ingen makt över mig, om den icke vore dig given ovanifrån.
Därför har den större synd, som har överlämnat mig åt dig.»
Från den stunden sökte Pilatus efter någon utväg att giva honom lös.
Men judarna ropade och sade: »Giver du honom lös, så är du icke kejsarens vän.
Vemhelst som gör sig till konung, han sätter sig upp mot kejsaren.»
När Pilatus hörde de orden, lät han föra ut Jesus och satte sig på domarsätet, på en plats som kallades Litostroton, på hebreiska Gabbata.
Och det var tillredelsedagen före påsken, vid sjätte timmen.
Och han sade till judarna: »Se här är eder konung!»
Då skriade de: »Bort med honom!
Bort med honom!
Korsfäst honom!»
Pilatus sade till dem: »Skall jag korsfästa eder konung?»
Översteprästerna svarade: »Vi hava ingen annan konung än kejsaren.»
Då gjorde han dem till viljes och bjöd att han skulle korsfästas.
Och de togo Jesus med sig.
Och han bar själv sitt kors och kom så ut till det ställe som kallades Huvudskalleplatsen, på hebreiska Golgata.
Där korsfäste de honom, och med honom två andra, en på vardera sidan, och Jesus i mitten.
Men Pilatus lät ock göra en överskrift och sätta upp den på korset; och den lydde så: »Jesus från Nasaret, judarnas konung.»
Den överskriften läste många av judarna, ty det ställe där Jesus var korsfäst låg nära staden: och den var avfattad på hebreiska, på latin och på grekiska.
Då sade judarnas överstepräster till Pilatus: »Skriv icke: 'Judarnas konung', utan skriv att han har sagt sig vara judarnas konung.»
Pilatus svarade: »Vad jag har skrivit, det har jag skrivit.»
Då nu krigsmännen hade korsfäst Jesus, togo de hans kläder och delade dem i fyra delar, en del åt var krigsman.
Också livklädnaden togo de.
Men livklädnaden hade inga sömmar, utan var vävd i ett stycke, uppifrån och alltigenom.
Därför sade de till varandra: »Låt oss icke skära sönder den, utan kasta lott om vilken den skall tillhöra.»
Ty skriftens ord skulle fullbordas: »De delade mina kläder mellan sig och kastade lott om min klädnad.»
Så gjorde nu krigsmännen.
Men vid Jesu kors stodo hans moder och hans moders syster, Maria, Klopas' hustru, och Maria från Magdala.
När Jesus nu fick se sin moder och bredvid henne den lärjunge som han älskade, sade han till sin moder: »Moder, se din son.»
Sedan sade han till lärjungen: »Se din moder.»
Och från den stunden tog lärjungen henne hem till sig.
Eftersom nu Jesus visste att allt annat redan var fullbordat, sade han därefter, då ju skriften skulle i allt uppfyllas: »Jag törstar.»
Där stod då en kärl som var fullt av ättikvin.
Med det vinet fyllde de en svamp, som de satte på en isopsstängel och förde till hans mun.
Och när Jesus hade tagit emot vinet, sade han: »Det är fullbordat.»
Sedan böjde han ned huvudet och gav upp andan.
Men eftersom det var tillredelsedag och judarna icke ville att kropparna skulle bliva kvar på korset över sabbaten (det var nämligen en stor sabbatsdag), bådo de Pilatus att han skulle låta sönderslå de korsfästas ben och taga bort kropparna.
Så kommo då krigsmännen och slogo sönder den förstes ben och sedan den andres som var korsfäst med honom.
När de därefter kommo till Jesus och sågo honom redan vara död, slogo de icke sönder hans ben;
men en av krigsmännen stack upp han sida med ett spjut, och strax kom därifrån ut blod och vatten.
Och den som har sett detta, han har vittnat därom, för att ock I skolen tro; och hans vittnesbörd är sant, och han vet att han talar sanning.
Ty detta skedde, för att skriftens ord skulle fullbordas: »Intet ben skall sönderslås på honom.»
Och åter ett annat skriftens ord lyder så: »De skola se upp till honom som de hava stungit.»
Men Josef från Arimatea, som var en Jesu lärjunge -- fastän i hemlighet, av fruktan för judarna -- kom därefter och bad Pilatus att få taga Jesu kropp; och Pilatus tillstadde honom det.
Då gick han åstad och tog hans kropp.
Och jämväl Nikodemus kom dit, han som första gången hade besökt honom om natten; denne förde med sig en blandning av myrra och aloe, vid pass hundra skålpund.
Och de togo Jesu kropp och omlindade den med linnebindlar och lade dit de välluktande kryddorna, såsom judarna hava för sed vid tillredelse till begravning.
Men invid det ställe där han hade blivit korsfäst var en örtagård, och i örtagården fanns en ny grav, som ännu ingen hade varit lagd i.
Där lade de nu Jesus, eftersom det var judarnas tillredelsedag och graven låg nära.
Men på första veckodagen, medan det ännu var mörkt, kom Maria från Magdala dit till graven och fick se stenen vara borttagen från graven.
Då skyndade hon därifrån och kom till Simon Petrus och till den andre lärjungen, den som Jesus älskade, och sade till dem: »De hava tagit Herren bort ur graven, och vi veta icke var de hava lagt honom.»
Då begåvo sig Petrus och den andre lärjungen åstad på väg till graven.
Och de sprungo båda på samma gång; men den andre lärjungen sprang fortare än Petrus och kom först fram till graven.
Och när han lutade sig ditin, så han linnebindlarna ligga där; dock gick han icke in.
Sedan, efter honom, kom ock Simon Petrus dit.
Han gick in i graven och fick så se huru bindlarna lågo där,
och huru duken som hade varit höljd över hans huvud icke låg tillsammans med bindlarna, utan för sig själv på ett särskilt ställe, hopvecklad.
Då gick ock den andre lärjungen ditin, han som först hade kommit till graven; och han såg och trodde.
De hade nämligen ännu icke förstått skriftens ord, att han skulle uppstå från de döda.
Och lärjungarna gingo så hem till sitt igen.
Men Maria stod och grät utanför graven.
Och under det hon grät, lutade hon sig in i graven
och fick då se två änglar i vita kläder sitta där Jesu kropp hade legat, den ene vid huvudets plats, den andre vid fötternas.
Och de sade till henne: »Kvinna, varför gråter du?»
Hon svarade dem: »De hava tagit bort min Herre, och jag vet icke var de hava lagt honom.»
Vid det hon sade detta, vände hon sig om och fick se Jesus stå där; men hon visste icke att det var Jesus.
Jesus sade till henne: »Kvinna, varför gråter du?
Vem söker du?»
Hon trodde att det var örtagårdsmästaren och svarade honom: »Herre, om det är du som har burit bort honom, så säg mig var du har lagt honom, så att jag kan hämta honom.»
Jesus sade till henne: »Maria!»
Då vände hon sig om och sade till honom på hebreiska: »Rabbuni!» (det betyder mästare).
Jesus sade till henne: »Rör icke vid mig; jag har ju ännu icke farit upp till Fadern.
Men gå till mina bröder, och säg till dem att jag far upp till min Fader och eder Fader, till min Gud och eder Gud.»
Maria från Magdala gick då och omtalade för lärjungarna att hon hade sett Herren, och att han hade sagt detta till henne.
På aftonen samma dag, den första veckodagen, medan lärjungarna av fruktan för judarna voro samlade inom stängda dörrar, kom Jesus och stod mitt ibland dem och sade till dem: »Frid vare med eder!»
Och när han hade sagt detta, visade han dem sina händer och sin sida.
Och lärjungarna blevo glada, när de sågo Herren.
Åter sade Jesus till dem: »Frid vare med eder!
Såsom Fadern har sänt mig, så sänder ock jag eder.»
Och när han hade sagt detta, andades han på dem och sade till dem: »Tagen emot helig ande!
Om I förlåten någon hans synder, så äro de honom förlåtna; och om I binden någon i hans synder, så är han bunden i dem.»
Men Tomas, en av de tolv, han som kallades Didymus, var icke med dem, när Jesus kom.
Då nu de andra lärjungarna sade till honom att de hade sett Herren, svarade han dem: »Om jag icke ser hålen efter spikarna i hans händer och sticker mitt finger i hålen efter spikarna och sticker min hand i hans sida, så kan jag icke tro det.»
Åtta dagar därefter voro hans lärjungar åter därinne, och Tomas var med bland dem.
Då kom Jesus, medan dörrarna voro stängda, och stod mitt ibland de, och sade: »Frid vare med eder!»
Sedan sade han till Tomas: »Räck hit dit finger, se här äro mina händer; och räck hit din hand, och stick den i min sida.
Och tvivla icke, utan tro.»
Tomas svarade och sade till honom: »Min Herre och min Gud!»
Jesus sade till honom: »Eftersom du har sett mig, tror du?
Saliga äro de som icke se och dock tro.»
Ännu många andra tecken, som icke äro uppskrivna i denna bok, gjorde Jesus i sina lärjungars åsyn.
Men dessa hava blivit uppskrivna, för att I skolen tro att Jesus är Messias, Guds Son, och för att I genom tron skolen hava liv i hans namn.
Därefter uppenbarade sig Jesus åter för lärjungarna, vid Tiberias' sjö; och vid den uppenbarelsen gick så till:
Simon Petrus och Tomas, som kallades Didymus, och Natanael, han som var från Kana i Galileen, och Sebedeus' söner voro tillsammans, och med dem två andra av hans lärjungar.
Simon Petrus sade då till dem: »Jag vill gå åstad och fiska.»
De sade till honom: »Vi gå också med dig.»
Så begåvo de sig åstad och stego i båten.
Men den natten fingo de intet.
När det sedan hade blivit morgon, stod Jesus där på stranden; dock visste lärjungarna icke att det var Jesus.
Och Jesus sade till dem: »Mina barn, haven I något att äta?»
De svarade honom: »Nej.»
Han sade till dem: »Kasten ut nätet på högra sidan om båten, så skolen I få.»
Då kastade de ut; och nu fingo de en så stor hop fiskar, att de icke förmådde draga upp nätet.
Den lärjunge som Jesus älskade sade då till Petrus: »Det är Herren.»
När Simon Petrus hörde att det var Herren, tog han på sig sin överklädnad -- ty han var oklädd -- och gav sig i sjön.
Men de andra lärjungarna kommo med båten och drogo efter sig nätet med fiskarna; de voro nämligen icke längre från land än vid pass två hundra alnar.
När de sedan hade stigit i land, sågo de glöd ligga där och fisk, som låg därpå, och bröd.
Jesus sade till dem: »Tagen hit av de fiskar som I nu fingen.»
Då steg Simon Petrus i båten och drog nätet upp på land, och det var fullt av stora fiskar, ett hundra femtiotre stycken.
Och fastän de voro så många, hade nätet icke gått sönder.
Därefter sade Jesus till dem: »Kommen hit och äten.»
Och ingen av lärjungarna dristade sig att fråga honom vem han var, ty de förstodo att det var Herren.
Jesus gick då fram och tog brödet och gav dem, likaledes ock av fiskarna.
Detta var nu tredje gången som Jesus uppenbarade sig för sina lärjungar, sedan han hade uppstått från de döda.
När de hade ätit, sade Jesus till Simon Petrus: »Simon, Johannes' son, älskar du mig mer än dessa göra?»
Han svarade honom: »Ja, Herre; du vet att jag har dig kär.»
Då sade han till honom: »Föd mina lamm.»
Åter frågade han honom, för andra gången: »Simon, Johannes' son, älskar du mig?»
Han svarade honom: »Ja, Herre; du vet att jag har dig kär.»
Då sade han till honom: »Var en herde för mina får.»
För tredje gången frågade han honom: »Simon, Johannes' son, har du mig kär?»
Petrus blev bedrövad över att han för tredje gången frågade honom: »Har du mig kär?»
Och han svarade honom: »Herre, du vet allting; du vet att jag har dig kär.»
Då sade Jesus till honom: »Föd mina får.
Sannerligen, sannerligen säger jag dig: När du var yngre, omgjordade du dig själv och gick vart du ville; men när du bliver gammal, skall du nödgas sträcka ut dina händer, och en annan skall omgjorda dig och föra dig dit du icke vill.»
Detta sade han för att giva till känna med hurudan död Petrus skulle förhärliga Gud.
Och sedan han hade sagt detta, sade han till honom: »Följ mig.»
När Petrus vände sig om, fick han se att den lärjunge som Jesus älskade följde med, densamme som under aftonmåltiden hade lutat sig mot hans bröst och frågat honom: »Herre, vilken är det som skall förråda dig?»
Då nu Petrus såg den lärjungen, frågade han Jesus: »Herre, huru bliver det då med denne?»
Jesus svarade honom: »Om jag vill att han skall leva kvar, till dess jag kommer, vad kommer det dig vid?
Följ du mig.»
Så kom det talet ut ibland bröderna, att den lärjungen icke skulle dö.
Men Jesus hade icke sagt till honom att han icke skulle dö, utan allenast: »Om jag vill att han skall leva kvar, till dess jag kommer, vad kommer det dig vid?»
Det är den lärjungen som vittnar om detta, och som har skrivit detta; och vi veta att hans vittnesbörd är sant.
Ännu mycket annat var det som Jesus gjorde; och om allt detta skulle uppskrivas, det ena med det andra, så tror jag att icke ens hela världen skulle kunna rymma de böcker som då bleve skrivna.
I min förra skrift, gode Teofilus, har jag berättat om allt vad Jesus gjorde och lärde,
ända till den dag då han blev upptagen, sedan han genom helig ande hade givit sina befallningar åt apostlarna som han hade utvalt.
För dem hade han ock genom många säkra bevis tett sig såsom levande, efter utståndet lidande; ty under fyrtio dagar lät han sig ses av dem och talade med dem om Guds rike.
När han då var tillsammans med dem, bjöd han dem och sade: »Lämnen icke Jerusalem, utan förbiden där vad Fadern har utlovat, det varom I haven hört av mig.
Ty Johannes döpte med vatten, men få dagar härefter skolen I bliva döpta i helig ande.»
Då de nu hade kommit tillhopa, frågade de honom och sade: »Herre, skall du nu i denna tid upprätta igen riket åt Israel?»
Han svarade dem: »Det tillkommer icke eder att få veta tider eller stunder som Fadern i sin makt har fastställt.
Men när den helige Ande kommer över eder, skolen I undfå kraft och bliva mina vittnen, både i Jerusalem och i hela Judeen och Samarien, och sedan intill jordens ända.»
När han hade sagt detta, lyftes han inför deras ögon upp i höjden, och en sky tog honom bort ur deras åsyn.
Och medan de skådade mot himmelen, under det han for upp, se, då stodo hos dem två män i vita kläder.
Och dessa sade: »I galileiske män, varför stån I och sen mot himmelen?
Denne Jesus, som har blivit upptagen från eder till himmelen, han skall komma igen på samma sätt som I haven sett honom fara upp till himmelen.»
Sedan vände de tillbaka till Jerusalem från det berg som kallas Oljeberget, vilket ligger nära Jerusalem, icke längre därifrån, än man får färdas på en sabbat.
Och när de hade kommit dit, gingo de upp i den sal i övre våningen, där de plägade vara tillsammans: Petrus och Johannes och Jakob och Andreas, Filippus och Tomas, Bartolomeus och Matteus, Jakob, Alfeus' son, och Simon ivraren och Judas, Jakobs son.
Alla dessa höllo endräktigt ut i bön tillika med Maria, Jesu moder, och några andra kvinnor samt Jesu bröder.
En av de dagarna stod Petrus upp och talade bland bröderna, som då voro församlade till ett antal av omkring etthundratjugu; han sade:
»Mina bröder, det skriftens ord skulle fullbordas, som den helige Ande genom Davids mun hade profetiskt talat om Judas, vilken blev vägvisare åt de män som grepo Jesus.
Han var ju räknad bland oss och hade också fått detta ämbete på sin lott.
Och med de penningar han hade fått såsom lön för sin ogärning förvärvade han sig en åker.
Men han störtade framstupa ned, och hans kropp brast mitt itu, så att alla hans inälvor gåvo sig ut.
Detta blev bekant för alla Jerusalems invånare, och så blev den åkern på deras tungomål kallad Akeldamak (det betyder Blodsåkern).
Så är ju skrivet i Psalmernas bok: 'Hans gård blive öde, och ingen må finnas, som bor däri'; och vidare: 'Hans ämbete tage en annan.'
Därför bör nu någon av de män som följde oss under hela den tid då Herren Jesus gick ut och in bland oss,
allt ifrån den dag då han döptes av Johannes ända till den dag då han blev upptagen och skildes ifrån oss -- någon av dessa män bör insättas till att jämte oss vittna om hans uppståndelse.»
Därefter ställde de fram två: Josef (som kallades Barsabbas och hade tillnamnet Justus) och Mattias.
Och de bådo och sade: »Herre, du som känner allas hjärtan, visa oss vilken av dessa två du har utvalt
till att få den plats såsom tjänare och apostel, vilken Judas övergav, för att gå till den plats som var hans.»
Och de drogo lott om dem, och lotten föll på Mattias.
Och så blev denne, jämte de elva, räknad såsom apostel.
När sedan pingstdagen var inne, voro de alla församlade med varandra.
Då kom plötsligt från himmelen ett dån, såsom om en våldsam storm hade dragit fram; och det uppfyllde hela huset där de sutto.
Och tungor såsom av eld visade sig för dem och fördelade sig och satte sig på dem, en på var av dem.
Och de blevo alla uppfyllda av helig ande och begynte tala andra tungomål, efter som Anden ingav dem att tala.
Nu bodde i Jerusalem fromma judiska män från allahanda folk under himmelen.
Och när dånet hördes, församlade sig hela hopen, och en stor rörelse uppstod, ty var och en hörde sitt eget tungomål talas av dem.
Och de uppfylldes av häpnad och förundran och sade: »Äro de icke galiléer, alla dessa som här tala?
Huru kommer det då till, att var och en av oss hör sitt eget modersmål talas?
Vi må vara parter eller meder eller elamiter, vi må hava vårt hem i Mesopotamien eller Judeen eller Kappadocien, i Pontus eller provinsen Asien,
i Frygien eller Pamfylien, i Egypten eller i Libyens bygder, åt Cyrene till, eller vara hitflyttade främlingar från Rom,
vi må vara judar eller proselyter, kretenser eller araber, alla höra vi dem på våra egna tungomål tala om Guds väldiga gärningar.»
Så uppfylldes de alla av häpnad och visste icke vad de skulle tänka.
Och de sade, den ene till den andre: »Vad kan detta betyda?»
Men somliga drevo gäck med dem och sade: »De äro fulla av sött vin.»
Då trädde Petrus fram, jämte de elva, och hov upp sin röst och talade till dem: »I judiske män och I alla Jerusalems invånare, detta mån I veta, och lyssnen nu till mina ord:
Det är icke så som I menen, att dessa äro druckna; det är ju blott tredje timmen på dagen.
Nej, här uppfylles det som är sagt genom profeten Joel:
'Och det skall ske i de yttersta dagarna, säger Gud, att jag skall utgjuta av min Ande över allt kött, och edra söner och edra döttrar skola profetera, och edra ynglingar skola se syner, och edra gamla män skola hava drömmar;
ja, över mina tjänare och mina tjänarinnor skall jag i de dagarna utgjuta av min Ande, och de skola profetera.
Och jag skall låta undertecken synas uppe på himmelen och tecken nere på jorden: blod och eld och rökmoln.
Solen skall vändas i mörker och månen i blod, förrän Herrens dag kommer, den stora och härliga.
Och det skall ske att var och en som åkallar Herrens namn, han skall varda frälst.'
I män av Israel, hören dessa ord: Jesus från Nasaret, en man som inför eder fick vittnesbörd av Gud genom kraftgärningar och under och tecken, vilka Gud genom honom gjorde bland eder, såsom I själva veten,
denne som blev given i edert våld, enligt vad Gud i sitt rådslut och sin försyn hade bestämt, honom haven I genom män som icke veta av lagen låtit fastnagla vid korset och döda.
Men Gud gjorde en ände på dödens vånda och lät honom uppstå, eftersom det icke var möjligt att han skulle kunna behållas av döden.
Ty David säger med tanke på honom: 'Jag har haft Herren för mina ögon alltid, ja, han är på min högra sida, för att jag icke skall vackla.
Fördenskull gläder sig mitt hjärta, och min tunga fröjdar sig, och jämväl min kropp får vila med en förhoppning:
den, att du icke skall lämna min själ åt dödsriket och icke låta din Helige se förgängelse.
Du har kungjort mig livets vägar; du skall uppfylla mig med glädje inför ditt ansikte.'
Mina bröder, jag kan väl fritt säga till eder om vår stamfader David att han är både död och begraven; hans grav finnes ju ibland oss ännu i dag.
Men eftersom han var en profet och visste att Gud med ed hade lovat honom att 'av hans livs frukt sätta en konung på hans tron',
därför förutsåg han att Messias skulle uppstå, och talade därom och sade att Messias icke skulle lämnas åt dödsriket, och att hans kropp icke skulle se förgängelse.
Denne -- Jesus -- har nu Gud låtit uppstå; därom kunna vi alla vittna.
Och sedan han genom Guds högra hand har blivit upphöjd och av Fadern undfått den utlovade helige Anden, har han utgjutit vad I här sen och hören.
Ty icke har David farit upp till himmelen; fastmer säger han själv: 'Herren sade till min herre: Sätt dig på min högra sida,
till dess jag har lagt dina fiender dig till en fotapall.
Så må nu hela Israels hus veta och vara förvissat om att denne Jesus som I haven korsfäst, honom har Gud gjort både till Herre och till Messias.»
När de hörde detta, kände de ett styng i hjärtat.
Och de sade till Petrus och de andra apostlarna: »Bröder, vad skola vi göra?»
Petrus svarade dem: »Gören bättring, och låten alla döpa eder i Jesu Kristi namn till edra synders förlåtelse; då skolen I såsom gåva undfå den helige Ande.
Ty eder gäller löftet och edra barn, jämväl alla dem som äro i fjärran, så många som Herren, vår Gud, kallar.»
Också med många andra ord bad och förmanade han dem, i det han sade: »Låten frälsa eder från detta vrånga släkte.»
De som då togo emot hans ort läto döpa sig; och så ökades församlingen på den dagen med vid pass tre tusen personer.
Och dessa höllo fast vid apostlarnas undervisning och brödragemenskapen, vid brödsbrytelsen och bönerna.
Och fruktan kom över var och en; och många under och tecken gjordes genom apostlarna.
Men alla de som trodde höllo sig tillsammans och hade allting gemensamt;
de sålde sina jordagods och vad de eljest ägde och delade med sig därav åt alla, eftersom var och en behövde.
Och ständigt, var dag, voro de endräktigt tillsammans i helgedomen; och hemma i husen bröto de bröd och åto med fröjd och i hjärtats enfald, och lovade Gud.
Och allt folket vad dem väl bevåget.
Och Herren ökade församlingen, dag efter dag, med dem som läto sig frälsas.
Och Petrus och Johannes gingo upp till helgedomen, till den bön som hölls vid nionde timmen.
Och där bars fram en man som hade varit ofärdig allt ifrån moderlivet, och som man var dag plägade sätta vid den port i helgedomen, som kallades Sköna porten, för att han skulle kunna begära allmosor av dem som gingo in i helgedomen.
När denne nu fick se Petrus och Johannes, då de skulle gå in i helgedomen, bad han dem om en allmosa.
Då fäste Petrus och Johannes sina ögon på honom, och Petrus sade: »Se på oss.»
När han då gav akt på dem, i förväntan att få något av dem,
sade Petrus: »Silver och guld har jag icke; men vad jag har, det giver jag dig.
I Jesu Kristi, nasaréens namn: stå upp och gå.»
Och så fattade han honom vid högra handen och reste upp honom.
Och strax fingo hans fötter och fotleder styrka,
och han sprang upp och stod upprätt och begynte gå och följde dem in i helgedomen, alltjämt gående och springande, under det att han lovade Gud.
Och allt folket såg honom, där han gick omkring och lovade Gud.
Och när de kände igen honom och sågo att det var samme man som plägade sitta och begära allmosor vid Sköna porten i helgedomen, blevo de uppfyllda av häpnad och bestörtning över det som hade vederfarits honom.
Då han nu höll sig till Petrus och Johannes, strömmade allt folket, utom sig av häpnad, tillsammans till dem på den plats som kallades Salomos pelargång.
När Petrus såg detta, tog han till orda och talade till folket så: »I män av Israel, varför undren I över denne man, och varför sen I så på oss, likasom hade vi genom någon vår kraft eller fromhet åstadkommit att han kan gå?
Nej, Abrahams och Isaks och Jakobs Gud, våra fäders Gud, har förhärligat sin tjänare Jesus, honom som I utlämnaden, och som I förnekaden inför Pilatus, när denne redan hade beslutit att giva honom lös.
Ja, I förnekaden honom, den helige och rättfärdige, och begärden att en dråpare skulle givas åt eder.
Och livets furste dräpten I, men Gud uppväckte honom från de döda; därom kunna vi själva vittna.
Och det är på grund av tron på hans namn som denne man, vilken I sen och kännen, har undfått styrka av hans namn; och den tro som verkas genom Jesus har, i allas eder åsyn, gjort att han nu kan bruka alla lemmar.
Nu vet jag väl, mina bröder, att I såväl som edra rådsherrar haven gjort detta, därför att I icke vissten bättre.
Men Gud har på detta sätt låtit det gå i fullbordan, som han förut genom alla sina profeters mun hade förkunnat, nämligen att hans Smorde skulle lida.
Gören därför bättring och omvänden eder, så att edra synder bliva utplånade,
på det att tider av vederkvickelse må komma från Herren, i det att han sänder den Messias som han har utsett åt eder, nämligen Jesus,
vilken dock himmelen måste behålla intill de tider nå allt skall bliva upprättat igen, varom Gud har talat genom sina forntida heliga profeters mun.
Moses har ju sagt: 'En profet skall Herren Gud låta uppstå åt eder, av edra bröder, en som är mig lik; honom skolen I lyssna till i allt vad han talar till eder.
Och det skall ske att var och en som icke lyssnar till den profeten, han skall utrotas ur folket.'
Och sedan hava alla profeterna, både Samuel och de som följde efter honom, så många som hava talat, också bebådat dessa tider.
I ären själva barn av profeterna och delaktiga i det förbund som Gud slöt med edra fäder, när han sade till Abraham: 'Och i din säd skola alla släkter på jorden varda välsignade.'
För eder först och främst har Gud låtit sin tjänare uppstå, och han har sänt honom för att välsigna eder, när I, en och var, omvänden eder från eder ondska.»
Medan de ännu talade till folket, kommo prästerna och tempelvaktens befälhavare och sadducéerna över dem.
Ty det förtröt dem att du undervisade folket och i Jesus förkunnade uppståndelsen från de döda.
Därför grepo de dem nu och satte dem i fängsligt förvar till följande dag, eftersom det redan var afton.
Men många av dem som hade hört vad som hade talats kommo till tro; och antalet av männen uppgick nu till vid pass fem tusen.
Dagen därefter församlade sig deras rådsherrar och äldste och skriftlärde i Jerusalem;
där voro då ock Hannas, översteprästen, och Kaifas och Johannes och Alexander och alla som voro av översteprästerlig släkt.
Och de läto föra fram dem inför sig och frågade dem: »Av vilken makt eller i genom vilket namn haven I gjort detta?»
Då sade Petrus till dem, uppfylld av helig ande: »I folkets rådsherrar och äldste,
eftersom vi i dag underkastas rannsakning för en god gärning mot en sjuk man och tillfrågas varigenom denne har blivit botad,
så mån I veta, I alla och hela Israels folk, att det är genom Jesu Kristi, nasaréens, namn, hans som I haven korsfäst, men som Gud har uppväckt från de döda -- att det är genom det namnet som denne man står inför eder frisk och färdig.
Han är 'den stenen som av byggningsmännen' -- av eder själva -- 'aktades för intet, men som har blivit en hörnsten'.
Och i ingen annan finnes frälsning; ej heller finnes under himmelen något annat namn, bland människor givet, genom vilket vi kunna bliva frälsta.»
När de sågo Petrus och Johannes vara så frimodiga och förnummo att de voro olärda män ur folket, förundrade de sig.
Men så kände de igen dem och påminde sig att de hade varit med Jesus.
Och när de sågo mannen som hade blivit botad stå där bredvid dem, kunde de icke säga något däremot.
De befallde dem alltså att gå ut från rådsförsamlingen.
Sedan överlade de med varandra
och sade: »Vad skola vi göra med dessa män?
Att ett märkligt tecken har blivit gjort av dem, det är ju uppenbart för alla Jerusalems invånare, och vi kunna icke förneka det.
Men för att detta icke ännu mer skall komma ut bland folket, må vi strängeligen förbjuda dem att hädanefter i det namnet tala för någon människa.»
Därefter kallade de in dem och förbjödo dem helt och hållet att tala eller undervisa i Jesu namn.
Men Petrus och Johannes svarade och sade till dem: »Om det är rätt inför Gud att vi hörsamma eder mer är Gud, därom mån I själva döma;
vi för vår del kunna icke underlåta att tala vad vi hava sett och hört.»
Då förbjödo de dem detsamma ännu strängare, men läto dem sedan gå.
Ty eftersom alla prisade Gud för det som hade skett, kunde de, för folkets skull, icke finna någon utväg genom att straffa dem.
Mannen som genom detta tecken hade blivit botad var nämligen över fyrtio år gammal.
När de alltså hade blivit lösgivna, kommo de till sina egna och omtalade för dem allt vad översteprästerna och de äldste hade sagt dem.
Då de hörde detta, ropade de endräktigt till Gud och sade: »Herre, det är du som har gjort himmelen och jorden och havet och allt vad i dem är.
Och du har genom vår fader Davids, din tjänares, mun sagt genom helig ande: 'Varför larmade hedningarna och tänkte folken fåfänglighet?
Jordens konungar trädde fram, och furstarna samlade sig tillhopa mot Herren och hans Smorde.'
Ja, i sanning, de församlade sig i denna stad mot din helige tjänare Jesus, mot honom som du har smort: Herodes och Pontius Pilatus med hedningarna och Israels folkstammar;
de församlade sig till att utföra allt vad din hand och ditt rådslut förut hade bestämt skola ske.
Och nu, Herre, se till deras hotelser, och giv dina tjänare att de med all frimodighet må förkunna ditt ord,
i det att du uträcker din hand till att bota de sjuka, och till att låta tecken och under ske genom din helige tjänare Jesu namn.»
När de hade slutat att bedja, skakades platsen där de voro församlade, och de blevo alla uppfyllda av den helige Ande, och de förkunnade Guds ord med frimodighet.
Och i hela skaran av dem som trodde var ett hjärta och en själ.
Ingen enda kallade något av det han ägde för sitt, utan du hade allting gemensamt.
Och med stor kraft framburo apostlarna vittnesbördet om Herren Jesu uppståndelse; och stor nåd var över dem alla.
Bland dem fanns ingen som led nöd; ty alla som ägde något jordstycke eller något hus sålde detta och buro fram betalningen för det sålda
och lade den för apostlarnas fötter, och man delade ut därav, så att var och en fick efter som han behövde.
Josef, som av apostlarna ock kallades Barnabas (det betyder förmanaren), en levit som var bördig från Cypern,
också han sålde en åker som han ägde och bar fram penningarna och lade dem för apostlarnas fötter.
Men en ung man vid namn Ananias och hans hustru Safira sålde ett jordagods,
och han tog därvid, med sin hustrus vetskap, undan något av betalningen därför; allenast en del bar han fram och lade för apostlarnas fötter.
Då sade Petrus: »Ananias, varför har Satan fått uppfylla ditt hjärta, så att du har velat bedraga den helige Ande och taga undan något av betalningen för jordstycket?
Detta var ju din egendom, medan du hade det kvar; och när det var sålt, voro ju penningarna i din makt.
Huru kunde du få något sådant i sinnet?
Du har ljugit, icke för människor, utan för Gud.»
När Ananias hörde dessa ord, föll han ned och gav upp andan.
Och stor fruktan kom över alla som hörde detta.
Och de yngre männen stodo upp och höljde in honom och buro ut honom och begrovo honom.
Vid pass tre timmar därefter kom hans hustru in, utan att veta om, vad som hade skett.
Petrus sade då till henne: »Säg mig, var det för den summan I sålden jordstycket?»
Hon svarade: »Ja, för den summan.»
Då sade Petrus till henne: »Huru kunden I vilja komma överens om att fresta Herrens Ande?
Se, härutanför dörren höras nu fotstegen av de män som hava begravt din man; och de skola bära ut också dig.»
Och strax föll hon ned vid hans fötter och gav upp andan; och när de unge männen kommo in, funno de henne död.
De buro då ut henne och begrovo henne bredvid hennes man.
Och stor fruktan kom över hela församlingen och över alla andra som hörde detta.
Och genom apostlarna gjordes många tecken och under bland folket; och de höllo sig alla endräktigt tillsammans i Salomos pelargång.
Av de andra dristade sig ingen att närma sig dem, men folket höll dem i ära.
Och ännu flera trodde och slöto sig till Herren, hela skaror av både män och kvinnor.
Ja, man bar de sjuka ut på gatorna och lade dem på bårar och i sängar, för att, när Petrus kom gående, åtminstone hans skugga måtte falla på någon av dem.
Och jämväl från städerna runt omkring Jerusalem kom folket i skaror och förde med sig sjuka och sådana som voro plågade av orena andar; och alla blevo botade.
Då stod översteprästen upp och alla som höllo med honom -- de som hörde till sadducéernas parti -- och de uppfylldes av nitälskan
och läto gripa apostlarna och sätta dem i allmänt häkte.
Men en Herrens ängel öppnade om natten fängelsets portar och förde ut dem och sade:
»Gån åstad och träden upp i helgedomen, och talen till folket alla det sanna livets ord.»
När de hade hört detta, gingo de inemot dagbräckningen in i helgedomen och undervisade.
Emellertid kommo översteprästen och de som höllo med honom och sammankallade Stora rådet, alla Israels barns äldste.
Därefter sände de åstad till fängelset för att hämta dem.
Men när rättstjänarna kommo dit, funno de dem icke i fängelset.
De vände då tillbaka och omtalade detta
och sade: »Fängelset funno vi stängt med all omsorg och väktarna stående utanför portarna, men då vi öppnade, funno vi ingen därinne.»
När tempelvaktens befälhavare och översteprästerna hörde detta, visst de icke vad de skulle tänka därom, eller vad som skulle bliva av detta.
Då kom någon och berättade för den: »De män som I haven insatt i fängelset, de stå nu i helgedomen och undervisa folket.»
Befälhavaren gick då med rättstjänarna åstad och hämtade dem; dock brukade de icke våld, ty de fruktade att bliva stenade av folket.
Och sedan de hade hämtat dem, förde de dem fram inför Stora rådet.
Och översteprästen anställde förhör med dem
och sade: »Vi hava ju allvarligen förbjudit eder att undervisa i det namnet, och likväl haven I uppfyllt Jerusalem med eder undervisning, och I viljen nu låta den mannens blod komma över oss.»
Men Petrus och de andra apostlarna svarade och sade: »Man måste lyda Gud mer än människor.
Våra fäders Gud har uppväckt Jesus, som I haden upphängt på trä och dödat.
Och Gud har med sin högra hand upphöjt honom till en hövding och frälsare, för att åt Israel förläna bättring och syndernas förlåtelse.
Om allt detta kunna vi själva vittna, så ock den helige Ande, vilken Gud har givit åt dem som äro honom lydiga.»
När de hörde detta, blevo de mycket förbittrade och ville döda dem.
Men en farisé, en laglärare vid namn Gamaliel, som var aktad av allt folket, stod då upp i Rådet och tillsade att man för en kort stund skulle föra ut männen.
Sedan sade han till de andra: »I män av Israel, sen eder för vad I tänken göra med dessa män.
För en tid sedan uppträdde ju Teudas och gav sig ut för att något vara, och till honom slöt sig en hop av vid pass fyra hundra män.
Och han blev dödad, och alla som hade trott på honom förskingrades och blevo till intet.
Efter honom uppträdde Judas från Galileen, vid den tid då skattskrivningen pågick; denne förledde en hop folk till avfall, så att de följde honom.
Också han förgicks, och alla som hade trott på honom blevo förskingrade.
Och nu säger jag eder: Befatten eder icke med dessa män, utan låten dem vara; ty skulle detta vara ett rådslag eller ett verk av människor, så kommer det att slås ned;
men är det av Gud, så kunnen I icke slå ned dessa män.
Sen till, att I icke mån befinnas strida mot Gud själv.»
Och de lydde hans råd; de kallade in apostlarna, och sedan de hade låtit gissla dem, förbjödo de dem att tala i Jesu namn och läto dem därefter gå.
Och de gingo ut från rådsförsamlingen, glada över att de hade aktats värdiga att lida smälek för det namnets skull.
Och de upphörde icke att var dag undervisa i helgedomen och hemma i husen och förkunna evangelium om Kristus Jesus.
Vid denna tid, då nu lärjungarnas antal förökades, begynte de grekiska judarna knorra mot de infödda hebréerna över att deras änkor blevo förbisedda vid den dagliga utdelningen.
Då sammankallade de tolv hela lärjungaskaran och sade: »Det är icke tillbörligt att vi försumma Guds ord för att göra tjänst vid borden.
Så utsen nu bland eder, I bröder, sju män som hava gott vittnesbörd om sig och äro fulla av ande och vishet, män som vi kunna sätta till att sköta denna syssla.
Vi skola då helt få ägna oss åt bönen och åt ordets tjänst.»
Det talet behagade hela menigheten.
Och de utvalde Stefanus, en man som var full av tro och helig ande, vidare Filippus och Prokorus och Nikanor och Timon och Parmenas, slutligen Nikolaus, en proselyt från Antiokia.
Dem läto de träda fram för apostlarna, och dessa bådo och lade händerna på dem.
Och Guds ord hade framgång, och lärjungarnas antal förökades mycket i Jerusalem; och en stor hop av prästerna blevo lydiga och trodde.
Och Stefanus var full av nåd och kraft och gjorde stora under och tecken bland folket.
Men av dem som hörde till den synagoga som kallades »De frigivnes och cyrenéernas och alexandrinernas synagoga», så ock av dem som voro från Cilicien och provinsen Asien, stodo några upp för att disputera med Stefanus.
Dock förmådde de icke stå emot den vishet och den ande som här talade.
Då skaffade de några män som föregåvo att de hade hört honom tala hädiska ord mot Moses och mot Gud.
De uppeggade så folket och de äldste och de skriftlärde och överföllo honom och grepo honom och förde honom inför Stora rådet.
Där läto de falska vittnen träda fram, vilka sade: »Denne man upphör icke att tala mot vår heliga plats och mot lagen.
Ty vi hava hört honom säga att Jesus, han från Nasaret, skall bryta ned denna byggnad och förändra de stadgar som Moses har givit oss.»
Då nu alla som sutto i Rådet fäste sina ögon på honom, syntes dem hans ansikte vara såsom en ängels ansikte.
Och översteprästen frågade: »Förhåller detta sig så?»
Då sade han: »Bröder och fäder, hören mig.
Härlighetens Gud uppenbarade sig för vår fader Abraham, medan han ännu var i Mesopotamien, och förrän han bosatte sig i Karran,
och sade till honom: 'Gå ut ur ditt land och från din släkt, och drag till det land som jag skall visa dig.'
Då gick han åstad ut ur kaldéernas land och bosatte sig i Karran.
Sedan, efter han faders död, bjöd Gud honom att flytta därifrån till detta land, där I nu bon.
Han gav honom ingen arvedel däri, icke ens så mycket som en fotsbredd, men lovade att giva det till besittning åt honom och åt hans säd efter honom; detta var på den tid då han ännu icke hade någon son.
Och vad Gud sade var detta, att hans säd skulle leva såsom främlingar i ett land som icke tillhörde dem, och att man skulle göra dem till trälar och förtrycka dem i fyra hundra år.
'Men det folk vars trälar de bliva skall jag döma', sade Gud; 'sedan skola de draga ut och hålla gudstjänst åt mig på denna plats.'
Och han upprättade ett omskärelsens förbund med honom.
Och så födde han Isak och omskar honom på åttonde dagen, och Isak födde Jakob, och Jakob födde våra tolv stamfäder.
Och våra stamfäder avundades Josef och sålde honom till Egypten.
Men Gud var med honom
och frälste honom ur allt hans betryck och lät honom finna nåd och gav honom vishet inför Farao, konungen i Egypten; och denne satte honom till herre över Egypten och över hela sitt hus.
Och hungersnöd kom över hela Egypten och Kanaan med stort betryck, och våra fäder kunde icke få något att äta.
Men när Jakob fick höra att bröd fanns i Egypten, sände han våra fäder åstad dit, en första gång.
Sedan, när de för andra gången kommo dit, blev Josef igenkänd av sina bröder, och Farao fick kunskap och Josefs släkt.
Därefter sände Josef åstad och kallade till sig sin fader Jakob och hela sin släkt, sjuttiofem personer.
Och Jakob for ned till Egypten; och han dog där, han såväl som våra fäder.
Och man förde dem därifrån till Sikem och lade dem i den grav som Abraham för en summa penningar hade köpt av Emmors barn i Sikem.
Och alltefter som tiden nalkades att det löfte skulle uppfyllas, som Gud hade givit Abraham, växte folket till och förökade sig i Egypten,
till dess en ny konung över Egypten uppstod, en som icke visste av Josef.
Denne konung gick listigt till väga mot vårt folk och förtryckte våra fäder och drev dem till att utsätta sina späda barn, för att dessa icke skulle bliva vid liv.
Vid den tiden föddes Moses, och han 'var ett vackert barn' inför Gud.
Under tre månader fostrades han i sin faders hus;
sedan, när han hade blivit utsatt, lät Faraos dotter hämta honom till sig och uppfostra honom såsom sin egen son.
Och Moses blev undervisad i all egyptiernas visdom och var mäktig i ord och gärningar.
Men när han blev fyrtio år gammal, fick han i sinnet att besöka sina bröder, Israels barn.
När han då såg att en av dem led orätt, tog han den misshandlade i försvar och hämnades honom, i det att han slog ihjäl egyptiern.
Nu menade han att hans bröder skulle förstå att Gud genom honom ville bereda dem frälsning; men de förstodo det icke.
Dagen därefter kom han åter fram till dem, där de tvistade, och ville förlika dem och sade: 'I män, I ären ju bröder; varför gören I då varandra orätt?'
Men den som gjorde orätt mot sin landsman stötte bort honom och sade: 'Vem har satt dig till hövding och domare över oss?
Kanske du vill döda mig, såsom du i går dödade egyptiern?'
Vid det talet flydde Moses bort och levde sedan såsom främling i Madiams land och födde där två söner.
Och när fyrtio är äter voro förlidna, uppenbarade sig för honom, i öknen vid berget Sinai, en ängel i en brinnande törnbuske.
När Moses såg detta, förundrade han sig över synen; och då han gick fram för att se vad det var, hördes Herrens röst:
'Jag är dina fäders Gud, Abrahams, Isaks och Jakobs Gud.'
Då greps Moses av bävan och dristade sig icke att se dit.
Och Herren sade till honom: 'Lös dina skor av dina fötter, ty platsen där du står är helig mark.
Jag har nogsamt sett mitt folks betryck i Egypten, och deras suckan har jag hört, och jag har stigit ned för att rädda dem.
Därför må du nu gå åstad; jag vill sända dig till Egypten.
Denne Moses, som de hade förnekat, i det de sade: 'Vem har satt dig till hövding och domare?', honom sände Gud att vara både en hövding och en förlossare, genom ängeln som uppenbarade sig för honom i törnbusken.
Det var han som förde ut dem, och som gjorde under och tecken i Egyptens land och i Röda havet och i öknen, under fyrtio år.
Det var samme Moses som sade till Israels barn: 'En profet skall Gud låta uppstå åt eder, av edra bröder, en som är mig lik.'
Det var och han, som under den tid då menigheten levde i öknen, både var hos ängeln, som talade med honom på berget Sinai, och tillika hos våra fäder; och han undfick levande ord för att giva dem åt eder.
Men våra fäder ville icke bliva honom lydiga, utan stötte bort honom och vände sig med sina hjärtan mot Egypten
och sade till Aron: 'Gör oss gudar, som kunna gå framför oss; ty vi veta icke vad som har vederfarits denne Moses, som förde oss ut ur Egyptens land.'
Och de gjorde i de dagarna en kalv och buro sedan fram offer åt avguden och gladde sig över sina händers verk.
Då vände Gud sig bort och prisgav dem till att dyrka himmelens härskara, såsom det är skrivet i Profeternas bok: 'Framburen I väl åt mig slaktoffer och spisoffer under de fyrtio åren i öknen, I av Israels hus?
Nej, I buren Moloks tält och guden Romfas stjärna, de bilder som I hade gjort för att tillbedja.
Därför skall jag låta eder föras åstad ända bortom Babylon.'
Våra fäder hade vittnesbördets tabernakel i öknen, så inrättat, som han som talade till Moses hade förordnat att denne skulle göra det, efter den mönsterbild som han hade fått se.
Och våra fäder togo det i arv och förde det sedan under Josua hitin, när de togo landet i besittning, efter de folk som Gud fördrev för våra fäder.
Så var det ända till Davids tid.
Denne fann nåd inför Gud och bad att han måtte finna 'ett rum till boning' åt Jakobs Gud.
Men det var Salomo som fick bygga ett hus åt honom.
Dock, den Högste bor icke i hus som äro gjorda med händer, ty det är såsom profeten säger:
'Himmelen är min tron, och jorden är min fotapall; vad för ett hus skullen I då kunna bygga åt mig, säger Herren, och vad för en plats skulle tjäna mig till vilostad?
Min hand har ju gjort allt detta.'
I hårdnackade, med oomskurna hjärtan och öron, I stån alltid emot den helige Ande, I likaväl som edra fäder.
Vilken av profeterna hava icke edra fäder förföljt?
De hava ju dräpt dem som förkunnade att den Rättfärdige skulle komma, han som I själva nu haven förrått och dräpt,
I som fingen lagen eder given genom änglars försorg, men icke haven hållit den.»
När de hörde detta, blevo de mycket förbittrade i sina hjärtan och beto sina tänder samman mot honom.
Men han, full av helig ande, skådade upp mot himmelen och fick se Guds härlighet och såg Jesus stå på Guds högra sida.
Och han sade: »Jag ser himmelen öppen och Människosonen stå på Guds högra sida.»
Då skriade de med hög röst och höllo för sina öron och stormade alla på en gång emot honom
och förde honom ut ur staden och stenade honom.
Och vittnena lade av sina mantlar vid en ung mans fötter, som hette Saulus.
Så stenade de Stefanus, under det att han åkallade och sade: »Herre Jesus, tag emot min ande.»
Och han föll ned på sina knän och ropade med hög röst: »Herre, tillräkna dem icke denna synd.»
Och när han hade sagt detta, avsomnade han.
Och jämväl Saulus hade gillat att man dödade honom.
Några fromma män begrovo dock Stefanus och höllo en stor dödsklagan efter honom.
Saulus åter for våldsamt fram mot församlingen; han gick omkring i husen och drog fram män och kvinnor och lät sätta dem i fängelse.
Men de som hade blivit kringspridda gingo omkring och förkunnade evangelii ord.
Och Filippus kom så ned till huvudstaden i Samarien och predikade Kristus för folket där.
Och när de hörde Filippus och sågo de tecken som han gjorde, aktade de endräktigt på det som han talade.
Ty från många som voro besatta av orena andar foro andarna ut under höga rop, och många lama och ofärdiga blevo botade.
Och det blev stor glädje i den staden.
Nu var där i staden före honom en man vid namn Simon, som hade övat trolldom, så att han hade slagit det samaritiska folket med häpnad, och som sade sig vara något stort.
Till honom höllo sig alla, både små och stora, och sade: »Denne är vad man kallar 'Guds stora kraft.'»
Och de höllo sig till honom, därför att han genom sina trollkonster under ganska lång tid hade slagit dem med häpnad.
Men nu, då de satte tro till Filippus, som förkunnade evangelium om Guds rike och om Jesu Kristi namn, läto de döpa sig, både män och kvinnor.
Ja, Simon själv kom till tro; och sedan han hade blivit döpt, höll han sig ständigt till Filippus.
Och när han såg de stora tecken och kraftgärningar som denne gjorde, betogs han av häpnad.
Då nu apostlarna i Jerusalem fingo höra att Samarien hade tagit emot Guds ord, sände de dit Petrus och Johannes.
Och när dessa kommo ditned, bådo de för dem, att de måtte undfå helig ande;
ty helig ande hade ännu icke fallit på någon av dem, utan de voro allenast döpta i Herren Jesu namn.
De lade då händerna på dem, och de undfingo helig ande.
När då Simon såg att det var genom apostlarnas handpåläggning som Anden blev given, bjöd han dem penningar
och sade: »Given ock mig den makten, så att var och en som jag lägger händerna på undfår helig ande.»
Då sade Petrus till honom: »Må dina penningar med dig själv gå i fördärvet, eftersom du menar att Guds gåva kan köpas för penningar.
Du har ingen del eller lott i det som här är fråga om, ty ditt hjärta är icke rättsinnigt inför Gud.
Gör fördenskull bättring och upphör med denna din ondska, och bed till Herren att den tanke som har uppstått i ditt hjärta må, om möjligt är, bliva dig förlåten.
Ty jag ser att du är förgiftad av ondska och fången i orättfärdighetens bojor.»
Då svarade Simon och sade: »Bedjen I till Herren för mig, att intet av det som I haven sagt må komma över mig.»
Och sedan de hade framburit sitt vittnesbörd och talat Herrens ord, begåvo de sig tillbaka till Jerusalem och förkunnade därvid evangelium i många samaritiska byar.
Men en Herrens ängel talade till Filippus och sade: »Stå upp och begiv dig vid middagstiden ut på den väg som leder ned från Jerusalem till Gasa; den är tom på folk.»
Då stod han upp och begav sig åstad.
Och se, en etiopisk man for där fram, en hovman som var en mäktig herre hos Kandace, drottningen i Etiopien, och var satt över hela hennes skattkammare.
Denne hade kommit till Jerusalem för att där tillbedja,
men var nu stadd på hemvägen och satt i sin vagn och läste profeten Esaias.
Då sade Anden till Filippus: »Gå fram och närma dig till denna vagn.»
Filippus skyndade fram och hörde att han läste profeten Esaias.
Då frågade han: »Förstår du vad du läser?»
Han svarade: »Huru skulle jag väl kunna förstå det, om ingen vägleder mig?»
Och han bad Filippus stiga upp och sätta sig bredvid honom.
Men det ställe i skriften som han läste var detta: »Såsom ett får fördes han bort till att slaktas; och såsom ett lamm som är tyst inför den som klipper det, så öppnade han icke sin mun.
Genom hans förnedring blev hans dom borttagen.
Vem kan räkna hans släkte?
Ty hans liv ryckes undan från jorden.»
Och hovmannen frågade Filippus och sade: »Jag beder dig, säg mig om vilken profeten talar detta, om sig själv eller om någon annan?»
Då öppnade Filippus sin mun och begynte med detta skriftens ord och förkunnade för honom evangelium om Jesus.
Och medan de färdades vägen fram, kommo de till ett vatten.
Då sade hovmannen: »Se, här finnes vatten.
Vad hindrar att jag döpes?»
272810
Och han lät vagnen stanna; och de stego båda ned i vattnet, Filippus och hovmannen, och han döpte honom.
Men när de hade stigit upp ur vattnet, ryckte Herrens Ande bort Filippus, och hovmannen såg honom icke mer, då han nu glad fortsatte sin färd.
Men Filippus blev efteråt sedd i Asdod.
Därefter vandrade han omkring och förkunnade evangelium i alla städer, till dess han kom till Cesarea.
Men Saulus, som alltjämt andades hot och mordlust mot Herrens lärjungar, gick till översteprästen
och utbad sig av honom brev till synagogorna i Damaskus, för att, om han funne några som voro på »den vägen», vare sig män eller kvinnor, han skulle kunna föra dem bundna till Jerusalem.
Men när han på sin färd nalkades Damaskus, hände sig att ett sken från himmelen plötsligt kringstrålade honom.
Och han föll ned till jorden och hörde då en röst som sade till honom: »Saul, Saul, varför förföljer du mig?»
Då sade han: »Vem är du, Herre?»
Han svarade: »Jag är Jesus, den som du förföljer.
Men stå nu upp och gå in i staden, så skall där bliva dig sagt vad du har att göra.»
Och männen som voro med honom på färden stodo mållösa av skräck, ty de hörde väl rösten, men sågo ingen.
Och Saulus reste sig upp från jorden, men när han öppnade sina ögon, kunde han icke mer se något.
De togo honom därför vid handen och ledde honom in i Damaskus.
Och under tre dagar såg han intet; och han varken åt eller drack.
Men i Damaskus fanns en lärjunge vid namn Ananias.
Till honom sade Herren i en syn: »Ananias!»
Han svarade: »Här är jag, Herre.»
Och Herren sade till honom: »Stå upp och gå till den gata som kallas Raka gatan och fråga i Judas' hus efter en man vid namn Saulus, från Tarsus.
Ty se, han beder.
Och i en syn har han sett huru en man vid namn Ananias kom in och lade händerna på honom, för att han skulle få sin syn igen.»
Då svarade Ananias: »Herre, jag har av många hört huru mycket ont den mannen har gjort dina heliga i Jerusalem.
Och han har nu här med sig fullmakt ifrån översteprästerna att fängsla alla dem som åkalla ditt namn.»
Men Herren sade till honom: »Gå åstad; ty denne man är mig ett utvalt redskap till att bära fram mitt namn inför hedningar och konungar och inför Israels barn;
och jag skall visa honom huru mycket han måste lida för mitt namns skull.»
Då gick Ananias åstad och kom in i huset; och han lade sina händer på honom och sade: »Saul, min broder, Herren har sänt mig, Jesus, som visade sig för dig på vägen där du färdades; han har sänt mig, för att du skall få din syn igen och bliva uppfylld av helig ande.»
Då var det strax såsom om fjäll föllo ifrån hans ögon, och han fick sin syn igen.
Och han stod upp och lät döpa sig.
Sedan tog han sig mat och blev därav stärkt.
Därefter var han någon tid tillsammans med lärjungarna i Damaskus.
Och strax begynte han i synagogorna predika om Jesus, att han var Guds Son.
Och alla som hörde honom blevo uppfyllda av häpnad och sade: »Var det icke denne som i Jerusalem förgjorde dem som åkallade det namnet?
Och hade han icke kommit hit, för att han skulle föra sådana människor bundna till översteprästerna?»
Men Saulus uppträdde med allt större kraft och gjorde de judar som bodde i Damaskus svarslösa, i det han bevisade att Jesus var Messias.
När så en längre tid hade förgått, rådslogo judarna om att röja honom ur vägen;
men deras anslag blev bekant för Saulus.
Och då de nu, för att kunna röja honom ur vägen, till och med höllo vakt vid stadsportarna både dag och natt,
togo hans lärjungar honom en natt och släppte honom ut genom muren, i det att de sänkte ned honom i en korg.
När han sedan kom till Jerusalem, försökte han att närma sig lärjungarna; men alla fruktade för honom, ty de trodde icke att han verkligen var en lärjunge.
Då tog Barnabas sig an honom och förde honom till apostlarna och förtäljde för dem huru han på vägen hade sett Herren, som hade talat till honom, och huru han i Damaskus hade frimodigt predikat i Jesu namn.
Sedan gick han fritt ut och in bland dem i Jerusalem och predikade frimodigt i Herrens namn;
och han talade och disputerade med de grekiska judarna.
Men de gjorde försök att röja honom ur vägen.
När bröderna förnummo detta, förde de honom ned till Cesarea och sände honom därifrån vidare till Tarsus.
Så hade nu församlingen frid i hela Judeen och Galileen och Samarien; och den blev uppbyggd och vandrade i Herrens fruktan och växte till genom den helige Andes tröst och förmaning.
Medan nu Petrus vandrade omkring bland dem alla, hände sig att han ock kom ned till de heliga som bodde i Lydda.
Där träffade han på en man vid namn Eneas, som i åtta år hade legat till sängs; han var nämligen lam.
Och Petrus sade till honom: »Eneas, Jesus Kristus botar dig.
Stå upp och lägg ihop din bädd.»
Då stod han strax upp.
Och alla som bodde i Lydda och i Saron sågo honom; och de omvände sig till Herren.
I Joppe bodde då en lärjunginna vid namn Tabita (det betyder detsamma som Dorkas).
Hon överflödade i goda gärningar och gav allmosor rikligen.
Men just i de dagarna hände sig att hon blev sjuk och dog.
Och man tvådde henne och lade henne i en sal i övre våningen.
Då nu Lydda låg nära Joppe och lärjungarna hade hört att Petrus var där, sände de två män till honom och bådo honom att utan dröjsmål komma till dem.
Petrus stod då upp och följde med dem.
Och när han kom dit, förde de honom upp i salen; och alla änkorna kommo där omkring honom gråtande och visade honom alla livklädnader och mantlar som Dorkas hade gjord, medan hon ännu levde ibland dem.
Då tillsade Petrus dem allasammans att gå ut och föll ned på sina knän och bad; sedan vände han sig mot den döda och sade: »Tabita, stå upp.»
Då slog hon upp ögonen, och när hon fick se Petrus, satte hon sig upp.
Och han räckte henne handen och reste upp henne och kallade sedan in de heliga, jämte änkorna, och ställde henne levande framför den.
Detta blev bekant i hela Joppe, och många kommo till tro på Herren.
Därefter stannade han en längre tid i Joppe hos en garvare vid namn Simon.
I Cesarea bodde en man vid namn Kornelius, en hövitsman vid den så kallade italiska krigsskaran.
Han var en from man, som »fruktade Gud» tillika med hela sitt hus; han utdelade rikligen allmosor åt folket och bad alltid till Gud.
En dag omkring nionde timmen såg denne tydligt i en syn en Guds ängel, som kom in till honom och sade till honom: »Kornelius!»
Han betraktade honom förskräckt och frågade: »Vad är det, herre?»
Då sade ängeln till honom: »Dina böner och dina allmosor hava uppstigit till Gud och äro i åminnelse hos honom.
Så sänd nu några män till Joppe och låt hämta en viss Simon, som ock kallas Petrus.
Han gästar hos en garvare vid namn Simon, som har ett hus vid havet.»
När ängeln som hade talat med honom var borta, kallade han till sig två av sina tjänare och en from krigsman, en av dem som hörde till hans närmaste följe,
och förtäljde alltsammans för dem och sände dem åstad till Joppe.
Men dagen därefter, medan dessa voro på vägen och nalkades staden, gick Petrus vid sjätte timmen upp på taket för att bedja.
Och han blev hungrig och ville hava något att äta.
Medan man nu tillredde maten, föll han i hänryckning.
Han såg himmelen öppen och någonting komma ned som liknade en stor linneduk, och som fasthölls vid de fyra hörnen och sänktes ned till jorden.
Och däri funnos alla slags fyrfota och krälande djur som leva på jorden, och alla slags himmelens fåglar.
Och en röst kom till honom: »Stå upp, Petrus, slakta och ät.»
Men Petrus svarade: »Bort det, Herre!
Jag har aldrig ätit något oheligt och orent.»
Åter, för andra gången, kom en röst till honom: »Vad Gud har förklarat för rent, det må du icke hålla för oheligt.»
Detta skedde tre gånger efter varandra; sedan blev duken strax åter upptagen till Himmelen.
Medan Petrus i sitt sinne undrade över vad den syn han hade sett skulle betyda, hade de män som voro utsända av Kornelius redan frågat sig fram till Simons hus; och de stannade nu vid porten
och ropade på någon för att få veta om Simon, som ock kallades Petrus, gästade där.
Men under det Petrus alltjämt begrundade synen, sade Anden till honom: »Här äro ett par män som fråga efter dig.
Stå upp, och gå ditned och följ med dem, utan att tveka; ty det är jag som har sänt dem.»
Då steg Petrus ned till männen och sade: »Se här är jag, den som I frågen efter.
Av vilken orsak haven I kommit hit?»
De svarade: »Hövitsmannen Kornelius, en rättfärdig och gudfruktig man, som har gott vittnesbörd om sig av hela det judiska folket, har i en uppenbarelse fått befallning av en helig ängel att hämta dig till sig och höra vad du har att säga.»
Då bjöd han dem komma in och beredde dem härbärge.
Dagen därefter stod han upp och begav sig åstad med dem; och några av bröderna i Joppe följde med honom.
Följande dag kommo de fram till Cesarea.
Och Kornelius väntade på dem och hade kallat tillhopa sina fränder och närmaste vänner.
Då nu Petrus skulle träda in, gick Kornelius emot honom och betygade honom sin vördnad, i det att han föll ned för hans fötter.
Men Petrus reste upp honom och sade: »Stå upp; också jag är en människa.»
Och under samtal med honom trädde Petrus in och fann många vara där församlade.
Och han sade till dem: »I veten själva att det är en judisk man förbjudet att hava något umgänge med en utlänning eller att besöka en sådan; men mig har Gud lärt att icke räkna någon människa för ohelig eller oren.
Därför kom jag ock utan invändning hit, när jag blev hämtad.
Och nu frågar jag eder av vilket skäl I haven låtit hämta mig.»
Då svarade Kornelius: »Det är nu fjärde dagen sedan jag, just vid denna timme, förrättade i mitt hus den bön som man beder vid nionde timmen.
Då fick jag se en man i skinande klädnad stå framför mig,
och han sade: 'Kornelius, din bön är hörd, och dina allmosor hava kommit i åminnelse inför Gud.
Så sänd nu bud till Joppe och kalla till dig Simon, som ock kallas Petrus: han gästar i garvaren Simons hus vid havet.'
Då sände jag strax bud till dig, och du gjorde väl i att du kom.
Och nu äro vi alla här tillstädes inför Gud för att höra allt som har blivit dig befallt av Herren.»
Då öppnade Petrus sin mun och sade: »Nu förnimmer jag i sanning att 'Gud icke har anseende till personen',
utan att den som fruktar honom och övar rättfärdighet, han tages emot av honom, vilket folk han än må tillhöra.
Det ord som han har sänt till Israels barn för att genom Jesus Kristus, som är allas Herre, förkunna det glada budskapet om frid, det ordet kännen I,
den förkunnelse som gick ut över hela Judeen, sedan den hade begynt i Galileen efter den döpelse Johannes predikade --
förkunnelsen om Jesus från Nasaret och om huru Gud hade smort honom med helig ande och kraft, honom som vandrade omkring och gjorde gott och botade alla som voro under djävulens våld; ty Gud var med honom.
Vi kunna själva vittna om allt vad han gjorde både på den judiska landsbygden och i Jerusalem; likväl upphängde man honom på trä och dödade honom.
Men honom har Gud uppväckt på tredje dagen och låtit honom bliva uppenbar,
väl icke för allt folket, men för oss, som redan förut av Gud hade blivit utvalda till vittnen, och som åto och drucko med honom, sedan han hade uppstått från de döda.
Och han bjöd oss predika för folket och betyga att han är den som av Gud har blivit bestämd till att vara domare över levande och döda.
Om honom bära alla profeterna vittnesbörd och betyga att var och en som tror på honom skall få syndernas förlåtelse genom hans namn.»
Medan Petrus ännu så talade, föll den helige Ande på alla dem som hörde hans tal.
Och alla de omskurna troende män som hade kommit dit med Petrus blevo uppfyllda av häpnad över att den helige Ande hade blivit utgjuten jämväl över hedningarna, såsom en gåva åt dem.
De hörde dem nämligen tala tungomål och storligen prisa Gud.
Då tog Petrus till orda och sade: »Icke kan väl någon hindra att dessa döpas med vatten, då de hava undfått den helige Ande, de likaväl som vi?»
Och så bjöd han att man skulle döpa dem i Jesu Kristi namn.
Därefter bådo de honom att han skulle stanna hos dem några dagar.
Men apostlarna och de bröder som voro i Judeen fingo höra att också hedningarna hade tagit emot Guds ord.
När så Petrus kom upp till Jerusalem, begynte de som voro omskurna gå till rätta med honom;
de sade: »Du har ju besökt oomskurna män och ätit med dem.»
Då begynte Petrus från början och omtalade för dem allt i följd och ordning; han sade:
»Jag var i staden Joppe, stadd i bön; då såg jag under hänryckning i en syn någonting komma ned, som liknade en stor linneduk, vilken fasthölls vid de fyra hörnen och sänktes ned från himmelen; och det kom ända ned till mig.
Och jag betraktade det och gav akt därpå; då fick jag däri se fyrfota djur, sådana som leva på jorden, tama och vilda, så ock krälande djur och himmelens fåglar.
Jag hörde ock en röst säga till mig: 'Stå upp, Petrus, slakta och ät.'
Men jag svarade: 'Bort det, Herre!
Aldrig har något oheligt eller orent kommit i min mun.'
För andra gången talade en röst från himmelen: 'Vad Gud har förklarat för rent, det må du icke hålla för oheligt.'
Detta skedde tre gånger efter varandra; sedan drogs alltsammans åter upp till himmelen.
Och i detsamma kommo tre män, som hade blivit sända till mig från Cesarea, och stannade framför huset där vi voro.
Och Anden sade till mig att jag skulle följa med dem, utan att göra någon åtskillnad mellan folk och folk.
Också de sex bröder som äro här kommo med mig; och vi gingo in i mannens hus.
Och han berättade för oss huru han hade sett ängeln träda in i hans hus, och att denne hade sagt: 'Sänd åstad till Joppe och låt hämta Simon, som ock kallas Petrus.
Han skall tala till dig ord genom vilka du skall bliva frälst, du själv och hela ditt hus.'
Och när jag hade begynt tala, föll den helige Ande på dem, alldeles såsom det under den första tiden skedde med oss.
Då kom jag ihåg Herrens ord, huru han hade sagt: 'Johannes döpte med vatten, men I skolen bliva döpta i helig ande.'
Då alltså Gud åt dem hade givit samma gåva som åt oss, som hava kommit till tro på Herren Jesus Kristus, huru skulle då jag hava kunnat sätta mig emot Gud?»
När de hade hört detta, gåvo de sig till freds och prisade Gud och sade: »Så har då Gud också åt hedningarna förlänat den bättring som för till liv.»
De som hade blivit kringspridda genom den förföljelse som utbröt för Stefanus' skull drogo emellertid omkring ända till Fenicien och Cypern och Antiokia, men förkunnade icke ordet för andra än för judar.
Dock funnos bland dem några män från Cypern och Cyrene, som när de kommo till Antiokia, också talade till grekerna och för dem förkunnade evangelium om Herren Jesus.
Och Herrens hand var med dem, och en stor skara kom till tro och omvände sig till Herren.
Ryktet härom nådde församlingen i Jerusalem; och de sände då Barnabas till Antiokia.
När han kom dit och fick se vad Guds nåd hade verkat, blev han glad och förmanade dem alla att med hjärtats fasta föresats stadigt hålla sig till Herren.
Ty han var en god man och full av helig ande och tro.
Och ganska mycket folk blev ytterligare fört till Herren.
Sedan begav han sig åstad till Tarsus för att uppsöka Saulus.
Och när han hade träffat honom, tog han honom med sig till Antiokia.
Ett helt år hade de sedan sin umgängelse inom församlingen och undervisade ganska mycket folk.
Och det var i Antiokia som lärjungarna först begynte kallas »kristna».
Vid den tiden kommo några profeter från Jerusalem ned till Antiokia.
Och en av dem, vid namn Agabus, trädde upp och gav genom Andens ingivelse till känna att en stor hungersnöd skulle komma över hela världen; den kom också på Klaudius' tid.
Då bestämde lärjungarna att de, var och en efter sin förmåga, skulle sända något till understöd åt de bröder som bodde i Judeen.
Detta gjorde de också, och genom Barnabas och Saulus översände de det till de äldste.
Vid den tiden lät konung Herodes gripa och misshandla några av dem som hörde till församlingen.
Och Jakob, Johannes' broder, lät han avrätta med svärd.
När han såg att detta behagade judarna, fortsatte han och lät fasttaga också Petrus.
Detta skedde under det osyrade brödets högtid.
Och sedan han hade gripit honom, satte han honom i fängelse och uppdrog åt fyra vaktavdelningar krigsmän, vardera på fyra man, att bevaka honom; och hans avsikt var att efter påsken ställa honom fram inför folket.
Under tiden förvarades Petrus i fängelset, men församlingen bad enträget till Gud för honom.
Natten före den dag då Herodes tänkte draga honom inför rätta låg Petrus och sov mellan två krigsmän, fängslad med två kedjor; och utanför dörren voro väktare utsatta till att bevaka fängelset.
Då stod plötsligt en Herrens ängel där, och ett sken lyste i rummet.
Och han stötte Petrus i sidan och väckte honom och sade: »Stå nu strax upp»; och kedjorna föllo ifrån hans händer.
Ängeln sade ytterligare till honom: »Omgjorda dig, och tag på dig dina sandaler.»
Och han gjorde så. därefter sade ängeln till honom: »Tag din mantel på dig och följ mig.»
Och Petrus gick ut och följde honom; men han förstod icke att det som skedde genom ängeln var något verkligt, utan trodde att det var en syn han såg.
När de så hade gått genom första och andra vakten, kommo de till järnporten som ledde ut till staden.
Den öppnade sig för dem av sig själv, och de trädde ut och gingo en gata fram; och i detsamma försvann ängeln ifrån honom.
När sedan Petrus kom till sig igen, sade han: »Nu vet jag och är förvissad om att Herren har utsänt sin ängel och räddat mig ur Herodes' hand och undan allt det som det judiska folket hade väntat sig.»
När han alltså hade förstått huru det var, gick han till det hus där Maria bodde, hon som var moder till den Johannes som ock kallades Markus; där voro ganska många församlade och bådo.
Då han nu klappade på portdörren, kom en tjänsteflicka, vid namn Rode, för att höra vem det var.
Och när hon kände igen Petrus' röst, öppnade hon i sin glädje icke porten, utan skyndade in och berättade att Petrus stod utanför porten.
Då sade de till henne: »Du är från dina sinnen.»
Men hon bedyrade att det var såsom hon hade sagt.
Då sade de: »Det är väl hans ängel.»
Men Petrus fortfor att klappa; och när de öppnade, sågo de med häpnad att det var han.
Och han gav tecken åt dem med handen att de skulle tiga, och förtäljde för dem huru Herren hade fört honom ut ur fängelset.
Och han tillade: »Låten Jakob och de andra bröderna få veta detta.»
Sedan gick han därifrån och begav sig till en annan ort.
Men när det hade blivit dag, uppstod bland krigsmännen en ganska stor oro och undran över vad som hade blivit av Petrus.
När så Herodes ville hämta honom, men icke fann honom, anställde han rannsakning med väktarna och bjöd att de skulle föras bort till bestraffning.
Därefter for han ned från Judeen till Cesarea och vistades sedan där.
Men han hade fattat stor ovilja mot tyrierna och sidonierna.
Dessa infunno sig nu gemensamt hos honom; och sedan de hade fått Blastus, konungens kammarherre, på sin sida, bådo de om fred, ty deras land hade sin näring av konungens.
På utsatt dag klädde sig då Herodes i konungslig skrud och satte sig på tronen och höll ett tal till dem.
Då ropade folket: »En guds röst är detta, och icke en människas.»
Men i detsamma slog honom en Herrens ängel, därför att han icke gav Gud äran.
Och han föll i en sjukdom som bestod däri att han uppfrättes av maskar, och så gav han upp andan.
Men Guds ord hade framgång och utbredde sig.
Och sedan Barnabas och Saulus hade fullgjort sitt uppdrag i Jerusalem och avlämnat understödet, vände de tillbaka och togo då med sig Johannes, som ock kallades Markus.
I den församling som fanns i Antiokia verkade nu såsom profeter och lärare Barnabas och Simeon, som kallades Niger, och Lucius från Cyrene, så ock Manaen, landsfursten Herodes' fosterbroder, och Saulus.
När dessa förrättade Herrens tjänst och fastade, sade den helige Ande: »Avskiljen åt mig Barnabas och Saulus för det verk som jag har kallat dem till.»
Då fastade de och bådo och lade händerna på dem och läto dem begiva sig åstad.
Dessa, som så hade blivit utsända av den helige Ande, foro nu ned till Seleucia och seglade därifrån till Cypern.
Och när de hade kommit till Salamis, förkunnade de Guds ord i judarnas synagogor.
De hade också med sig Johannes såsom tjänare.
Och sedan de hade färdats över hela ön ända till Pafos, träffade de där på en judisk trollkarl och falsk profet, vid namn Barjesus,
som vistades hos landshövdingen Sergius Paulus.
Denne var en förståndig man.
Han kallade till sig Barnabas och Saulus och begärde att få höra Guds ord.
Men Elymas (eller trollkarlen, ty namnet har den betydelsen) stod emot dem och ville hindra landshövdingen från att komma till tro.
Saulus, som ock kallades Paulus, uppfylldes då av helig ande och fäste ögonen på honom
och sade: »O du djävulens barn, du som är full av allt slags svek och arglistighet och en fiende till allt vad rätt är, skall du då icke upphöra att förvrida Herrens raka vägar?
Se, nu kommer Herrens hand över dig, och du skall till en tid bliva blind och icke kunna se solen.»
Och strax föll töcken och mörker över honom; och han gick omkring och sökte efter någon som kunde leda honom.
När då landshövdingen såg vad som hade skett, häpnade han över Herrens lära och kom till tro.
Paulus och hans följeslagare lade sedan ut ifrån Pafos och foro till Perge i Pamfylien.
Där skilde sig Johannes ifrån dem och vände tillbaka till Jerusalem.
Men själva foro de vidare från Perge och kommo till Antiokia i Pisidien.
Och på sabbatsdagen gingo de in i synagogan och satte sig där.
Och sedan man hade föreläst ur lagen och profeterna, sände synagogföreståndarna till dem och läto säga: »Bröder, haven I något förmaningens ord att säga till folket, så sägen det.»
Då stod Paulus upp och gav tecken med handen och sade: »I män av Israels hus och I som 'frukten Gud', hören mig.
Detta folks, Israels, Gud utvalde våra fäder, och han upphöjde detta folk, medan de ännu bodde såsom främlingar i Egyptens land, och förde dem sedan ut därifrån 'med upplyft arm'.
Och under en tid av vid pass fyrtio år hade han fördrag med dem i öknen.
Och sedan han hade utrotat sju folk i Kanaans land, utskiftade han dessas land till arvedelar åt dem.
Därunder förgick en tid av vid pass fyra hundra femtio år.
Sedan gav han dem domare, ända till profeten Samuels tid.
Därefter begärde de en konung; och Gud gav dem Saul, Kis' son, en man av Benjamins stam, för en tid av fyrtio år.
Men denne avsatte han och gjorde David till konung över dem.
Honom gav han ock sitt vittnesbörd, i det han sade: 'Jag har funnit David, Jessais son, en man efter mitt hjärta.
Han skall i alla stycken göra min vilja.'
Av dennes säd har Gud efter sitt löfte låtit Jesus komma, såsom Frälsare åt Israel.
Men redan innan han uppträdde, hade Johannes predikat bättringens döpelse för hela Israels folk.
Och när Johannes höll på att fullborda sitt lopp, sade han: 'Vad I menen mig vara, det är jag icke.
Men se, efter mig kommer den vilkens skor jag icke är värdig att lösa av han fötter.'
Mina bröder, I som ären barn av Abrahams släkt, så ock I andra här, I som 'frukten Gud', till oss har ordet om denna frälsning blivit sänt.
Ty eftersom Jerusalems invånare och deras rådsherrar icke kände honom, uppfyllde de ock genom sin dom över honom profeternas utsagor, vilka var sabbat föreläses;
och fastän de icke funno honom skyldig till något som förtjänade döden, bådo de likväl Pilatus att han skulle låta döda honom.
När de så hade fört till fullbordan allt som var skrivet om honom, togo de honom ned från korsets trä och lade honom i en grav.
Men Gud uppväckte honom från de döda.
Sedan visade han sig under många dagar för dem som med honom hade gått upp från Galileen till Jerusalem, och som nu äro hans vittnen inför folket.
Och vi förkunna för eder det glada budskapet, att det löfte som gavs åt våra fäder, det har Gud låtit gå i fullbordan för oss, deras barn, därigenom att han har låtit Jesus uppstå,
såsom ock är skrivet i andra psalmen: 'Du är min Son, jag har i dag fött dig.'
Och att han har låtit honom uppstå från de döda, så att han icke mer skall vända tillbaka till förgängelsen, det har han sagt med dessa ord: 'Jag skall uppfylla åt eder de heliga löften som jag i trofasthet har givit åt David.'
Därför säger han ock i en annan psalm: 'Du skall icke låta din Helige se förgängelsen.'
När David i sin tid hade tjänat Guds vilja, avsomnade han ju och blev samlad till sina fäder och såg förgängelsen;
men den som Gud har uppväckt, han har icke sett förgängelsen.
Så mån I nu veta, mena bröder, att genom honom syndernas förlåtelse förkunnas för eder,
och att i honom var och en som tror bliver rättfärdig och friad ifrån allt det varifrån I icke under Moses' lag kunden bliva friade.
Sen därför till, att över eder icke må komma det som är sagt hos profeterna:
'Sen här, I föraktare, och förundren eder, och bliven till intet; ty en gärning utför jag i edra dagar, en gärning som I alls icke skullen tro, om den förtäljdes för eder.'»
När de sedan gingo därifrån, bad men dem att de nästa sabbat skulle tala för dem om samma sak.
Och när församlingen åtskildes, följde många judar och gudfruktiga proselyter med Paulus och Barnabas.
Dessa talade då till dem och förmanade dem att stadigt hålla sig till Guds nåd.
Följande sabbat kom nästan hela staden tillsammans för att höra Guds ord.
Då nu judarna sågo det myckna folket, uppfylldes de av nitälskan och foro ut i smädelser och motsade det som Paulus talade.
Då togo Paulus och Barnabas mod till sig och sade: »Guds ord måste i första rummet förkunnas för eder.
Men eftersom I stöten det bort ifrån eder och icke akten eder själva värdiga det eviga livet, så vända vi oss nu till hedningarna.
Ty så har Herren bjudit oss: 'Jag har satt dig till ett ljus för hednafolken, för att du skall bliva till frälsning intill jordens ända.'»
När hedningarna hörde detta, blevo de glada och prisade Herrens ord; och de kommo till tro, så många det var beskärt att få evigt liv.
Och Herrens ord utbredde sig över hela landet.
Men judarna uppeggade de ansedda kvinnor som »fruktade Gud», så ock de förnämsta männen i staden, och uppväckte en förföljelse mot Paulus och Barnabas och drevo dem bort ifrån sin stads område.
Dessa skuddade då stoftet av sina fötter mot dem och begåvo sig till Ikonium.
Och lärjungarna uppfylldes alltmer av glädje och helig ande.
På samma sätt tillgick det i Ikonium: de gingo in i judarnas synagoga och talade så, att en stor hop av både judar och greker kommo till tro;
men de judar som voro ohörsamma retade upp hedningarna och väckte deras förbittring mot bröderna.
Så vistades de där en längre tid och predikade frimodigt, i förtröstan på Herren, och han gav vittnesbörd åt sitt nådesord, i det att han lät tecken och under ske genom dem.
Men folket i staden delade sig, så att somliga höllo med judarna, andra åter med apostlarna.
Och när sedan, både ibland hedningar och ibland judar med deras föreståndare, en storm hade blivit uppväckt emot dem, och man ville misshandla och stena dem,
flydde de, så snart de förstodo huru det var, till städerna Lystra och Derbe i Lykaonien och till trakten omkring dem.
Och där förkunnade de evangelium.
I Lystra fanns nu en man som satt där oförmögen att bruka sina fötter, ty allt ifrån sin moders liv hade han varit ofärdig och hade aldrig kunnat gå.
Denne hörde på, när Paulus talade.
Och då Paulus fäste sina ögon på honom och såg att han hade tro, så att han kunde bliva botad,
sade han med hög röst: »Res dig upp och stå på dina fötter.»
Då sprang mannen upp och begynte gå.
När folket såg vad Paulus hade gjort, hovo de upp sin röst och ropade på lykaoniskt tungomål: »Gudarna hava stigit ned till oss i människogestalt.»
Och de kallade Barnabas för Jupiter, men Paulus kallade de för Merkurius, eftersom det var han som förde ordet.
Och prästen vid det Jupiterstempel som låg utanför staden förde fram tjurar och kransar till portarna och ville jämte folket anställa ett offer.
Men när apostlarna, Barnabas och Paulus, fingo höra detta, revo de sönder sina kläder och sprungo ut bland folket och ropade
och sade: »I män, vad är det I gören?
Också vi äro människor, av samma natur som I, och vi förkunna för eder evangelium, att I måsten omvända eder från dessa fåfängliga avgudar till den levande Guden, 'som har gjort himmelen och jorden och havet och allt vad i dem är'.
Han har under framfarna släktens tider tillstatt alla hedningar att gå sina egna vägar.
Dock har han icke låtit sig vara utan vittnesbörd, ty han har bevisat eder välgärningar, i det han har givit eder regn och fruktbara tider från himmelen och så vederkvickt edra hjärtan med mat och glädje.»
Genom sådana ord stillade de med knapp nöd folket, så att man icke offrade åt dem.
Men några judar kommo dit från Antiokia och Ikonium.
Dessa drogo folket över på sin sida och stenade Paulus och släpade honom ut ur staden, i tanke att han var död.
Men sedan lärjungarna hade samlat sig omkring honom, reste han sig upp och gick in i staden.
Dagen därefter begav han sig med Barnabas åstad därifrån till Derbe.
Och de förkunnade evangelium i den staden och vunno ganska många lärjungar.
Sedan vände de tillbaka till Lystra och Ikonium och Antiokia
och styrkte lärjungarnas själar, i det de förmanade dem att stå fasta i tron och sade dem, att det är genom mycken bedrövelse som vi måste ingå i Guds rike.
Därefter utvalde de åt dem »äldste» för var särskild församling och anbefallde dem efter bön och fastor åt Herren, som de nu trodde på.
Sedan färdades de vidare genom Pisidien och kommo till Pamfylien.
Där förkunnade de ordet i Perge och foro sedan ned till Attalia.
Därifrån avseglade de till Antiokia, samma ort varifrån de hade blivit utsända, sedan man hade anbefallt dem åt Guds nåd, för det verk som de nu hade fullbordat.
Och när de hade kommit dit, kallade de tillhopa församlingen och omtalade för dem huru stora ting Gud hade gjort med dem, och huru han för hedningarna hade öppnat en dörr till tro.
Sedan vistades de där hos lärjungarna en ganska lång tid.
Men från Judeen kommo några män ditned och lärde bröderna så: »Om I icke låten omskära eder, såsom Moses har stadgat, så kunnen I icke bliva frälsta.»
Då uppstod söndring, och Paulus och Barnabas kommo i ett ganska skarpt ordskifte med dem.
Det bestämdes därför, att Paulus och Barnabas och några andra av dem skulle, för denna tvistefrågas skull, fara upp till apostlarna och de äldste i Jerusalem.
Och församlingen utrustade dem för resan, och de foro genom Fenicien och Samarien och förtäljde utförligt om hedningarnas omvändelse och gjorde därmed alla bröderna stor glädje.
När de sedan kommo fram till Jerusalem, mottogos de av församlingen och av apostlarna och de äldste och omtalade huru stora ting Gud hade gjort med dem.
Men några ifrån fariséernas parti, vilka hade kommit till tro, stodo upp och sade att man borde omskära dem och bjuda dem att hålla Moses' lag.
Då trädde apostlarna och de äldste tillsammans för att överlägga om denna sak.
Och sedan man länge hade förhandlat därom, stod Petrus upp och sade till dem: »Mina bröder, I veten själva att Gud, för lång tid sedan, bland eder utvalde mig att vara den genom vilkens mun hedningarna skulle få höra evangelii ord och komma till tro.
Och Gud, som känner allas hjärtan, gav dem sitt vittnesbörd, därigenom att han lät dem, likaväl som oss, undfå den helige Ande.
Och han gjorde ingen åtskillnad mellan oss och dem, i det att han genom tron renade deras hjärtan.
Varför fresten I då nu Gud, genom att på lärjungarnas hals vilja lägga ett ok som varken våra fäder eller vi hava förmått bära?
Vi tro ju fastmer att det är genom Herren Jesu nåd som vi bliva frälsta, vi likaväl som de.»
Då teg hela menigheten, och man hörde på Barnabas och Paulus, som förtäljde om huru stora tecken och under Gud genom dem hade gjort bland hedningarna.
När de hade slutat att tala, tog Jakob till orda och sade: »Mina bröder, hören mig.
Simeon har förtäljt huru Gud först så skickade, att han bland hedningarna fick ett folk som kunde kallas efter hans namn.
Därmed stämmer ock överens vad profeterna hava talat; ty så är skrivet:
'Därefter skall jag komma tillbaka och åter bygga upp Davids förfallna hydda; ja, dess ruiner skall jag bygga upp och så upprätta den igen,
för att ock övriga människor skola söka Herren, alla hedningar som hava uppkallats efter mitt namn.
Så säger Herren, han som skall göra detta,
såsom han ock har vetat det förut av evighet.'
Därför är min mening att man icke bör betunga sådana som hava varit hedningar, men omvänt sig till Gud,
utan allenast skriva till dem att de skola avhålla sig från avgudastyggelser och från otukt och från köttet av förkvävda djur och från blod.
Ty Moses har av ålder sina förkunnare i alla städer, då han ju var sabbat föreläses i synagogorna.»
Därefter beslöto apostlarna och de äldste, tillika med hela församlingen, att bland sig utvälja några män, som jämte Paulus och Barnabas skulle sändas till Antiokia; och de valde Judas, som kallades Barsabbas, och Silas, vilka bland bröderna voro ledande män.
Och man översände genom dem följande skrivelse: »Apostlarna och de äldste, edra bröder, hälsa eder, I bröder av hednisk börd, som bon i Antiokia, Syrien och Cilicien.
Alldenstund vi hava hört att några som hava kommit från oss hava förvirrat eder med sitt tal och väckt oro i edra själar, utan att de hava haft något uppdrag av oss,
så hava vi enhälligt kommit till det beslutet att utvälja några män, som vi skulle sända till eder jämte Barnabas och Paulus, våra älskade bröder,
vilka hava vågat sina liv för vår Herres, Jesu Kristi, namns skull.
Alltså sända vi nu Judas och Silas, vilka ock muntligen skola kungöra detsamma för eder.
Den helige Ande och vi hava nämligen beslutit att icke pålägga eder någon ytterligare börda, utöver följande nödvändiga föreskrifter:
att I skolen avhålla eder från avgudaofferskött och från blod och från köttet av förkvävda djur och från otukt.
Om I noga tagen eder till vara för detta, så skall det gå eder väl.
Faren väl.»
De fingo så begiva sig åstad och kommo ned till Antiokia.
Där kallade de tillsammans menigheten och lämnade fram brevet.
Och när menigheten läste detta, blevo de glada över det hugnesamma budskapet.
Judas och Silas, som själva voro profeter, talade därefter många förmaningens ord till bröderna och styrkte dem.
Och sedan de hade uppehållit sig där någon tid, fingo de i frid fara ifrån bröderna tillbaka till dem som hade sänt dem.
275440
Men Paulus och Barnabas vistades fortfarande i Antiokia, där de undervisade och, jämte många andra förkunnade evangelii ord från Herren.
Efter någon tid sade Paulus till Barnabas: »Låt oss nu fara tillbaka och besöka våra bröder, i alla de städer där vi hava förkunnat Herrens ord, och se till, huru det är med dem.»
Barnabas ville då att de skulle taga med sig Johannes, som ock kallades Markus.
Men Paulus fann icke skäligt att taga med sig en man som hade övergivit dem i Pamfylien och icke följt med dem till deras arbete.
Och så skarp blev deras tvist att de skilde sig ifrån varandra; och Barnabas tog med sig Markus och avseglade till Cypern.
Men Paulus utvalde åt sig Silas; och sedan han av bröderna hade blivit anbefalld åt Herrens nåd, begav han sig åstad
och färdades genom Syrien och Cilicien och styrkte församlingarna.
Han kom då också till Derbe och till Lystra.
Där fanns en lärjunge vid namn Timoteus, som var son av en troende judisk kvinna och en grekisk fader,
och som hade gott vittnesbörd om sig av bröderna i Lystra och Ikonium.
Paulus ville nu att denne skulle fara med honom.
För de judars skull som bodde i dessa trakter tog han honom därför till sig och omskar honom, ty alla visste att hans fader var grek.
Och när de sedan foro genom städerna, meddelade de församlingarna till efterföljd de stadgar som voro fastställda av apostlarna och de äldste i Jerusalem.
Så styrktes nu församlingarna i tron, och brödernas antal förökades för var dag.
Sedan togo de vägen genom Frygien och det galatiska landet; de förhindrades nämligen av den helige Ande att förkunna ordet i provinsen Asien.
Och när de hade kommit fram emot Mysien, försökte de att fara in i Bitynien, men Jesu Ande tillstadde dem det icke.
Då begåvo de sig över Mysien ned till Troas.
Här visade sig för Paulus i en syn om natten en macedonisk man, som stod där och bad honom och sade: »Far över till Macedonien och hjälp oss.»
När han hade sett denna syn, sökte vi strax någon lägenhet att fara därifrån till Macedonien, ty vi förstodo nu att Gud hade kallat oss att förkunna evangelium för dem.
Vi lade alltså ut från Troas och foro raka vägen till Samotrace och dagen därefter till Neapolis
och sedan därifrån till Filippi.
Denna stad, en romersk koloni, är den första i denna del av Macedonien.
I den staden vistades vi någon tid.
På sabbatsdagen gingo vi utom stadsporten, längs med en flod, till en plats som gällde såsom böneställe.
Där satte vi oss ned och talade med de kvinnor som hade samlats dit.
Och en kvinna som »fruktade Gud», en purpurkrämerska från staden Tyatira, vid namn Lydia, lyssnade till samtalet; och Herren öppnade hennes hjärta, så att hon aktade på det som Paulus talade.
Och sedan hon jämte sitt husfolk hade låtit döpa sig, bad hon oss och sade: »Eftersom I ansen mig vara en kvinna som tror på Herren, så kommen in i mitt hus och stannen där.»
Och hon nödgade oss därtill.
Och det hände sig en gång, då vi gingo ned till bönestället, att vi mötte en tjänsteflicka, som hade en spådomsande i sig och genom sina spådomar skaffade sina herrar mycken inkomst.
Denne följde efter Paulus och oss andra och ropade och sade: »Dessa män äro Guds, den Högstes, tjänare, och de förkunna för eder frälsningens väg.»
Så gjorde hon under många dagar.
Men Paulus tog illa vid sig och vände sig om och sade till anden: »I Jesu Kristi namn bjuder jag dig att fara ut ur henne.»
Och anden for ut i samma stund.
Men när hennes herrar sågo att det för dem var slut med allt hopp om vidare inkomst, grepo de Paulus och Silas och släpade dem till torget inför överhetspersonerna.
Och sedan de hade fört dem tid fram, till domarna, sade de: »Dessa män uppväcka stor oro i vår stad; de äro judar
och vilja införa stadgar som det för oss, såsom romerska medborgare, icke är lovligt att antaga eller hålla.»
Också folket reste sig upp emot dem, och domarna läto slita av dem deras kläder och bjödo att man skulle piska dem med spön.
Och sedan de hade låtit giva dem många slag, kastade de dem i fängelse och bjödo fångvaktaren att hålla dem i säkert förvar.
Då denne fick en så sträng befallning, satte han in dem i det innersta fängelserummet och fastgjorde deras fötter i stocken.
Vid midnattstiden voro Paulus och Silas stadda i bön och lovade Gud med sång, och de andra fångarna hörde på dem.
Då kom plötsligt en stark jordstöt, så att fängelsets grundvalar skakades; och i detsamma öppnades alla dörrar, och allas bojor löstes.
Då vaknade fångvaktaren; och när han fick se fängelsets dörrar öppna, drog han sitt svärd och ville döda sig själv, i tanke att fångarna hade kommit undan.
Men Paulus ropade med hög röst och sade: »Gör dig intet ont; ty vi äro alla här.»
Då lät han hämta ljus och sprang in och föll ned för Paulus och Silas, bävande.
Därefter förde han ut dem och sade: »I herrar, vad skall jag göra för att bliva frälst?»
De svarade: »Tro på Herren Jesus, så bliver du med ditt hus frälst.»
Och de förkunnade Guds ord för honom och för alla dem som voro i hans hus.
Och redan under samma timme på natten tog han dem till sig och tvådde deras sår och lät strax döpa sig med allt sitt husfolk.
Och han förde dem upp i sitt hus och dukade ett bord åt dem och fröjdade sig över att han med allt sitt hus hade kommit till tro på Gud.
Men när det hade blivit dag, sände domarna åstad rättstjänarna och läto säga: »Släpp ut männen.»
Fångvaktaren underrättade då Paulus härom och sade: »Domarna hava sänt bud att I skolen släppas ut.
Gån därför nu eder väg i frid.»
Men Paulus sade till dem: »De hava offentligen låtit gissla oss, utan dom och rannsakning, oss som äro romerska medborgare, och hava kastat oss i fängelse; nu vilja de också i tysthet släppa oss ut!
Nej, icke så; de måste själva komma och taga oss ut.»
Rättstjänarna inberättade detta för domarna.
När dessa hörde att de voro romerska medborgare, blevo de förskräckta.
Och de gingo dit och talade goda ord till dem och togo dem ut och bådo dem lämna staden.
När de så hade kommit ut ur fängelset, begåvo de sig hem till Lydia.
Och sedan de där hade träffat bröderna och talat förmaningens ord till dem, drogo de vidare.
Och de foro över Amfipolis och Apollonia och kommo så till Tessalonika.
Där hade judarna en synagoga;
i den gick Paulus in, såsom hans sed var.
Och under tre sabbater talade han där med dem, i det han utgick ifrån skrifterna
och utlade dem och bevisade att Messias måste lida och uppstå från de döda; och han sade: »Denne Jesus som jag förkunnar för eder är Messias.»
Och några av dem läto övertyga sig och slöto sig till Paulus och Silas; så gjorde ock en stor hop greker som »fruktade Gud», likaså ganska många av de förnämsta kvinnorna.
Då grepos judarna av nitälskan och togo med sig allahanda dåligt folk ifrån gatan och ställde till folkskockning och oroligheter i staden och trängde fram mot Jasons hus och ville draga dem ut inför folket.
Men när de icke funno dem, släpade de Jason och några av bröderna inför stadens styresmän och ropade: »Dessa män, som hava uppviglat hela världen, hava nu också kommit hit;
och Jason har tagit emot dem i sitt hus.
De göra alla tvärtemot kejsarens påbud och säga att en annan, en som heter Jesus, är konung.
Så väckte de oro bland folket och hos stadens styresmän, när de hörde detta.
Dessa läto då Jason och de andra ställa borgen för sig och släppte dem därefter lösa.
Men strax om natten blevo Paulus och Silas av bröderna sända åstad till Berea.
Och när de hade kommit dit, gingo de till judarnas synagoga.
Dessa voro ädlare till sinnes än judarna i Tessalonika; de togo emot ordet med all villighet och rannsakade var dag skrifterna, för att se om det förhölle sig såsom nu sades.
Många av dem kommo därigenom till tro, likaså ganska många ansedda grekiska kvinnor och jämväl män.
Men när judarna i Tessalonika fingo veta att Guds ord förkunnades av Paulus också i Berea, kommo de dit och uppviglade också där folket och väckte oro bland dem.
Strax sände då bröderna Paulus åstad ända ned till havet, men både Silas och Timoteus stannade kvar på platsen.
De som ledsagade Paulus förde honom vidare till Aten och foro så därifrån tillbaka, med bud till Silas och Timoteus att dessa med det snaraste skulle komma till honom.
Men, Paulus nu väntade på dem i Aten, upprördes han i sin ande, när han såg huru uppfylld staden var med avgudabilder.
Han höll därför i synagogan samtal med judarna och med dem som »fruktade Gud», så ock på torget, var dag, med dem som han träffade där
Också några filosofer, dels av epikuréernas skola, dels av stoikernas, gåvo sig i ordskifte med honom.
Och somliga sade: »Vad kan väl denne pratmakare vilja säga?»
Andra åter: »Han tyckes vara en förkunnare av främmande gudar.»
De evangelium om Jesus och om uppståndelsen.
Och de grepo honom och förde honom till Areopagen och sade: »Kunna vi få veta vad det är för en ny lära som du förkunnar?
Ty det är förunderliga ting som du talar oss i öronen.
Vi vilja nu veta vad detta skall betyda.»
Det var nämligen så med alla atenare, likasom ock med de främlingar som hade bosatt sig bland dem, att de icke hade tid och håg för annat än att tala om eller höra på något nytt för dagen.
Då trädde Paulus fram mitt på Areopagen och sade: »Atenare, jag ser av allting att I ären mycket ivriga gudsdyrkare.
Ty medan jag har gått omkring och betraktat edra helgedomar, har jag ock funnit ett altare med den inskriften: 'Åt en okänd Gud.'
Om just detta väsende, som I sålunda dyrken utan att känna det, är det jag nu kommer med budskap till eder.
Den Gud som har gjort världen och allt vad däri är, han som är Herre över himmel och jord, han bor icke i tempel som äro gjorda med händer,
ej heller låter han betjäna sig av människohänder, såsom vore han i behov av något, han som själv åt alla giver liv, anda och allt.
Och han har skapat människosläktets alla folk, alla från en enda stamfader, till att bosätta sig utöver hela jorden; och han har fastställt för dem bestämda tider och utstakat de gränser inom vilka de skola bo --
detta för att de skola söka Gud, om de till äventyrs skulle kunna treva sig fram till honom och finna honom; fastän han ju icke är långt ifrån någon enda av oss.
Ty i honom är det som vi leva och röra oss och äro till, såsom ock några av edra egna skalder hava sagt: 'Vi äro ju ock av hans släkt.'
Äro vi nu av Guds släkt, så böra vi icke mena att gudomen är lik någonting av guld eller silver eller sten, något som är danat genom mänsklig konst och uppfinning.
Med sådana okunnighetens tider har Gud hittills haft fördrag, men nu bjuder han människorna att de alla allestädes skola göra bättring.
Ty han har fastställt en dag då han skall 'döma världen med rättfärdighet', genom en man som han har bestämt därtill; och han har åt alla givit en bekräftelse härpå, i det att han har låtit honom uppstå från de döda.»
När de hörde talas om att »uppstå från de döda», drevo somliga gäck därmed, andra åter sade: »Vi vilja höra dig tala härom ännu en gång.»
Med detta besked gick Paulus bort ifrån dem.
Dock slöto sig några män till honom och kommo till tro.
Bland dessa var Dionysius, han som tillhörde Areopagens domstol, så ock en kvinna vid namn Damaris och några andra jämte dem.
Därefter lämnade Paulus Aten och kom till Korint.
Där träffade han en jude vid namn Akvila, bördig från Pontus, vilken nyligen hade kommit från Italien med sin hustru Priscilla.
(Klaudius hade nämligen påbjudit att alla judar skulle lämna Rom.)
Till dessa båda slöt han sig nu,
och eftersom han hade samma hantverk som de, stannade han kvar hos dem, och de arbetade tillsammans; de voro nämligen till yrket tältmakare.
Och i synagogan höll han var sabbat samtal och övertygade både judar och greker.
När sedan Silas och Timoteus kommo ditned från Macedonien, var Paulus helt upptagen av att förkunna ordet, i det att han betygade för judarna att Jesus var Messias.
Men när dessa stodo emot honom och foro ut i smädelser, skakade han stoftet av sina kläder och sade till dem: »Edert blod komme över edra egna huvuden.
Jag är utan skuld och går nu till hedningarna.»
Och han gick därifrån och tog in hos en man vid namn Titius Justus, som »fruktade Gud»; denne hade sitt hus invid synagogan.
Men Krispus, synagogföreståndaren, kom med hela sitt hus till tro på Herren; också många andra korintier som hörde honom trodde och läto döpa sig.
Och i en syn om natten sade Herren till Paulus: »Frukta icke, utan tala och tig icke;
ty jag är med dig, och ingen skall komma vid dig och göra dig skada.
Jag har ock mycket folk i denna stad.»
Så uppehöll han sig där bland dem ett år och sex månader och undervisade i Guds ord.
Men när Gallio var landshövding i Akaja, reste sig judarna, alla tillhopa, upp mot Paulus och förde honom inför domstolen
och sade: »Denne man förleder människorna att dyrka Gud på ett sätt som är emot lagen.»
När då Paulus ville öppna sin mun och tala, sade Gallio till judarna: »Vore något brott eller något ont och arglistigt dåd begånget, då kunde väl vara skäligt att jag tålmodigt hörde på eder, I judar.
Men är det någon tvistefråga om ord och namn eller om eder egen lag, så mån I själva avgöra saken; i sådana mål vill jag icke vara domare.»
Och så visade han bort dem från domstolen.
Då grepo de alla gemensamt Sostenes, synagogföreståndaren, och slogo honom inför domstolen; och Gallio frågade alls icke därefter.
Men Paulus stannade där ännu ganska länge.
Därpå tog han avsked av bröderna och avseglade till Syrien, åtföljd av Priscilla och Akvila, sedan han i Kenkrea hade låtit raka sitt huvud; han hade nämligen bundit sig genom ett löfte.
Så kommo de till Efesus, och där lämnade Paulus dem.
Själv gick han in i synagogan och gav sig i samtal med judarna.
Och de bådo honom att han skulle stanna där något längre; men han samtyckte icke därtill,
utan tog avsked av dem med de orden: »Om Gud vill, skall jag vända tillbaka till eder.»
Och så lämnade han Efesus.
Och när han hade kommit till Cesarea, begav han sig upp och hälsade på hos församlingen och for därefter ned till Antiokia.
Sedan han hade uppehållit sig där någon tid, for han vidare, och färdades först genom det galatiska landet och därefter genom Frygien och styrkte alla lärjungarna.
Men till Efesus kom en jude vid namn Apollos, bördig från Alexandria, en lärd man, mycket förfaren i skrifterna.
Denne sade blivit undervisad om »Herrens väg» och talade, brinnande i anden, och undervisade grundligt om Jesus, fastän han allenast hade kunskap om Johannes' döpelse.
Han begynte ock att frimodigt tala i synagogan.
När Priscilla och Akvila hörde honom, togo de honom till sig och undervisade honom grundligare om »Guds väg».
Och då han sedan ville fara till Akaja, skrevo bröderna till lärjungarna där och uppmanade dem att taga vänligt emot honom.
Och när han hade kommit fram, blev han dem som trodde till mycken hjälp, genom den nåd han hade undfått.
Ty med stor kraft vederlade han judarna offentligen och bevisade genom skrifterna att Jesus var Messias.
Medan Apollos var i Korint, kom Paulus, sedan han hade farit genom de övre delarna av landet, ned till Efesus.
Där träffade han några lärjungar.
Och han frågade dessa: »Undfingen I helig ande, när I kommen till tro?»
De svarade honom: »Nej, vi hava icke ens hört att helig ande är given.»
Han frågade: »Vilken döpelse bleven I då döpta med?»
De svarade: »Vi döptes med Johannes' döpelse»
Då sade Paulus: »Johannes' döpelse var en döpelse till bättring; och han sade därvid till folket, att det var på den som skulle komma efter honom, det är på Jesus, som de skulle tro.»
Sedan de hade hört detta, läto de döpa sig i Herren Jesu namn.
Och när Paulus lade händerna på dem, kom den helige Ande över dem, och de talade tungomål och profeterade.
Och tillsammans voro de vid pass tolv män.
Därefter gick han in i synagogan; och under tre månader samtalade han där, frimodigt och övertygande, med dem om Guds rike.
Men när några av dem förhärdade sig och voro ohörsamma och inför menigheten talade illa om »den vägen», vände han sig ifrån dem och avskilde lärjungarna och samtalade sedan dagligen med dessa i Tyrannus' lärosal.
Så fortgick det i två år, och alla provinsen Asiens inbyggare, både judar och greker, fingo på detta sätt höra Herrens ord.
Och Gud gjorde genom Paulus kraftgärningar av icke vanligt slag.
Man till och med tog handkläden och förkläden, som hade varit i beröring med hans kropp, och lade dem på de sjuka; och sjukdomarna veko då ifrån dem, och de onda andarna foro ut.
Men också några kringvandrande judiska besvärjare företogo sig nu att över dem som voro besatta av onda andar nämna Herren Jesu namn; de sade: »Jag besvär eder vid den Jesus som Paulus predikar.
Bland dem som så gjorde voro sju söner av en viss Skevas, en judisk överstepräst.
Men den onde anden svarade då och sade till dem: »Jesus känner jag, Paulus är mig ock väl bekant men vilka ären I?»
Och mannen som var besatt av den onde anden störtade sig på dem och övermannade både den ene och den andre; han betedde sig så våldsamt mot dem, att de måste fly ut ur huset, nakna och sargade.
Och detta blev bekant för alla Efesus' invånare, både judar och greker, och fruktan föll över dem alla, och Herren Jesu namn blev storligen prisat.
Och många av dem som hade kommit till tro trädde fram och bekände sin synd och omtalade vad de hade gjort.
Och ganska många av dem som hade övat vidskepliga konster samlade ihop sina böcker och brände upp dem i allas åsyn.
Och när man räknade tillsammans vad böckerna voro värda, fann man att värdet uppgick till femtio tusen silverpenningar.
På detta sätt hade Herrens ord mäktig framgång och visade sin kraft.
Efter allt detta bestämde sig Paulus genom Andens tillskyndelse, att över Macedonien och Akaja fara till Jerusalem.
Och han sade: »Sedan jag har varit där, måste jag ock se Rom.»
Han sände då två av sina medhjälpare, Timoteus och Erastus, åstad till Macedonien, men själv stannade han ännu någon tid i provinsen Asien.
Vid den tiden uppstod ganska mycket oväsen angående »den vägen».
Där fanns nämligen en guldsmed, vid namn Demetrius, som förfärdigade Dianatempel av silver och därmed skaffade hantverkarna en ganska stor inkomst.
Han kallade tillhopa dessa, jämte andra som hade liknande arbete, och sade: »I man, I veten att det är detta arbete som giver oss vår goda bärgning;
men nu sen och hören I att denne Paulus icke allenast i Efesus, utan i nästan hela provinsen Asien genom sitt tal har förlett ganska mycket folk, i det han säger att de gudar som göras med människohänder icke äro gudar.
Och det är fara värt, icke allenast att denna vår hantering kommer i missaktning, utan ock att den stora gudinnan Dianas helgedom bliver räknad för intet, och att jämväl denna gudinna, som hela provinsen Asien, ja, hela världen dyrkar, kommer att lida avbräck i sitt stora anseende.»
När de hörde detta, blevo de fulla av vrede och skriade: »Stor är efesiernas Diana!»
Och hela staden kom i rörelse, och alla stormade på en gång till skådebanan och släpade med sig Gajus och Aristarkus, två macedonier som voro Paulus' följeslagare
Paulus ville då gå in bland folket men lärjungarna tillstadde honom det icke.
Också några asiarker, som voro hans vänner, sände bud till honom och bådo honom att han icke skulle giva sig in på skådebanan.
Och de skriade, den ene så och den andre så; ty menigheten var upprörd, och de flesta visste icke varför de hade kommit tillsammans.
Då drog man ur folkhopen fram Alexander, som judarna sköto framför sig.
Och Alexander gav tecken med handen att han ville hålla ett försvarstal inför folket.
Men när de märkte att han var jude, begynte de ropa, alla med en mun, och skriade under ett par timmars tid: »Stor är efesiernas Diana!»
Men stadens kansler lugnade folket och sade: »Efesier, finnes då någon människa som icke vet, att efesiernas stad är vårdare av den stora Dianas tempel och den bild av henne, som har fallit ned från himmelen?
Eftersom ju ingen kan bestrida detta, bören I hålla eder lugna och icke företaga eder något förhastat.
Emellertid haven I dragit fram dessa män, som icke äro helgerånare, ej heller smäda vår gudinna,
Om nu Demetrius och de hantverkare som hålla ihop med honom hava sak mot någon, så finnas ju domstolssammanträden och landshövdingar.
Må de alltså göra upp saken med varandra inför rätta.
Och haven I något att andraga som går därutöver, så må sådant avgöras i den lagliga folkförsamlingen.
På grund av det som i dag har skett löpa vi ju till och med fara att bliva anklagade för upplopp, fastän vi icke hava gjort något ont; och någon giltig anledning till denna folkskockning kunna vi icke heller uppgiva.»
Med dessa ord fick han menigheten att skiljas åt.
Då nu oroligheterna voro stillade, kallade Paulus lärjungarna till sig och talade till dem förmaningens ord; och sedan han hade tagit avsked av dem, begav han sig åstad för att fara till Macedonien.
Och när han hade färdats genom det landet och jämväl där talat många förmaningens ord, kom han till Grekland.
Där uppehöll han sig i tre månader.
När han sedan tänkte avsegla därifrån till Syrien, beslöt han, eftersom judarna förehade något anslag mot honom, att göra återfärden genom Macedonien.
Och med honom följde Sopater, Pyrrus' son, från Berea, och av tessalonikerna Aristarkus och Sekundus, vidare Gajus från Derbe och Timoteus, slutligen Tykikus och Trofimus från provinsen Asien.
Men dessa foro i förväg och inväntade oss i Troas.
Sedan, efter det osyrade brödets högtid, avseglade vi andra ifrån Filippi och träffade dem på femte dagen åter i Troas; och där vistades vi i sju dagar.
På första veckodagen voro vi församlade till brödsbrytelse, och Paulus, som tänkte fara vidare dagen därefter, samtalade med bröderna.
Och samtalet drog ut ända till midnattstiden;
och ganska många lampor voro tända i den sal i övre våningen, där vi voro församlade.
Invid fönstret satt då en yngling vid namn Eutykus, och när Paulus talade så länge, föll denne i djup sömn och blev så överväldigad av sömnen, att han störtade ned från tredje våningen; och när man tog upp honom, var han död
Då gick Paulus ned och lade sig över honom och fattade om honom och sade: »Klagen icke så; ty livet är ännu kvar i honom.»
Sedan gick han åter upp, och bröt brödet och åt, och samtalade ytterligare ganska länge med dem, ända till dess att det dagades; först då begav han sig i väg.
Och de förde ynglingen hem levande och kände sig nu icke litet tröstade.
Men vi andra gingo i förväg ombord på skeppet och avseglade till Assos, där vi tänkte taga Paulus ombord; ty så hade han förordnat, eftersom han själv tänkte fara land vägen.
Och när han sammanträffade med oss i Assos, togo vi honom ombord och kommo sedan till Mitylene.
Därifrån seglade vi vidare och kommo följande dag mitt för Kios.
Dagen därefter lade vi till vid Samos; och sedan vi hade legat över i Trogyllium, kommo vi nästföljande dag till Miletus.
Paulus hade nämligen beslutit att segla förbi Efesus, för att icke fördröja sig i provinsen Asien; ty han påskyndade sin färd, för att, om det bleve honom möjligt, till pingstdagen kunna vara i Jerusalem.
Men från Miletus sände han bud till Efesus och kallade till sig församlingens äldste.
Och när de hade kommit till honom, sade han till dem: »I veten själva på vad sätt jag hela tiden, ifrån första dagen då jag kom till provinsen Asien, har umgåtts med eder:
huru jag har tjänat Herren i all ödmjukhet, under tårar och prövningar, som hava vållats mig genom judarnas anslag.
Och I veten att jag icke har dragit mig undan, när det gällde något som kunde vara eder nyttigt, och att jag icke har försummat att offentligen och hemma i husen predika för eder och undervisa eder.
Ty jag har allvarligt uppmanat både judar och greker att göra bättring och vända sig till Gud och tro på vår Herre Jesus.
Och se, bunden i anden begiver jag mig nu till Jerusalem, utan att veta vad där skall vederfaras mig;
allenast det vet jag, att den helige Ande i den ene staden efter den andra betygar för mig och säger att bojor och bedrövelser vänta mig.
Dock anser jag mitt liv icke vara av något värde för mig själv, om jag blott får väl fullborda mitt lopp och vad som hör till det ämbete jag har mottagit av Herren Jesus: att vittna om Guds nåds evangelium.
Och se, jag vet nu att I icke mer skolen få se mitt ansikte, I alla bland vilka jag har gått omkring och predikat om riket.
Därför betygar jag för eder nu i dag att jag icke bär skuld för någons blod.
Ty jag har icke undandragit mig att förkunna för eder allt Guds rådslut.
Så haven nu akt på eder själva och på hela den hjord i vilken den helige Ande har satt eder till föreståndare, till att vara herdar för Guds församling, som han har vunnit med sitt eget blod.
Jag vet, att sedan jag har skilts från eder svåra ulvar skola komma in bland eder, och att de icke skola skona hjorden.
Ja, bland eder själva skola män uppträda, som tala vad förvänt är, för att locka lärjungarna att följa sig.
Vaken därför, och kommen ihåg att jag i tre års tid, natt och dag, oavlåtligen under tårar har förmanat var och en särskild av eder.
Och nu anbefaller jag eder åt Gud och hans nådesord, åt honom som förmår uppbygga eder och giva åt eder eder arvedel bland alla som äro helgade.
Silver eller guld eller kläder har jag icke åstundat av någon.
I veten själva att dessa mina händer hava gjort tjänst, för att skaffa nödtorftigt uppehälle åt mig och åt dem som hava varit med mig.
I allt har jag genom mitt föredöme visat eder att man så, under eget arbete, bör taga sig an de svaga och komma ihåg Herren Jesu ord, huru han själv sade: 'Saligare är att giva än att taga.'»
När han hade sagt detta, föll han ned på sina knän och bad med dem alla.
Och de begynte alla att gråta bitterligen och föllo Paulus om halsen och kysste honom innerligt;
och mest sörjde de för det ordets skull som han hade sagt, att de icke mer skulle få se hans ansikte.
Och så ledsagade de honom till skeppet.
Sedan vi hade skilts ifrån dem, lade vi ut och foro raka vägen till Kos och kommo dagen därefter till Rodus och därifrån till Patara.
Där funno vi ett skepp som skulle fara över till Fenicien; på det gingo vi ombord och lade ut.
Och när vi hade fått Cypern i sikte, lämnade vi denna ö på vänster hand och seglade till Syrien och landade vid Tyrus; ty där skulle skeppet lossa sin last.
Och vi uppsökte där lärjungarna och stannade hos dem i sju dagar.
Dessa sade nu genom Andens tillskyndelse till Paulus att han icke borde begiva sig till Jerusalem.
Men när vi hade stannat där de dagarna ut, bröto vi upp därifrån och gåvo oss i väg, ledsagade av dem alla, med hustrur och barn, ända utom staden.
Och på stranden föllo vi ned på våra knän och bådo
och togo sedan avsked av varandra.
Därefter stego vi ombord på skeppet, och de andra vände tillbaka hem igen.
Från Tyrus kommo vi till Ptolemais, och därmed avslutade vi sjöresan.
Och vi hälsade på hos bröderna där och stannade hos dem en dag.
Men följande dag begåvo vi oss därifrån och kommo till Cesarea.
Där togo vi in hos evangelisten Filippus, en av de sju, och stannade kvar hos honom.
Denne hade fyra ogifta döttrar, som ägde profetisk gåva.
Under den tid av flera dagar, som vi stannade där, kom en profet, vid namn Agabus, dit ned från Judeen.
När denne hade kommit till oss, tog han Paulus' bälte och band därmed sina händer och fötter och sade: »Så säger den helige Ande: 'Den man som detta bälte tillhör, honom skola judarna så binda i Jerusalem, och sedan skola de överlämna honom i hedningarnas händer.'»
När vi hörde detta, bådo såväl vi själva som bröderna i staden honom att han icke skulle begiva sig upp till Jerusalem.
Men då svarade Paulus: »Varför gråten I så och sargen mitt hjärta?
Jag är ju redo icke allenast att låta mig bindas, utan ock att dö i Jerusalem, för Herren Jesu namns skull.»
Då han alltså icke lät övertala sig, gåvo vi oss till freds och sade: »Ske Herrens vilja.»
Efter de dagarnas förlopp gjorde vi oss i ordning och begåvo oss upp till Jerusalem.
Från Cesarea följde också några av lärjungarna med oss, och dessa förde oss till en viss Mnason från Cypern, en gammal lärjunge, som vi skulle gästa hos.
Och när vi kommo till Jerusalem, togo bröderna emot oss med glädje.
Dagen därefter gick Paulus med oss andra till Jakob; dit kommo ock alla de äldste.
Och sedan han hade hälsat dem förtäljde han för dem alltsammans, det ena med det andra, som Gud genom hans arbete hade gjort bland hedningarna.
När de hörde detta, prisade de Gud.
Och de sade till honom: »Du ser, käre broder, huru många tusen judar det är som hava kommit till tro, och alla nitälska de för lagen.
Nu har det blivit dem sagt om dig, att du lär alla judar som bo spridda bland hedningarna att avfalla från Moses, i det du säger att de icke behöva omskära sina barn, ej heller i övrigt vandra efter vad stadgat är.
Vad är då att göra?
Helt visst skall man få höra att du har kommit hit.
Gör därför såsom vi nu vilja säga dig.
Vi hava här fyra män som hava bundit sig genom ett löfte.
Tag med dig dessa, och låt helga dig tillsammans med dem, och åtag dig omkostnaderna för dem, så att de kunna låta raka sina huvuden.
Då skola alla förstå att intet av allt det som har blivit dem sagt om dig äger någon grund, utan att också du vandrar efter lagen och håller den.
Vad åter angår de hedningar som hava kommit till tro, så hava vi här beslutit och jämväl skrivit till dem, att de böra taga sig till vara för kött från avgudaoffer och för blod och för köttet av förkvävda djur och för otukt.»
Så tog då Paulus männen med sig och lät följande dag helga sig tillsammans med dem; sedan gick han in i helgedomen och gav till känna när den tid skulle gå till ända, för vilken de hade låtit helga sig, den tid före vars utgång offer skulle frambäras för var och en särskild av dem.
När de sju dagarna nästan voro ute, fingo judarna från provinsen Asien se honom i helgedomen och uppviglade då allt folket.
Och de grepo honom
och ropade: »I män av Israel, kommen till hjälp!
Här är den man som allestädes lär alla sådant som är emot vårt folk och emot lagen och emot denna plats.
Därtill har han nu ock fört greker in i helgedomen och oskärat denna heliga plats.»
De hade nämligen förut sett efesiern Trofimus i staden tillsammans med honom och menade att Paulus hade fört denne in i helgedomen.
Och hela staden kom i rörelse, och folket skockade sig tillsammans.
Och då de nu hade gripit Paulus, släpade de honom ut ur helgedomen, varefter portarna genast stängdes igen.
Men just som de stodo färdiga att dräpa honom, anmäldes det hos översten för den romerska vakten att hela Jerusalem var i uppror.
Denne tog då strax med sig krigsmän och hövitsmän och skyndade ned till dem.
Och när de fingo se översten och krigsmännen, upphörde de att slå Paulus
Översten gick då fram och tog honom i förvar och bjöd att man skulle fängsla honom med två kedjor.
Och han frågade vem han var och vad han hade gjort.
Men bland folket ropade den ene så, den andre så.
Då han alltså för larmets skull icke kunde få något säkert besked, bjöd han att man skulle föra honom till kasernen.
Och när han kom fram till trappan, trängde folket så våldsamt på, att han måste bäras av krigsmännen,
ty folkhopen följde efter och skriade: »Bort med honom!»
Då nu Paulus skulle föras in i kasernen, sade han till översten: »Tillstädjes det mig att säga något till dig?»
Han svarade: »Kan du tala grekiska?
Är du då icke den egyptier som för en tid sedan ställde till 'dolkmännens' uppror, de fyra tusens, och förde dem ut i öknen?»
Då svarade Paulus: »Nej, jag är en judisk man från Tarsus, medborgare alltså i en betydande stad i Cilicien.
Men jag beder dig, tillstäd mig att tala till folket.»
Och han tillstadde honom det.
Då gav Paulus från trappan, där han stod, med handen ett tecken åt folket.
Och sedan där hade blivit helt tyst, talade han till dem på hebreiska och sade:
»Bröder och fäder, hören vad jag nu inför eder vill tala till mitt försvar.»
När de hörde att han talade till dem på hebreiska, blevo de ännu mer stilla.
Och han fortsatte:
»Jag är en judisk man, född i Tarsus i Cilicien, men uppfostrad här i staden och undervisad vid Gamaliels fötter, efter fädernas lag i all dess stränghet.
Och jag var en man som nitälskade för Gud, såsom I allasammans i dag gören.
Jag förföljde 'den vägen' ända till döds, och både män och kvinnor lät jag binda och sätta i fängelse;
det vittnesbördet kan översteprästen och de äldstes hela råd giva mig.
Också fick jag av dem brev till bröderna i Damaskus; och jag begav mig dit, för att fängsla jämväl dem som voro där och föra dem till Jerusalem, så att de kunde bliva straffade.
Men när jag var på vägen och nalkades Damaskus, hände sig vid middagstiden att ett starkt sken från himmelen plötsligt kringstrålade mig.
Och jag föll ned till marken och hörde då en röst som sade till mig: 'Saul, Saul, varför förföljer du mig?'
Då svarade jag: 'Vem är du, Herre?'
Han sade till mig: 'Jag är Jesus från Nasaret, den som du förföljer.'
Och de som voro med mig sågo väl skenet, men hörde icke rösten av den som talade till mig.
Då frågade jag: 'Vad skall jag göra, Herre?'
Och Herren svarade mig: 'Stå upp och gå in i Damaskus; där skall allt det bliva dig sagt, som är dig förelagt att göra.'
Men eftersom jag, till följd av det starka skenet, icke mer kunde se togo mina följeslagare mig vid handen och ledde mig, så att jag kom in i Damaskus.
Där fanns en efter lagen fram man, Ananias, vilken hade gott vittnesbörd om sig av alla judar som bodde där.
Denne kom nu och trädde fram till mig och sade: 'Saul, min broder, hav din syn igen.'
Och i samma stund fick jag min syn igen och såg upp på honom.
Då sade han: 'Våra fäders Gud har utsett dig till att känna hans vilja och till att se den Rättfärdige och höra ord från hans mun.
Ty du skall vara hans vittne inför alla människor och vittna om vad du har sett och hört.
Varför dröjer du då nu?
Stå upp och låt döpa dig och avtvå dina synder, och åkalla därvid hans namn.'
Men när jag hade kommit tillbaka till Jerusalem, hände sig, medan jag bad i helgedomen, att jag föll i hänryckning
och såg honom och hörde honom säga till mig: 'Skynda dig med hast bort ifrån Jerusalem; ty de skola icke här taga emot ditt vittnesbörd om mig.'
Men jag sade: 'Herre, de veta själva att det var jag som överallt i synagogorna lät fängsla och gissla dem som trodde på dig.
Och när Stefanus', ditt vittnes, blod utgöts, var ock jag tillstädes och gillade vad som skedde och vaktade de mäns kläder, som dödade honom.'
Då sade han till mig: Gå; jag vill sända dig åstad långt bort till hedningarna.'»
Ända till dess att han sade detta hade de hört på honom.
Men nu hovo de upp sin röst och ropade: »Bort ifrån jorden med den människan!
Det är icke tillbörligt att en sådan får leva.»
Då de så skriade och därvid revo av sig sina kläder och kastade stoft upp i luften,
bjöd översten att man skulle föra in honom i kasernen, och gav befallning om att man skulle förhöra honom under gisselslag, så att han finge veta varför de så ropade mot honom.
Men när de redan hade sträckt ut honom till gissling, sade Paulus till den hövitsman som stod där: »Är det lovligt för eder att gissla en romersk medborgare, och det utan dom och rannsakning?»
När hövitsmannen hörde detta, gick han till översten och underrättade honom härom och sade: »Vad är det du tänker göra?
Mannen är ju romersk medborgare.»
Då gick översten dit och frågade honom: »Säg mig, är du verkligen romersk medborgare?»
Han svarade: »Ja.»
Översten sade då: Mig har det kostat en stor summa penningar att köpa den medborgarrätten.»
Men Paulus sade: »Jag däremot har den redan genom födelsen.»
Männen som skulle hava förhört honom drogo sig då strax undan och lämnade honom.
Och när översten nu hade fått veta att han var romersk medborgare, blev också han förskräckt, vid tanken på att han hade låtit fängsla honom.
Då han emellertid ville få säkert besked om varför Paulus anklagades av judarna, låt han dagen därefter taga av honom bojorna och bjöd översteprästerna och hela Stora rådet att komma tillsammans.
Sedan lät han föra Paulus ditned och ställde honom inför dem.
Och Paulus fäste ögonen på Rådet och sade: »Mina bröder, allt intill denna dag har jag vandrat inför Gud med ett i allo gott samvete.»
Då befallde översteprästen Ananias dem som stodo bredvid honom, att de skulle slå honom på munnen.
Paulus sade då till honom: »Gud skall slå dig, du vitmenade vägg.
Du sitter här för att döma mig efter lagen, och ändå bjuder du, tvärtemot lagen, att man skall slå mig!»
Då sade de som stodo därbredvid: »Smädar du Guds överstepräst?»
Paulus svarade: »Jag visste icke, mina bröder, att han var överstepräst.
Det är ju skrivet: 'Mot en hövding i ditt folk skall du icke tala onda ord.'»
Nu hade Paulus märkt att den ena delen av dem utgjordes av sadducéer och den andra av fariséer.
Därför sade han med ljudelig röst inför Rådet: »Mina bröder, jag är farisé, en avkomling av fariséer.
Det är för vårt hopps skull, för de dödas uppståndelses skull, som jag står här inför rätta.»
Knappt hade han sagt detta, förrän en strid uppstod mellan fariséerna och sadducéerna, så att hopen blev delad.
Sadducéerna säga nämligen att det icke finnes någon uppståndelse, ej heller någon ängel eller ande, men fariséerna bekänna sig tro på både det ena och det andra.
Och man begynte ropa och larma; och några skriftlärde som hörde till fariséernas parti stodo upp och begynte ivrigt disputera med de andra och sade: »Vi finna intet ont hos denne man.
Kanhända har en ande eller en ängel verkligen talat med honom.»
Då nu en så häftig strid hade uppstått, fruktade översten att de skulle slita Paulus i stycken, och bjöd manskapet gå ned och rycka honom undan dem och föra honom till kasernen.
Natten därefter kom Herren och stod framför honom och sade: »Var vid gott mod; ty såsom du har vittnat om mig i Jerusalem, så måste du ock vittna i Rom.»
När det sedan hade blivit dag, sammangaddade sig judarna och förpliktade sig med dyr ed att varken äta eller dricka, förrän de hade dräpt Paulus.
Och det var mer än fyrtio män som så hade sammansvurit sig.
Dessa gingo till översteprästerna och de äldste och sade: »Vi hava med dyr ed förpliktat oss att ingenting smaka, förrän vi hava dräpt Paulus.
Så mån I nu, tillsammans med Rådet, hemställa hos översten att han låter föra honom ned till eder, detta under föregivande att I tänken grundligare undersöka hans sak.
Vi skola då vara redo att röja honom ur vägen, innan han hinner fram.»
Men Paulus' systerson fick höra om försåtet.
Han kom därför till kasernen och gick ditin och omtalade för Paulus vad han hade hört.
Paulus bad då att en av hövitsmännen skulle komma till honom, och sade: »För denne yngling till översten; ty han har en underrättelse att lämna honom.»
Denne tog honom då med sig och förde honom till översten och sade: »Fången Paulus har kallat mig till sig och bett mig föra denne yngling till dig, ty han har något att säga dig.»
Då tog översten honom vid handen och gick avsides med honom och frågade honom: »Vad är det för en underrättelse du har att lämna mig?»
Han svarade: »Judarna hava kommit överens om att bedja dig att du i morgon låter föra Paulus ned till Rådet, detta under föregivande att det tänker skaffa sig grundligare kunskap om honom.
Gör dem nu icke till viljes häri; ty mer än fyrtio av dem ligga i försåt för honom och hava med dyr ed förpliktat sig att varken äta eller dricka, förrän de hava röjt honom ur vägen.
Och nu äro de redo och vänta allenast på att du skall bevilja deras begäran.»
Översten bjöd då ynglingen att icke för någon omtala att han hade yppat detta för honom, och lät honom sedan gå.
Därefter kallade han till sig två av hövitsmännen och sade till dem: »Låten två hundra krigsmän göra sig redo att i natt vid tredje timmen avgå till Cesarea, så ock sjuttio ryttare och två hundra spjutbärare.»
Och han tillsade dem att skaffa åsnor, som de skulle låta Paulus rida på så att han oskadd kunde föras till landshövdingen Felix.
Och han skrev ett brev, så lydande:
»Klaudius Lysias hälsar den ädle landshövdingen Felix.
Denne man blev gripen av judarna, och det var nära att han hade blivit dödad av dem.
Då kom jag tillstädes med mitt manskap och tog honom ifrån dem, sedan jag hade fått veta att han var romersk medborgare.
Men då jag också ville veta vad de anklagade honom för, lät jag ställa honom inför deras Stora råd.
Jag fann då att anklagelsen mot honom gällde några tvistefrågor i deras lag, men att han icke var anklagad för något som förtjänade död eller fängelse.
Sedan har jag fått kännedom om att något anslag förehaves mot honom, och därför sänder jag honom nu strax till dig.
Jag har jämväl bjudit hans anklagare att inför dig föra sin talan mot honom.»
Så togo nu krigsmännen Paulus, såsom det hade blivit dem befallt, och förde honom om natten till Antipatris.
Dagen därefter vände de själva tillbaka till kasernen och läto ryttarna färdas vidare med honom.
När dessa kommo till Cesarea, lämnade de fram brevet till landshövdingen och förde jämväl Paulus fram inför honom.
Sedan han hade läst brevet, frågade han från vilket landskap han var; och när han hade fått veta att han var från Cilicien, sade han:
»Jag skall höra vad du har att säga, när också dina anklagare hava kommit tillstädes.»
Och så bjöd han att man skulle förvara honom i Herodes' borg.
Fem dagar därefter for översteprästen Ananias ditned med några av de äldste och en sakförare, Tertullus; dessa anmälde inför landshövdingen klagomål mot Paulus.
Och sedan denne hade blivit förekallad, begynte Tertullus sitt anklagelsetal; han sade:
»Att vi genom dig åtnjuta mycken frid och ro, och att genom din försorg, ädle Felix, goda åtgärder hava blivit vidtagna för detta folk, det erkänna vi på allt sätt och allestädes, med många tacksägelser.
Men för att icke alltför länge besvära dig beder jag att du, i din mildhet, ville höra allenast några få ord av oss.
Vi hava funnit att denne är en fördärvlig man, som uppväcker strid bland alla judar i hela världen, och att han är en huvudman för nasaréernas parti.
Han har ock försökt att oskära helgedomen; därför grepo vi honom,
278430
och du kan nu själv anställa rannsakning med honom och så skaffa dig kännedom om allt det som vi anklaga honom för.»
De andra judarna instämde häri och påstodo att det förhöll sig så.
Då landshövdingen nu gav tecken åt Paulus att han skulle tala, tog han till orda och sade: »Eftersom jag vet att du nu i många år har varit domare över detta folk, försvarar jag min sak med frimodighet.
Du kan själv lätt förvissa dig om att det icke är mer än tolv dagar sedan jag kom upp till Jerusalem för att tillbedja.
Och varken i helgedomen eller i synagogorna eller ute i staden har man funnit mig tvista med någon eller ställa till folkskockning.
Ej heller kunna de inför dig bevisa det som de nu anklaga mig för.
Men det bekänner jag för dig att jag, i enlighet med 'den vägen', vilken de kalla en partimening, så tjänar mina fäders Gud, att jag tror allt vad som är skrivet i lagen och i profeterna,
och att jag har samma hopp till Gud som dessa hysa, att de döda skola uppstå, både rättfärdiga och orättfärdiga.
Därför lägger också jag mig vinn om att alltid hava ett okränkt samvete inför Gud och människor.
Så kom jag nu, efter flera års förlopp, tillbaka för att överlämna några allmosor till mitt folk och för att frambära offer.
Därunder påträffades jag i helgedomen, sedan jag hade låtit helga mig, utan att hava vållat någon folkskockning eller något larm,
av några judar från provinsen Asien, vilka nu borde vara här tillstädes inför dig och framställa sina klagomål, om de hava något att anklaga mig för.
Eller ock må dessa som äro här tillstädes säga vad orätt de funno mig skyldig till, när jag stod inför Stora rådet,
om det icke skulle vara i fråga om detta enda ord, som jag ljudeligen uttalade, där jag stod ibland dem: 'Det är för de dödas uppståndelses skull som jag i dag står inför rätta här bland eder.'»
Men Felix, som mycket väl kände till »den vägen», uppsköt målet och sade: »När översten Lysias kommer hit ned, vill jag undersöka eder sak.»
Och han befallde hövitsmannen att hålla honom i förvar, dock så, att man skulle behandla honom milt och icke hindra någon av hans närmaste från att vara honom till tjänst.
Någon tid därefter infann sig Felix tillsammans med sin hustru Drusilla, som var judinna; och han lät hämta Paulus och hörde honom om tron på Kristus Jesus.
Men när Paulus talade med dem om rättfärdighet och återhållsamhet och om den tillstundande domen, blev Felix förskräckt och sade: »Gå din väg för denna gång; när jag får läglig tid, vill jag kalla dig till mig.»
Han hoppades också att han skulle få penningar av Paulus, varför han ock ganska ofta lät hämta honom och samtalade med honom.
När två år voro förlidna, fick Felix till efterträdare Porcius Festus.
Och eftersom Felix ville göra judarna sig bevågna, lämnade han Paulus kvar i fängelset.
Tre dagar efter det att Festus hade tillträtt hövdingdömet for han från Cesarea upp till Jerusalem.
Översteprästerna och de förnämsta bland judarna anmälde då inför honom klagomål mot Paulus.
För att få denne i sitt våld anhöllo de hos Festus och begärde såsom en ynnest, att han skulle låta hämta honom till Jerusalem.
De ville nämligen lägga försåt för honom, så att de kunde döda honom under vägen.
Festus svarade då att Paulus hölls i förvar i Cesarea, och att han själv tänkte inom kort fara dit tillbaka.
Och han tillade: »De bland eder som det vederbör må alltså fara dit ned med mig och framlägga sin anklagelse mot mannen, om han är skyldig till något ont.»
Sedan han hade vistats hos dem högst åtta eller tio dagar, kom han åter ned till Cesarea.
Dagen därefter satte han sig på domarsätet och bjöd att Paulus skulle föras fram.
När denne hade infunnit sig, omringades han av de judar som hade kommit ned från Jerusalem, och dessa framställde nu många svåra beskyllningar.
Men de förmådde icke bevisa dem,
ty Paulus försvarade sig och visade att han icke på något sätt hade försyndat sig, vare sig mot judarnas lag eller mot helgedomen eller mot kejsaren.
Men Festus ville göra judarna sig bevågna och frågade Paulus och sade: »Vill du fara upp till Jerusalem och där stå till rätta inför mig i denna sak?»
Paulus svarade: »Jag står här inför kejserlig domstol, och av sådan domstol bör jag dömas.
Mot judarna har jag intet orätt gjort, såsom du själv mycket väl vet.
Om jag nu eljest är skyldig till något orätt och har gjort något som förtjänar döden, så vill jag icke undandraga mig att dö; men om deras anklagelser mot mig äro utan grund, så kan ingen giva mig till pris åt dem.
Jag vädjar till kejsaren.» --
Sedan Festus därefter hade överlagt med sitt råd, svarade han: »Till kejsaren har du vädjat, till kejsaren skall du ock få fara.»
Efter några dagars förlopp kommo konung Agrippa och Bernice till Cesarea och hälsade på hos Festus.
Medan de nu i flera dagar vistades där, framlade Festus Paulus' sak för konungen och sade: »Felix har här lämnat efter sig en man såsom fånge;
och när jag var i Jerusalem, anmälde judarnas överstepräster och äldste klagomål mot honom och begärde att han skulle dömas skyldig.
Men jag svarade dem att det icke var romersk sed att prisgiva någon människa, förrän den anklagade hade fått stå ansikte mot ansikte med sina anklagare och haft tillfälle att försvara sig mot anklagelsen.
Sedan de hade kommit med mig hit, satte jag mig alltså utan uppskov, dagen därefter, på domarsätet och bjöd att mannen skulle föras fram.
Men när hans anklagare uppträdde, anförde de mot honom ingen beskyllning för sådana förbrytelser som jag hade tänkt mig;
de voro allenast i tvist med honom om några frågor som rörde deras särskilda gudsdyrkan, och angående en viss Jesus, som är död, men om vilken Paulus påstod att han lever.
Då jag var villrådig huru jag skulle göra med undersökningen härom, frågade jag om han ville fara till Jerusalem och där stå till rätta i denna sak.
När Paulus då sade sig vilja vädja till kejsaren och begärde att bliva hållen i förvar, för att sedan undergå rannsakning inför honom, bjöd jag att han skulle hållas i förvar, till dess jag kunde sända honom till kejsaren.»
Då sade Agrippa till Festus: »Jag skulle också själv gärna vilja höra den mannen.»
Han svarade: »I morgon skall du få höra honom.»
Dagen därefter kommo alltså Agrippa och Bernice, med stor ståt, och gingo in i domsalen, tillika med överstarna och de förnämsta männen i staden; och på Festus' befallning blev Paulus införd.
Då sade Festus: »Konung Agrippa, och alla I andra som ären har tillstädes med oss, I sen här den man för vilkens skull hela hopen av judar, både i Jerusalem och här, har legat över mig med sina rop att han icke borde få leva längre.
Jag för min del har kommit till insikt om att han icke har gjort något som förtjänar döden;
men då han nu själv har vädjat till kejsaren, har jag beslutit att sända honom till denne.
Jag har emellertid icke något säkert besked om honom att giva min höge herre, när jag skriver.
Därför har jag fört honom fram inför eder, och först och främst inför dig, konung Agrippa, för att jag, efter det att rannsakning har; blivit hållen, skall få veta vad jag bör skriva.
Ty det synes mig vara orimligt att sända åstad en fånge, utan att på samma gång giva till känna vad han är anklagad för.»
Agrippa sade nu till Paulus: »Det tillstädjes dig att tala för din sak.»
Då räckte Paulus ut handen och talade så till sitt försvar:
»Jag skattar mig lycklig att jag, i fråga om allt det som judarna anklaga mig för, i dag skall försvara mig inför dig, konung Agrippa,
som så väl känner judarnas alla stadgar och tvistefrågor.
Därför beder jag dig höra mig med tålamod.
Hurudant mitt liv allt ifrån ungdomen har varit, det veta alla judar, ty jag har ju från tidiga år framlevat det bland mitt folk och i Jerusalem.
Och sedan lång tid tillbaka känna de om mig -- såframt de nu vilja tillstå det -- att jag har tillhört det strängaste partiet i vår gudsdyrkan och levat såsom farisé.
Och nu står jag här till rätta för vårt hopp om det som Gud har lovat våra fäder,
det vartill ock våra tolv stammar, under det de tjäna Gud med iver både natt och dag, hoppas att nå fram.
För det hoppets skull, o konung, är jag anklagad av judarna.
Varför hålles det då bland eder för otroligt att Gud uppväcker döda?
Jag för min del menade alltså att jag med all makt borde strida mot Jesu, nasaréens, namn;
så gjorde jag ock i Jerusalem.
Och många av de heliga inspärrade jag i fängelse, sedan jag av översteprästerna hade fått fullmakt därtill; och när man ville döda dem, röstade ock jag därför.
Och överallt i synagogorna försökte jag, gång på gång, att genom straff tvinga dem till hädelse.
I mitt raseri mot dem gick jag så långt, att jag förföljde dem till och med ända in i utländska städer.
När jag nu i detta ärende var på väg till Damaskus, med fullmakt och uppdrag från översteprästerna,
fick jag under min färd, o konung, mitt på dagen se ett sken från himmelen, klarare än solens glans, kringstråla mig och mina följeslagare.
Och vi föllo alla ned till jorden, och jag hörde då en röst säga till mig på hebreiska: 'Saul, Saul, varför förföljer du mig'?
Det är dig svårt att spjärna mot udden.'
Då sade jag: 'Vem är du, Herre?'
Herren svarade: 'Jag är Jesus, den som du förföljer.
Men res dig upp och stå på dina fötter; ty därför har jag visat mig för dig, att jag har velat utse dig till en tjänare och ett vittne, som skall vittna både om huru du nu har sett mig, och om huru jag vidare skall uppenbara mig för dig.
Och jag skall rädda dig såväl från ditt eget folk som från hedningarna.
Ty till dem sänder jag dig,
för att du skall öppna deras ögon, så att de omvända sig från mörkret till ljuset, och från Satans makt till Gud, på det att de må, genom tron på mig, undfå syndernas förlåtelse och få sin lott bland dem som äro helgade.'
Så blev jag då, konung Agrippa, icke ohörsam mot den himmelska synen,
utan predikade först för dem som voro i Damaskus och i Jerusalem, och sedan över hela judiska landet och för hedningarna, att de skulle göra bättring och omvända sig till Gud och göra sådana gärningar som tillhöra bättringen.
För denna saks skull var det som judarna grepo mig i helgedomen och försökte att döda mig.
Genom den hjälp som jag har undfått av Gud står jag alltså ännu i dag såsom ett vittne inför både små och stora; och jag säger intet annat, än vad profeterna och Moses hava sagt skola ske,
nämligen att Messias skulle lida och, såsom förstlingen av dem som uppstå från de döda, bära budskap om ljuset, såväl till vårt eget folk som till hedningarna.»
När han på detta satt försvarade sig, utropade Festus: »Du är från dina sinnen, Paulus; den myckna lärdomen gör dig förryckt.»
Men Paulus svarade: »Jag är icke från mina sinnen, ädle Festus; jag talar sanna ord med lugn besinning.
Konungen känner väl till dessa ting; därför talar jag också frimodigt inför honom.
Ty jag kan icke tro att något av detta är honom obekant; det har ju icke tilldragit sig i någon undangömd vrå.
Tror du profeterna, konung Agrippa?
Jag vet att du tror dem.»
Då sade Agrippa till Paulus: »Föga fattas att du övertalar mig och gör mig till kristen.»
Paulus svarade: »Vare sig det fattas litet eller fattas mycket, skulle jag önska inför Gud att icke allenast du, utan alla som i dag höra mig, måtte bliva sådana som jag är, dock med undantag av dessa bojor.»
Därefter stod konungen upp, och med honom landshövdingen och Bernice och de som sutto där tillsammans med dem.
Och när de gingo därifrån, talade de med varandra och sade: »Den mannen har icke gjort något som förtjänar död eller fängelse.»
Och Agrippa sade till Festus: »Denne man hade väl kunnat frigivas, om han icke hade vädjat till kejsaren.»
När det nu var beslutet att vi skulle avsegla till Italien, blev Paulus jämte några andra fångar överlämnad åt en hövitsman, vid namn Julius, som tillhörde den kejserliga vakten.
Och vi gingo ombord på ett skepp från Adramyttium, som skulle anlöpa provinsen Asiens kuststäder.
Så lade vi ut, och vi hade med oss Aristarkus, en macedonier från Tessalonika.
Dagen därefter lade vi till vid Sidon.
Och Julius, som bemötte Paulus med välvilja, tillstadde honom att besöka sina vänner där och åtnjuta deras omvårdnad.
När vi hade lagt ut därifrån, seglade vi under Cypern, eftersom vinden låg emot.
Och sedan vi hade seglat över havet, utanför Cilicien och Pamfylien, landade vi vid Myrra i Lycien.
Där träffade hövitsmannen på ett skepp från Alexandria, som skulle segla till Italien, och på det förde han oss ombord.
Under en längre tid gick nu seglingen långsamt, och vi kommo med knapp nöd inemot Knidus.
Och då vinden icke var oss gynnsam, seglade vi in under Kreta vid Salmone.
Det var med knapp nöd som vi kommo där förbi och hunno fram till en ort som kallades Goda hamnarna, icke långt från staden Lasea.
Härunder hade ganska lång tid hunnit förflyta, och sjöfarten begynte redan vara osäker; fastedagen var nämligen redan förbi.
Paulus varnade dem då
och sade: »I mån, jag ser att denna sjöresa kommer att medföra vedervärdigheter och stor olycka, icke allenast för last och skepp, utan ock för våra liv.»
Men hövitsmannen trodde mer på styrmannen och skepparen än på det som Paulus sade.
Och då hamnen icke låg väl till för övervintring, var flertalet av den meningen att man borde lägga ut därifrån och försöka om man kunde komma fram till Fenix, en hamn på Kreta, som ligger skyddad mot sydväst och nordväst; där skulle de sedan stanna över vintern.
Och då nu en lindrig sunnanvind blåste upp, menade de sig hava målet vunnet, och lyfte ankar och foro tätt utmed Kreta.
Men icke långt därefter kom en våldsam stormvind farande ned från ön; det var den så kallade nordostorkanen.
Då skeppet av denna rycktes med och icke kunde hållas upp mot vinden, gåvo vi efter och läto det driva.
När vi kommo under en liten ö som hette Kauda, förmådde vi dock, fastän med knapp nöd, bärga skeppsbåten.
Sedan manskapet hade dragit upp den, tillgrepo de nödhjälpsmedel och slogo tåg om skeppet.
Och då de fruktade att bliva kastade på Syrtenrevlarna, lade de ut drivankare och läto skeppet så driva.
Och eftersom vi alltjämt hårt ansattes av stormen, vräkte de dagen därefter en del av lasten över bord.
På tredje dagen kastade de med egna händer ut skeppsredskapen.
Och då under flera dagar varken sol eller stjärnor hade synts, och stormen låg ganska hårt på, hade vi icke mer något hopp om räddning.
Då nu många funnos som ingenting ville förtära, trädde Paulus upp mitt ibland dem och sade: »I män, I haden bort lyda mig och icke avsegla från Kreta; I haden då kunnat spara eder dessa vedervärdigheter och denna olycka.
Men nu uppmanar jag eder att vara vid gott mod, ty ingen av eder skall förlora sitt liv; allenast skeppet skall gå förlorat.
Ty i natt kom en ängel från den Gud som jag tillhör, och som jag också tjänar, och stod bredvid mig och sade:
'Frukta icke, Paulus.
Du skall komma att stå inför kejsaren; och se, Gud har skänkt dig alla dem som segla med dig.'
Varen därför vid gott mod, I män; ty jag har den förtröstan till Gud, att så skall ske som mig är sagt.
Men på en ö måste vi bliva kastade.»
När vi nu den fjortonde natten drevo omkring på Adriatiska havet, tyckte sjömännen sig vid midnattstiden finna att de närmade sig något land.
De lodade då och funno tjugu famnars djup.
När de hade kommit ett litet stycke längre fram lodade de åter och funno femton famnars djup.
Då fruktade de att vi skulle stöta på något skarpt grund, och kastade därför ut fyra ankaren från akterskeppet och längtade efter att det skulle dagas.
Sjömännen ville emellertid fly ifrån skeppet och firade ned skeppsbåten i havet, under föregivande att de tänkte föra ut ankaren ifrån förskeppet.
Då sade Paulus till hövitsmannen och krigsmännen: »Om icke dessa stanna kvar på skeppet, så kunnen I icke räddas.»
Då höggo krigsmännen av de tåg som höllo skeppsbåten, och läto den fara.
Medan det nu höll på att dagas, uppmanade Paulus alla att taga sig mat och sade: »Det är i dag fjorton dagar som I haven väntat och förblivit fastande, utan att förtära något.
Därför uppmanar jag eder att taga eder mat; detta skall förhjälpa eder till räddning.
Ty på ingen av eder skall ett huvudhår gå förlorat.
När han hade sagt detta, tog han ett bröd och tackade Gud i allas åsyn och bröt det och begynte äta.
Då blevo alla de andra vid gott mod och togo sig mat, också de.
Och vi voro på skeppet tillsammans två hundra sjuttiosex personer.
Sedan de hade ätit sig mätta, lättade de skeppet genom att kasta vetelasten i havet.
När det blev dag, kände de icke igen landet; men de blevo varse en vik med låg strand och beslöto då att, om möjligt, låta skeppet driva upp på denna.
De kapade så ankartågen på båda sidor och lämnade ankarna kvar i havet; tillika lösgjorde de rodren och hissade förseglet för vinden och styrde mot stranden.
De stötte då på ett rev och läto skeppet gå upp på det.
Där fastnade förskeppet och blev stående orörligt, men akterskeppet begynte brytas sönder av vågsvallet.
Då ville krigsmännen döda fångarna, för att ingen skulle kunna fly undan simmande.
Men hövitsmannen ville rädda Paulus och hindrade dem därför i deras uppsåt, och bjöd att de simkunniga först skulle kasta sig i vattnet och söka komma i land,
och att därefter de övriga skulle giva sig ut, somliga på plankor, andra på spillror av skeppet.
Så lyckades det för alla att komma välbehållna i land.
Först sedan vi hade blivit räddade, fingo vi veta att ön hette Malta.
Och infödingarna visade oss en icke vanlig välvilja; de tände upp en eld och togo oss alla med sig dit, för det påkommande regnets och för köldens skull.
När Paulus då tog upp ett fång torra kvistar som han lade på elden, kom, i följd av hettan, en huggorm fram därur och högg sig fast vid hans hand.
Då infödingarna fingo se ormen hänga där vid hans hand, sade de till varandra: »Helt visst är denne man en dråpare, som rättvisans gudinna icke tillstädjer att leva, om han nu ock har blivit räddad undan havet.»
Men han skakade ormen ifrån sig i elden och led ingen skada.
De väntade att han skulle svälla upp eller helt plötsligt falla ned död; men när de efter lång väntan fingo se att intet ont vederfors honom, ändrade de mening och sade att han var en gud.
I närheten av detta ställe var en lantgård, som tillhörde den förnämste mannen på ön, en som hette Publius; denne tog välvilligt emot oss och gav oss härbärge i tre dagar.
Nu hände sig att Publius' fader låg sjuk i en magsjukdom med feberanfall.
Paulus gick då in till honom och bad och lade händerna på honom och gjorde honom frisk.
Men när detta hade skett, kommo också de av öns övriga inbyggare som hade någon sjukdom till honom och blevo botade.
Och de bevisade oss ära på mångahanda sätt; och när vi skulle avsegla, försågo de oss med vad vi behövde.
Då tre månader voro förlidna, avseglade vi på ett skepp som hade legat vid ön över vintern; det var från Alexandria och bar Tvillinggudarnas bilder.
Och vi lade till vid Syrakusa och stannade där i tre dagar.
Därifrån foro vi längs kusten och kommo till Regium.
Dagen därefter fingo vi sunnanvind, och vi kommo så redan på andra dagen till Puteoli.
Där träffade vi på bröder, och hos dem stannade vi, på deras inbjudning, i sju dagar.
På detta sätt kommo vi till Rom.
Så snart bröderna där fingo höra om oss, gingo de oss till mötes ända till Forum Appii och Tres Taberne.
När Paulus fick se dem, tackade han Gud och fick nytt mod.
Och då vi hade kommit in i Rom, tillstaddes det Paulus att bo för sig själv, med den krigsman som skulle bevaka honom.
Tre dagar därefter kallade han tillhopa de förnämsta av judarna; och när de hade kommit tillsammans, sade han till dem: »Mina bröder, fastän jag icke har gjort något mot vårt folk eller mot fädernas stadgar, blev jag likväl i Jerusalem överlämnad i romarnas händer och fördes bort därifrån såsom fånge.
Och när de hade anställt rannsakning med mig, ville de giva mig lös, eftersom jag icke hade gjort något som förtjänade döden.
Men då judarna satte sig däremot, nödgades jag vädja till kejsaren; dock, icke som om jag hade någon anklagelse att göra mot mitt folk.
Av denna orsak har jag kallat eder hit till mig, för att få se eder och tala med eder, ty det är för Israels hopps skull som jag är bunden med denna kedja.»
Då svarade de honom: »Vi hava icke från Judeen mottagit någon skrivelse om dig, ej heller har någon av våra bröder kommit och berättat eller sagt något ont om dig.
Men vi finna skäligt att du låter oss höra huru du tänker.
Ty om det partiet är oss bekant att det allestädes mötes med gensägelse.
Sedan utsatte de en viss dag för honom, och på den kommo ännu flera till honom i hans härbärge.
Då vittnade han för dem om Guds rike och utlade vad därtill hör, och försökte att övertyga dem i fråga om Jesus, med bevis både ur Moses' lag och ur profeterna; därmed höll han på från morgonen ända till aftonen.
Och somliga läto övertyga sig av det som han sade, men andra trodde icke.
Och då de icke kunde komma överens med varandra, gingo de sin väg, och därvid sade Paulus allenast detta ord: »Rätt talade den helige Ande genom profeten Esaias till edra fäder,
när han sade: 'Gå åstad och säg till detta folk: Med hörande öron skolen I höra, och dock alls intet förstå, och med seende ögon skolen I se, och dock alls intet förnimma.
Ty detta folks hjärta har blivit förstockat; och med öronen höra de illa, och sina ögon hava de tillslutit, så att de icke se med sina ögon eller höra med sina öron eller förstå med sina hjärtan och omvända sig och bliva helade av mig'
Det mån I därför veta: till hedningarna bar denna Guds frälsning blivit sänd; de skola ock akta därpå.»
I två hela år bodde han sedan kvar i en bostad som han själv hade hyrt.