I begynnelsen skapade Gud himmel och jord.
Och jorden var öde och tom, och mörker var över djupet, och Guds Ande svävade över vattnet.
Och Gud sade: »Varde ljus»; och det vart ljus.
Och Gud såg att ljuset var gott; och Gud skilde ljuset från mörkret.
Och Gud kallade ljuset dag, och mörkret kallade han natt.
Och det vart afton, och det vart morgon, den första dagen.
Och Gud sade: »Varde mitt i vattnet ett fäste som skiljer vatten från vatten.»
Och Gud gjorde fästet, och skilde vattnet under fästet från vattnet ovan fästet; och det skedde så.
Och Gud kallade fästet himmel.
Och det vart afton, och det vart morgon, den andra dagen.
Och Gud sade: »Samle sig det vatten som är under himmelen till en särskild plats, så att det torra bliver synligt.»
Och det skedde så.
Och Gud kallade det torra jord, och vattensamlingen kallade han hav.
Och Gud såg att det var gott.
Och Gud sade: »Frambringe jorden grönska, fröbärande örter och fruktträd, som efter sina arter bära frukt, vari de hava sitt frö, på jorden.»
Och det skedde så;
jorden frambragte grönska, fröbärande örter, efter deras arter, och träd som efter sina arter buro frukt, vari de hade sitt frö.
Och Gud såg att det var gott.
Och det vart afton, och det vart morgon, den tredje dagen.
Och Gud sade: »Varde på himmelens fäste ljus som skilja dagen från natten, och vare de till tecken och till att utmärka särskilda tider, dagar och år,
och vare de på himmelens fäste till ljus som lysa över jorden.»
Och det skedde så;
Gud gjorde de två stora ljusen, det större ljuset till att råda över dagen, och det mindre ljuset till att råda över natten, så ock stjärnorna.
Och Gud satte dem på himmelens fäste till att lysa över jorden,
och till att råda över dagen och över natten, och till att skilja ljuset från mörkret.
Och Gud såg att det var gott.
Och det vart afton, och det vart morgon, den fjärde dagen.
Och Gud sade: »Frambringe vattnet ett vimmel av levande varelser; flyge ock fåglar över jorden under himmelens fäste.»
Och Gud skapade de stora havsdjuren och hela det stim av levande varelser, som vattnet vimlar av, efter deras arter, så ock alla bevingade fåglar, efter deras arter.
Och Gud såg att det var gott.
Och Gud välsignade dem och sade: »Varen fruktsamma och föröken eder, och uppfyllen vattnet i haven; föröke sig ock fåglarna på jorden.»
Och det vart afton, och det vart morgon, den femte dagen.
Och Gud sade: »Frambringe jorden levande varelser, efter deras arter, boskapsdjur och kräldjur och vilda djur, efter deras arter.»
Och det skedde så;
Gud gjorde de vilda djuren, efter deras arter, och boskapsdjuren, efter deras arter, och alla kräldjur på marken, efter deras arter.
Och Gud såg att det var gott.
Och Gud sade: »Låt oss göra människor till vår avbild, till att vara oss lika; och må de råda över fiskarna i havet och över fåglarna under himmelen och över boskapsdjuren och över hela jorden och över alla kräldjur som röra sig på jorden.»
Och Gud skapade människan till sin avbild, till Guds avbild skapade han henne, till man och kvinna skapade han dem.
Och Gud välsignade dem; Gud sade till dem: »Varen fruktsamma och föröken eder, och uppfyllen jorden och läggen den under eder; och råden över fiskarna i havet och över fåglarna under himmelen och över alla djur som röra sig på jorden.»
Och Gud sade: »Se, jag giver eder alla fröbärande örter på hela jorden och alla träd med fröbärande trädfrukt; detta skolen I hava till föda.
Men åt alla djur på jorden och åt alla fåglar under himmelen och åt allt som krälar på jorden, vad som i sig har en levande själ, åt dessa giver jag alla gröna örter till föda.»
Och det skedde så.
Och Gud såg på allt som han hade gjort, och se, det var mycket gott.
Och det vart afton, och det vart morgon, den sjätte dagen.
Så blevo nu himmelen och jorden fullbordade med hela sin härskara.
Och Gud fullbordade på sjunde dagen det verk som han hade gjort; och han vilade på sjunde dagen från allt det verk som han hade gjort.
Och Gud välsignade den sjunde dagen och helgade den, därför att han på den dagen vilade från allt sitt verk, det som Gud hade gjort, när han skapade.
Detta är berättelsen om den ordning i vilken allt blev till på himmelen och jorden, när de skapades, då när HERREN Gud gjorde jord och himmel.
Då bar jorden ännu ingen buske på marken, och ingen ört hade ännu skjutit upp på marken, ty HERREN Gud hade icke låtit regna på jorden, och ingen människa fanns, som kunde bruka jorden;
men en dimma steg upp från jorden och vattnade hela marken.
Och HERREN Gud danade människan av stoft från jorden och inblåste livsande i hennes näsa, och så blev människan en levande varelse.
Och HERREN Gud planterade en lustgård i Eden österut och satte däri människan som han hade danat.
HERREN Gud lät nämligen alla slags träd som voro ljuvliga att se på och goda att äta av växa upp ur marken, och livets träd mitt i lustgården, så ock kunskapens träd på gott och ont.
Och från Eden gick en flod ut, som vattnade lustgården; sedan delade den sig i fyra grenar.
Den första heter Pison; det är den som flyter omkring hela landet Havila, där guld finnes,
och det landets guld är gott; där finnes ock bdelliumharts och onyxsten.
Den andra floden heter Gihon; det är den som flyter omkring hela landet Kus.
Den tredje floden heter Hiddekel; det är den som har sitt lopp öster om Assyrien.
Den fjärde floden är Frat.
Så tog nu HERREN Gud mannen och satte honom i Edens lustgård, till att bruka och bevara den.
Och HERREN Gud bjöd mannen och sade: »Av alla andra träd i lustgården må du fritt äta,
men av kunskapens träd på gott och ont skall du icke äta, ty när du äter därav, skall du döden dö.»
Och HERREN Gud sade: »Det är icke gott att mannen är allena.
Jag vill göra åt honom en hjälp, en sådan som honom höves.»
Och HERREN Gud danade av jord alla markens djur och alla himmelens fåglar, och förde dem fram till mannen för att se huru denne skulle kalla dem; ty såsom mannen kallade var levande varelse, så skulle den heta.
Och mannen gav namn åt alla boskapsdjur, åt fåglarna under himmelen och åt alla markens djur.
Men för Adam fann han icke någon hjälp, sådan som honom hövdes.
Då lät HERREN Gud en tung sömn falla på mannen, och när han hade somnat, tog han ut ett av hans revben och fyllde dess plats med kött.
Och HERREN Gud byggde en kvinna av revbenet som han hade tagit av mannen, och förde henne fram till mannen.
Då sade mannen: »Ja, denna är nu ben av mina ben och kött av mitt kött.
Hon skall heta maninna, ty av man är hon tagen.»
Fördenskull skall en man övergiva sin fader och sin moder och hålla sig till sin hustru, och de skola varda ett kött.
Och mannen och hans hustru voro båda nakna och blygdes icke för varandra.
Men ormen var listigare än alla andra markens djur som HERREN Gud hade gjort; och han sade till kvinnan: »Skulle då Gud hava sagt: 'I skolen icke äta av något träd i lustgården'?»
Kvinnan svarade ormen: »Vi få äta av frukten på de andra träden i lustgården,
men om frukten på det träd som står mitt i lustgården har Gud sagt: 'I skolen icke äta därav, ej heller komma därvid, på det att I icke mån dö.'»
Då sade ormen till kvinnan: »Ingalunda skolen I dö;
men Gud vet, att när I äten därav, skola edra ögon öppnas, så att I bliven såsom Gud och förstån vad gott och ont är.»
Och kvinnan såg att trädet var gott att äta av, och att det var en lust för ögonen, och att det var ett ljuvligt träd, eftersom man därav fick förstånd, och hon tog av dess frukt och åt; och hon gav jämväl åt sin man, som var med henne, och han åt.
Då öppnades bådas ögon, och de blevo varse att de voro nakna; och de fäste ihop fikonlöv och bundo omkring sig.
Och de hörde HERREN Gud vandra i lustgården, när dagen begynte svalkas; då gömde sig mannen med sin hustru för HERREN Guds ansikte bland träden i lustgården.
Men HERREN Gud kallade på mannen och sade till honom: »Var är du?»
Han svarade: »Jag hörde dig i lustgården; då blev jag förskräckt, eftersom jag är naken; därför gömde jag mig.»
Då sade han: »Vem har låtit dig förstå att du är naken?
Har du icke ätit av det träd som jag förbjöd dig att äta av?»
Mannen svarade: »Kvinnan som du har givit mig till att vara med mig, hon gav mig av trädet, så att jag åt.»
Då sade HERREN Gud till kvinnan: »Vad är det du har gjort!»
Kvinnan svarade: »Ormen bedrog mig, så att jag åt.»
Då sade HERREN Gud till ormen: »Eftersom du har gjort detta, vare du förbannad bland alla djur, boskapsdjur och vilda djur.
På din buk skall du gå, och stoft skall du äta i alla dina livsdagar.
Och jag skall sätta fiendskap mellan dig och kvinnan, och mellan din säd och hennes säd.
Denna skall söndertrampa ditt huvud, och du skall stinga den i hälen.»
Och till kvinnan sade han: »Jag skall låta dig utstå mycken vedermöda, när du bliver havande; med smärta skall du föda dina barn.
Men till din man skall din åtrå vara, och han skall råda över dig.»
Och till Adam sade han: »Eftersom du lyssnade till din hustrus ord och åt av det träd om vilket jag hade bjudit dig och sagt: 'Du skall icke äta därav', därför vare marken förbannad för din skull.
Med vedermöda skall du nära dig av den i alla dina livsdagar;
törne och tistel skall den bära åt dig, men markens örter skola vara din föda.
I ditt anletes svett skall du äta ditt bröd, till dess du vänder åter till jorden; ty av den är du tagen.
Ty du är stoft, och till stoft skall du åter varda.»
Och mannen gav sin hustru namnet Eva, ty hon blev en moder åt allt levande.
Och HERREN Gud gjorde åt Adam och hans hustru kläder av skinn och satte på dem.
Och HERREN Gud sade: »Se, mannen har blivit såsom en av oss, så att han förstår vad gott och ont är.
Må han nu icke räcka ut sin hand och taga jämväl av livets träd och äta, och så leva evinnerligen.»
Och HERREN Gud förvisade honom ur Edens lustgård, för att han skulle bruka jorden, varav han var tagen.
Och han drev ut mannen, och satte öster om Edens lustgård keruberna jämte det ljungande svärdets lågor, för att bevaka vägen till livets träd.
Och mannen kände sin hustru Eva, och hon blev havande och födde Kain; då sade hon: »Jag har fött en man genom HERRENS hjälp.»
Och hon födde åter en son, Abel, den förres broder.
Och Abel blev en fårherde, men Kain blev en åkerman.
Och efter någon tid hände sig att Kain av markens frukt bar fram en offergåva åt HERREN.
Också Abel bar fram sin gåva, av det förstfödda i hans hjord, av djurens fett.
Och HERREN såg till Abel och hans offergåva;
men till Kain och hans offergåva såg han icke.
Då blev Kain mycket vred, och hans blick blev mörk.
Och HERREN sade till Kain: »Varför är du vred, och varför är din blick så mörk?
Är det icke så: om du har gott i sinnet, då ser du frimodigt upp; men om du icke har gott i sinnet, då lurar synden vid dörren; till dig står hennes åtrå, men du bör råda över henne.»
Och Kain talade med sin broder Abel; och när de voro ute på marken, överföll Kain sin broder Abel och dräpte honom.
Då sade HERREN till Kain: »Var är din broder Abel?»
Han svarade: »Jag vet icke; skall jag taga vara på min broder?»
Då sade han: »Vad har du gjort!
Hör, din broders blod ropar till mig från jorden.
Så vare du nu förbannad och förvisad ifrån åkerjorden, som har öppnat sin mun för att mottaga din broders blod av din hand.
När du brukar jorden, skall den icke mer giva dig sin gröda.
Ostadig och flyktig skall du bliva på jorden.»
Då sade Kain till HERREN: »Min missgärning är större än att jag kan bära den.
Se, du driver mig nu bort ifrån åkerjorden, och jag måste gömma mig undan för ditt ansikte.
Ostadig och flyktig skall jag bliva på jorden, och så skall ske att vemhelst som möter mig, han dräper mig.»
Men HERREN sade till honom: »Nej, ty Kain skall bliva hämnad sjufalt, vemhelst som dräper honom.»
Och HERREN satte ett tecken till skydd för Kain, så att ingen som mötte honom skulle slå honom ihjäl.
Så gick Kain bort ifrån HERRENS ansikte och bosatte sig i landet Nod, öster om Eden.
Och Kain kände sin hustru, och hon blev havande och födde Hanok.
Och han byggde en stad och kallade den staden Hanok, efter sin sons namn.
Och åt Hanok föddes Irad, och Irad födde Mehujael, och Mehujael födde Metusael, och Metusael födde Lemek.
Men Lemek tog sig två hustrur; den ena hette Ada, den andra Silla.
Och Ada födde Jabal; han blev stamfader för dem som bo i tält och idka boskapsskötsel.
Och hans broder hette Jubal; han blev stamfader för alla dem som hantera harpa och pipa.
Men Silla födde ock en son, Tubal-Kain; han var smed och gjorde alla slags redskap av koppar och järn.
Och Tubal-Kains syster var Naama.
Och Lemek sade till sina hustrur: »Ada och Silla, hören mina ord; I Lemeks hustrur, lyssnen till mitt tal: Se, en man dräper jag för vart sår jag får, och en yngling för var blånad jag får.
Ja, sjufalt hämnad bliver Kain, men Lemek sju- och sjuttiofalt.»
Och Adam kände åter sin hustru, och hon födde en son och gav honom namnet Set, i det hon sade: »Gud har beskärt mig en annan livsfrukt, till ersättning för Abel, eftersom Kain dräpte honom.»
Men åt Set föddes ock en son, och han gav honom namnet Enos.
Vid denna tid begynte man åkalla HERRENS namn.
Detta är stycket om Adams släkt.
När Gud skapade människor, gjorde han dem lika Gud.
Till man och kvinna skapade han dem; och han välsignade dem och gav dem namnet människa, när de blevo skapade.
När Adam var ett hundra trettio år gammal, födde han en son som var honom lik, hans avbild, och gav honom namnet Set.
Och sedan Adam hade fött Set, levde han åtta hundra år och födde söner och döttrar.
Alltså blev Adams hela levnadsålder nio hundra trettio år; därefter dog han.
När Set var ett hundra fem år gammal, födde han Enos.
Och sedan Set hade fött Enos, levde han åtta hundra sju år och födde söner och döttrar.
Alltså blev Sets hela ålder nio hundra tolv år; därefter dog han.
När Enos var nittio år gammal, födde han Kenan.
Och sedan Enos hade fött Kenan, levde han åtta hundra femton år och födde söner och döttrar.
Alltså blev Enos' hela ålder nio hundra fem år; därefter dog han.
När Kenan var sjuttio år gammal, födde han Mahalalel.
Och sedan Kenan fött Mahalalel, levde han åtta hundra fyrtio år och födde söner och döttrar.
Alltså blev Kenans hela ålder nio hundra tio år; därefter dog han.
När Mahalalel var sextiofem år gammal, födde han Jered.
Och sedan Mahalalel hade fött Jered, levde han åtta hundra trettio år och födde söner och döttrar.
Alltså blev Mahalalels hela ålder åtta hundra nittiofem år; därefter dog han.
När Jered var ett hundra sextiotvå år gammal, födde han Hanok.
Och sedan Jered hade fött Hanok, levde han åtta hundra år och födde söner och döttrar.
Alltså blev Jereds hela ålder nio hundra sextiotvå år; därefter dog han.
När Hanok var sextiofem år gammal, födde han Metusela.
Och Hanok vandrade i umgängelse med Gud i tre hundra år, sedan han hade fött Metusela, och han födde söner och döttrar.
Alltså blev Hanoks hela ålder tre hundra sextiofem år.
Sedan Hanok så hade vandrat i umgängelse med Gud, såg man honom icke mer, ty Gud tog honom bort.
När Metusela var ett hundra åttiosju år gammal, födde han Lemek.
Och sedan Metusela hade fött Lemek, levde han sju hundra åttiotvå år och födde söner och döttrar.
Alltså blev Metuselas hela ålder nio hundra sextionio år; därefter dog han.
När Lemek var ett hundra åttiotvå år gammal, födde han en son.
Och han gav honom namnet Noa, i det han sade: »Denne skall trösta oss vid vårt arbete och våra händers möda, när vi bruka jorden, som HERREN har förbannat.»
Och sedan Lemek hade fött Noa, levde han fem hundra nittiofem år och födde söner och döttrar.
Alltså blev Lemeks hela ålder sju hundra sjuttiosju år; därefter dog han.
När Noa var fem hundra år gammal, födde han Sem, Ham och Jafet.
Då nu människorna begynte föröka sig på jorden och döttrar föddes åt dem
sågo Guds söner att människornas döttrar voro fagra, och de togo till hustrur dem som de funno mest behag i.
Då sade HERREN: »Min ande skall icke bliva kvar i människorna för beständigt, eftersom de dock äro kött; så vare nu deras tid bestämd till ett hundra tjugu år.»
Vid den tiden, likasom ock efteråt, levde jättarna på jorden, sedan Guds söner begynte gå in till människornas döttrar och dessa födde barn åt dem; detta var forntidens väldiga män, som voro så namnkunniga.
Men när HERREN såg att människornas ondska var stor på jorden, och att deras hjärtans alla uppsåt och tankar beständigt voro allenast onda,
då ångrade HERREN att han hade gjort människorna på jorden, och han blev bedrövad i sitt hjärta.
Och HERREN sade: »Människorna, som jag skapade, vill jag utplåna från jorden, ja, både människor och fyrfotadjur och kräldjur och himmelens fåglar; ty jag ångrar att jag har gjort dem.»
Men Noa hade funnit nåd för HERRENS ögon.
Detta är berättelsen om Noas släkt.
Noa var en rättfärdig man och ostrafflig bland sitt släkte; i umgängelse med Gud vandrade Noa.
Och Noa födde tre söner: Sem, Ham och Jafet.
Men jorden blev alltmer fördärvad för Guds åsyn, och jorden uppfylldes av våld.
Och Gud såg att jorden var fördärvad, eftersom allt kött vandrade i fördärv på jorden.
Då sade Gud till Noa: »Jag har beslutit att göra ände på allt kött, ty jorden är uppfylld av våld som de öva; se, jag vill fördärva dem tillika med jorden.
Så gör dig nu en ark av goferträ, och inred arken med kamrar, och bestryk den med jordbeck innan och utan.
Och så skall du göra arken: Den skall vara tre hundra alnar lång, femtio alnar bred och trettio alnar hög;
en öppning för ljuset, en aln hög alltigenom, skall du göra ovantill på arken; och en dörr till arken skall du sätta på dess sida; och du skall inreda den så, att den får en undervåning, en mellanvåning och en övervåning.
Ty se, jag skall låta floden komma med vatten över jorden, till att fördärva allt kött som har i sig någon livsande, under himmelen; allt som finnes på jorden skall förgås.
Men med dig vill jag upprätta ett förbund: du skall gå in i arken med dina söner och din hustru och dina söners hustrur.
Och av allt levande, vad kött det vara må, skall du föra in i arken ett par av vart slag, för att behålla dem vid liv med dig; hankön och honkön skola de vara.
Av fåglarna, efter deras arter, av fyrfotadjuren, efter deras arter, av alla kräldjur på marken, efter deras arter, skall ett par av vart slag gå in till dig, för att du må behålla dem vid liv.
Och du skall taga till dig alla slags livsmedel, sådant som kan ätas, och samla det till dig, för att det må vara dig och dem till föda.
Och Noa gjorde så; han gjorde i alla stycken såsom Gud hade bjudit honom.
Och HERREN sade till Noa: »Gå in i arken med hela ditt hus, ty dig har jag funnit rättfärdig inför mig bland detta släkte.
Av alla rena fyrfotadjur skall du taga till dig sju par, hanne och hona, men av sådana fyrfotadjur som icke äro rena ett par, hanne och hona,
sammalunda av himmelens fåglar sju par, hankön och honkön, för att behålla deras släkten vid liv på hela jorden.
Ty sju dagar härefter skall jag låta det regna på jorden, i fyrtio dagar och fyrtio nätter, och jag skall utplåna från jorden alla varelser som jag har gjort.»
Och Noa gjorde i alla stycken såsom HERREN hade bjudit honom.
Noa var sex hundra år gammal, när floden kom med sitt vatten över jorden.
Och Noa gick in i arken med sina söner och sin hustru och sina söners hustrur, undan flodens vatten.
Och av fyrfotadjur, både rena och orena, och av fåglar och av allt som krälar på marken
gingo två och två, hankön och honkön, in till Noa i arken, såsom Gud hade bjudit Noa.
Och efter de sju dagarna kom flodens vatten över jorden.
I det år då Noa var sex hundra år gammal, i andra månaden, på sjuttonde dagen i månaden, den dagen bröto alla det stora djupets källor fram, och himmelens fönster öppnade sig,
och ett regn kom över jorden i fyrtio dagar och fyrtio nätter.
På denna samma dag gick Noa in i arken, så ock Sem, Ham och Jafet, Noas söner, vidare Noas hustru och hans söners tre hustrur med dem,
därtill alla vilda djur, efter sina arter, och alla boskapsdjur, efter sina arter, och alla kräldjur som röra sig på jorden, efter sina arter, och alla flygande djur, efter sina arter, allt vad fåglar heter, av alla slag.
De gingo in till Noa i arken, två och två av allt kött som hade i sig någon livsande.
Och de som gingo ditin voro hankön och honkön av allt slags kött, såsom Gud hade bjudit honom.
Och HERREN stängde igen om honom.
Och floden kom över jorden i fyrtio dagar, och vattnet förökade sig och lyfte arken, så att den flöt högt uppe över jorden.
Och vattnet steg och förökade sig mycket på jorden, och arken drev på vattnet.
Och vattnet steg mer och mer över jorden, och alla höga berg allestädes under himmelen övertäcktes.
Femton alnar högt steg vattnet över bergen, så att de övertäcktes.
Då förgicks allt kött som rörde sig på jorden, fåglar och boskapsdjur och vilda djur och alla smådjur som rörde sig på jorden, så ock alla människor.
Allt som fanns på det torra omkom, allt som där hade en fläkt av livsande i sin näsa.
Så utplånade han alla varelser på jorden, både människor och fyrfotadjur och kräldjur och himmelens fåglar; de utplånades från jorden, och allenast Noa räddades, jämte det som var med honom i arken.
Och vattnet fortfor att stiga över jorden i hundra femtio dagar.
Då tänkte Gud på Noa och på alla de vilda djur och alla de boskapsdjur som voro med honom i arken.
Och Gud lät en vind gå fram över jorden, så att vattnet sjönk undan;
och djupets källor och himmelens fönster tillslötos, och regnet från himmelen upphörde.
Och vattnet vek bort ifrån jorden mer och mer; efter hundra femtio dagar begynte vattnet avtaga.
Och i sjunde månaden, på sjuttonde dagen i månaden, stannade arken på Ararats berg.
Och vattnet avtog mer och mer intill tionde månaden.
I tionde månaden, på första dagen i månaden, blevo bergstopparna synliga.
Och efter fyrtio dagar öppnade Noa fönstret som han hade gjort på arken,
och lät en korp flyga ut; denne flög fram och åter, till dess vattnet hade torkat bort ifrån jorden.
Sedan lät han en duva flyga ut, för att få se om vattnet hade sjunkit undan från marken.
Men duvan fann ingen plats där hon kunde vila sin fot, utan kom tillbaka till honom i arken, ty vatten betäckte hela jorden.
Då räckte han ut sin hand och tog henne in till sig i arken.
Sedan väntade han ännu ytterligare sju dagar och lät så duvan än en gång flyga ut ur arken.
Och duvan kom till honom mot aftonen, och se, då hade hon ett friskt olivlöv i sin näbb.
Då förstod Noa att vattnet hade sjunkit undan från jorden.
Men han väntade ännu ytterligare sju dagar och lät så duvan åter flyga ut; då kom hon icke mer tillbaka till honom.
I det sexhundraförsta året, i första månaden, på första dagen i månaden, hade vattnet sinat bort ifrån jorden.
Då tog Noa av taket på arken och såg nu att marken var fri ifrån vatten.
Och i andra månaden, på tjugusjunde dagen i månaden, var jorden alldeles torr.
Då talade Gud till Noa och sade:
»Gå ut ur arken med din hustru och dina söner och dina söners hustrur.
Alla djur som du har hos dig, vad slags kött det vara må, både fåglar och fyrfotadjur och alla kräldjur som röra sig på jorden, skall du låta gå ut med dig, för att de må växa till på jorden och vara fruktsamma och föröka sig på jorden.»
Så gick då Noa ut med sina söner och sin hustru och sina söners hustrur.
Och alla fyrfotadjur, alla kräldjur och alla fåglar, alla slags djur som röra sig på jorden, gingo ut ur arken, efter sina släkten.
Och Noa byggde ett altare åt HERREN och tog av alla rena fyrfotadjur och av alla rena fåglar och offrade brännoffer på altaret.
När HERREN kände den välbehagliga lukten, sade han vid sig själv: »Jag skall härefter icke mer förbanna marken för människans skull, eftersom ju människans hjärtas uppsåt är ont allt ifrån ungdomen.
Och jag skall härefter icke mer dräpa allt levande, såsom jag nu har gjort.
Så länge jorden består, skola härefter sådd och skörd, köld och värme, sommar och vinter, dag och natt aldrig upphöra.»
Och Gud välsignade Noa och hans söner och sade till dem: »Varen fruktsamma och föröken eder, och uppfyllen jorden.
Och må fruktan och förskräckelse för eder komma över alla djur på jorden och alla fåglar under himmelen; jämte allt som krälar på marken och alla fiskar i havet vare de givna i eder hand.
Allt som rör sig och har liv skolen I hava till föda; såsom jag har givit eder gröna örter, så giver jag eder allt detta.
Kött som har i sig sin själ, det är sitt blod, skolen I dock icke äta.
Men edert eget blod, vari eder själ är, skall jag utkräva.
Jag skall utkräva det av vilket djur det vara må.
Jag skall ock av den ena människan utkräva den andres själ;
den som utgjuter människoblod, hans blod skall av människor bliva utgjutet, ty Gud har gjort människan till sin avbild.
Och varen I fruktsamma och föröken eder; växen till på jorden och föröken eder på den.»
Ytterligare sade Gud till Noa och till hans söner med honom:
»Se, jag vill upprätta ett förbund med eder, och med edra efterkommande efter eder,
och med alla levande varelser som I haven hos eder: fåglar, boskapsdjur och alla vilda djur hos eder, alla jordens djur som hava gått ut ur arken.
Jag vill upprätta ett förbund med eder: härefter skall icke mer ske att allt kött utrotas genom flodens vatten; ingen flod skall mer komma och fördärva jorden.»
Och Gud sade: »Detta skall vara tecknet till det förbund som jag gör mellan mig och eder, jämte alla levande varelser hos eder, för eviga tider:
min båge sätter jag i skyn; den skall vara tecknet till förbundet mellan mig och jorden.
Och när jag härefter låter skyar stiga upp över jorden och bågen då synes i skyn,
skall jag tänka på det förbund som har blivit slutet mellan mig och eder, jämte alla levande varelser, vad slags kött det vara må; och vattnet skall då icke mer bliva en flod som fördärvar allt kött.
När alltså bågen synes i skyn och jag ser på den, skall jag tänka på det eviga förbund som har blivit slutet mellan Gud och alla levande varelser, vad slags kött det vara må på jorden.»
Så sade nu Gud till Noa: »Detta skall vara tecknet till det förbund som jag har upprättat mellan mig och allt kött på jorden.»
Noas söner, som gingo ut ur arken, voro Sem, Ham och Jafet; men Ham var Kanaans fader.
Dessa tre voro Noas söner och från dessa hava alla jordens folk utgrenat sig.
Och Noa var en åkerman och var den förste som planterade en vingård.
Men när han drack av vinet, blev han drucken och låg blottad i sitt tält.
Och Ham, Kanaans fader, såg då sin faders blygd och berättade det för sina båda bröder, som voro utanför.
Men Sem och Jafet togo en mantel och lade den på sina skuldror, båda tillsammans, och gingo så baklänges in och täckte över sin faders blygd; de höllo därvid sina ansikten bortvända, så att de icke sågo sin faders blygd.
När sedan Noa vaknade upp från ruset och fick veta vad hans yngste son hade gjort honom, sade han:
»Förbannad vare Kanaan, en trälars träl vare han åt sina bröder!»
Ytterligare sade han: »Välsignad vare HERREN, Sems Gud, och Kanaan vare deras träl!
Gud utvidge Jafet, han tage sin boning i Sems hyddor, och Kanaan vare deras träl.»
Och Noa levde efter floden tre hundra femtio år;
alltså blev Noas hela ålder nio hundra femtio år; därefter dog han.
Detta är berättelsen om Noas söners släkt.
De voro Sem, Ham och Jafet; och åt dem föddes söner efter floden.
Jafets söner voro Gomer, Magog, Madai, Javan, Tubal, Mesek och Tiras.
Gomers söner voro Askenas, Rifat och Togarma.
Javans söner voro Elisa och Tarsis, kittéerna och dodanéerna.
Från dessa hava inbyggarna i hedningarnas Havsländer utbrett sig i sina länder, var efter sitt tungomål, efter sina släkter, i sina folk.
Hams söner voro Kus, Misraim, Put och Kanaan.
Kus' söner voro Seba, Havila, Sabta, Raema och Sabteka.
Raemas söner voro Saba och Dedan.
Men Kus födde Nimrod; han var den förste som upprättade ett välde på jorden.
Han var ock en väldig jägare inför HERREN; därför plägar man säga: »En väldig jägare inför HERREN såsom Nimrod.»
Och hans rike hade sin begynnelse i Babel, Erek, Ackad och Kalne, i Sinears land.
Från det landet drog han sedan ut till Assyrien och byggde Nineve, Rehobot-Ir och Kela,
och därtill Resen mellan Nineve och Kela; detta är »den stora staden».
Och Misraim födde ludéerna, anaméerna, lehabéerna, naftuhéerna,
patroséerna, kasluhéerna, från vilka filistéerna hava utgått, och kaftoréerna.
Och Kanaan födde Sidon, som var hans förstfödde, och Het,
så ock jebuséerna, amoréerna, girgaséerna,
hivéerna, arkéerna, sinéerna,
arvadéerna, semaréerna och hamatéerna.
Sedan utgrenade sig kananéernas släkter allt vidare,
så att kananéernas område sträckte sig från Sidon fram emot Gerar ända till Gasa, och fram emot Sodom, Gomorra, Adma och Seboim ända till Lesa.
Dessa voro Hams söner, efter deras släkter och tungomål, i deras länder och folk.
Söner föddes ock åt Sem, Jafets äldre broder, som blev stamfader för alla Ebers söner.
Sems söner voro Elam, Assur, Arpaksad, Lud och Aram.
Arams söner voro Us, Hul, Geter och Mas.
Arpaksad födde Sela, och Sela födde Eber.
Men åt Eber föddes två söner; den ene hette Peleg, ty i hans tid blev jorden fördelad; och hans broder hette Joktan.
Och Joktan födde Almodad, Selef, Hasarmavet, Jera,
Hadoram, Usal, Dikla,
Obal, Abimael, Saba,
Ofir, Havila och Jobab; alla dessa voro Joktans söner.
Och de hade sina boningsorter från Mesa fram emot Sefar, emot Östra berget.
Dessa voro Sems söner, efter deras släkter och tungomål, i deras länder, efter deras folk.
Dessa voro Noas söners släkter, efter deras ättföljd, i deras folk.
Och från dem hava folken efter floden utbrett sig på jorden.
Och hela jorden hade enahanda tungomål och talade på enahanda sätt.
Men när de bröto upp och drogo österut, funno de en lågslätt i Sinears land och bosatte sig där.
Och de sade till varandra: »Kom, låt oss slå tegel och bränna det.»
Och teglet begagnade de såsom sten, och såsom murbruk begagnade de jordbeck.
Och de sade: »Kom, låt oss bygga en stad åt oss och ett torn vars spets räcker upp i himmelen, och så göra oss ett namn; vi kunde eljest bliva kringspridda över hela jorden.»
Då steg HERREN ned för att se staden och tornet som människobarnen byggde.
Och HERREN sade: »Se, de äro ett enda folk och hava alla enahanda tungomål, och detta är deras första tilltag; härefter skall intet bliva dem omöjligt, vad de än besluta att göra.
Välan, låt oss stiga dit ned och förbistra deras tungomål, så att den ene icke förstår den andres tungomål.»
Och så spridde HERREN dem därifrån ut över hela jorden, så att de måste upphöra att bygga på staden.
Därav fick den namnet Babel, eftersom HERREN där förbistrade hela jordens tungomål; därifrån spridde ock HERREN ut dem över hela jorden.
Detta är berättelsen om Sems släkt.
När Sem var hundra år gammal, födde han Arpaksad, två år efter floden.
Och sedan Sem hade fött Arpaksad, levde han fem hundra år och födde söner och döttrar.
När Arpaksad var trettiofem år gammal, födde han Sela.
Och sedan Arpaksad hade fött Sela, levde han fyra hundra tre år och födde söner och döttrar.
När Sela var trettio år gammal, födde han Eber.
Och sedan Sela hade fött Eber, levde han fyra hundra tre år och födde söner och döttrar.
När Eber var trettiofyra år gammal, födde han Peleg.
Och sedan Eber hade fött Peleg, levde han fyra hundra trettio år och födde söner och döttrar.
När Peleg var trettio år gammal, födde han Regu.
Och sedan Peleg hade fött Regu, levde han två hundra nio år och födde söner och döttrar.
När Regu var trettiotvå år gammal, födde han Serug.
Och sedan Regu hade fött Serug, levde han två hundra sju år och födde söner och döttrar.
När Serug var trettio år gammal, födde han Nahor.
Och sedan Serug hade fött Nahor, levde han två hundra år och födde söner och döttrar.
När Nahor var tjugunio år gammal, födde han Tera.
Och sedan Nahor hade fött Tera, levde han ett hundra nitton år och födde söner och döttrar.
När Tera var sjuttio år gammal, födde han Abram, Nahor och Haran.
Och detta är berättelsen om Teras släkt.
Tera födde Abram, Nahor och Haran.
Och Haran födde Lot.
Och Haran dog hos sin fader Tera i sitt fädernesland, i det kaldeiska Ur.
Och Abram och Nahor togo sig hustrur; Abrams hustru hette Sarai, och Nahors hustru hette Milka, dotter till Haran, som var fader till Milka och Jiska.
Men Sarai var ofruktsam och hade inga barn.
Och Tera tog med sig sin son Abram och sin sonson Lot, Harans son, och sin sonhustru Sarai, som var hans son Abrams hustru; och de drogo tillsammans ut från det kaldeiska Ur på väg till Kanaans land; men när de kommo till Haran, bosatte de sig där.
Och Teras ålder blev två hundra fem år; därefter dog Tera i Haran.
Och HERREN sade till Abram: »Gå ut ur ditt land och från din släkt och från din faders hus, bort till det land som jag skall visa dig.
Så skall jag göra dig till ett stort folk; jag skall välsigna dig och göra ditt namn stort, och du skall bliva en välsignelse.
Och jag skall välsigna dem som välsigna dig, och den som förbannar dig skall jag förbanna, och i dig skola alla släkter på jorden varda välsignade.»
Och Abram gick åstad, såsom HERREN hade tillsagt honom, och Lot gick med honom.
Och Abram var sjuttiofem år gammal, när han drog ut från Haran.
Och Abram tog sin hustru Sarai och sin brorson Lot och alla ägodelar som de hade förvärvat och tjänarna som de hade skaffat sig i Haran; och de drogo åstad på väg mot Kanaans land
och kommo så till Kanaans land.
Och Abram drog fram i landet ända till den heliga platsen vid Sikem, till Mores terebint.
Och på den tiden bodde kananéerna där i landet.
Men HERREN uppenbarade sig för Abram och sade: »Åt din säd skall jag giva detta land.»
Då byggde han där ett altare åt HERREN, som hade uppenbarat sig för honom.
Sedan flyttade han därifrån till bergsbygden öster om Betel och slog där upp sitt tält, så att han hade Betel i väster och Ai i öster; och han byggde där ett altare åt HERREN och åkallade HERRENS namn.
Sedan bröt Abram upp därifrån och drog sig allt längre mot Sydlandet.
Men hungersnöd uppstod i landet, och Abram drog ned till Egypten för att bo där någon tid, eftersom hungersnöden var så svår i landet.
Men när han nalkades Egypten sade han till sin hustru Sarai: »Jag vet ju att du är en skön kvinna.
Om nu egyptierna tänka, när de få se dig: 'Hon är hans hustru', så skola de dräpa mig, under det att de låta dig leva.
Säg därför att du är min syster, så att det går mig väl för din skull, och så att jag för din skull får leva.»
Då nu Abram kom till Egypten, sågo egyptierna att hon var en mycket skön kvinna.
Och när Faraos hövdingar fingo se henne, prisade de henne för Farao, och så blev kvinnan tagen in i Faraos hus.
Och Abram blev av honom väl behandlad för hennes skull, så att han fick får, fäkreatur och åsnor, tjänare och tjänarinnor, åsninnor och kameler.
Men HERREN hemsökte Farao och hans hus med stora plågor för Sarais, Abrams hustrus, skull.
Då kallade Farao Abram till sig och sade: »Vad har du gjort mot mig!
Varför lät du mig icke veta att hon var din hustru?
Varför sade du: 'Hon är min syster' och vållade så, att jag tog henne till hustru åt mig?
Se, här har du nu din hustru, tag henne och gå.»
Och Farao gav sina män befallning om honom, att de skulle ledsaga honom till vägs med hans hustru och allt vad han ägde.
Så drog då Abram upp från Egypten med sin hustru och allt vad han ägde, och Lot jämte honom, till Sydlandet.
Och Abram var mycket rik på boskap och på silver och guld.
Och han färdades ifrån lägerplats till lägerplats och kom så från Sydlandet ända till Betel, till det ställe där hans tält förut hade stått, mellan Betel och Ai,
dit där han förra gången hade rest ett altare.
Och där åkallade Abram HERRENS namn.
Men Lot, som drog med Abram, hade också får och fäkreatur och tält.
Och landet räckte icke till för dem, så att de kunde bo tillsammans; ty deras ägodelar voro för stora för att de skulle kunna bo tillsammans;
och tvister uppstodo mellan Abrams och Lots boskapsherdar.
Tillika bodde på den tiden kananéerna och perisséerna där i landet.
Då sade Abram till Lot: »Icke skall någon tvist vara mellan mig och dig, och mellan mina herdar och dina herdar; vi äro ju fränder.
Ligger icke hela landet öppet för dig?
Skilj dig ifrån mig; vill du åt vänster, så går jag åt höger, och vill du åt höger, så går jag åt vänster.»
Då lyfte Lot upp sina ögon och såg att hela Jordanslätten överallt var vattenrik.
Innan HERREN fördärvade Sodom och Gomorra, var den nämligen såsom HERRENS lustgård, såsom Egyptens land, ända fram emot Soar.
Så utvalde då Lot åt sig hela Jordanslätten.
Och Lot bröt upp och drog österut, och de skildes så från varandra.
Abram förblev boende i Kanaans land, och Lot bodde i städerna på Slätten och drog med sina tält ända inemot Sodom.
Men folket i Sodom var mycket ont och syndigt inför HERREN.
Och HERREN sade till Abram, sedan Lot hade skilt sig från honom: »Lyft upp dina ögon och se, från den plats där du står, mot norr och söder och öster och väster.»
Ty hela det land som du nu ser skall jag giva åt dig och din säd för evärdlig tid.
Och jag skall låta din säd bliva såsom stoftet på jorden; kan någon räkna stoftet på jorden, så skall ock din säd kunna räknas.
Stå upp och drag igenom landet efter dess längd och dess bredd, ty åt dig skall jag giva det.»
Och Abram drog åstad med sina tält och kom och bosatte sig vid Mamres terebintlund invid Hebron; och han byggde där ett altare åt HERREN.
På den tid då Amrafel var konung i Sinear, Arjok konung i Ellasar, Kedorlaomer konung i Elam och Tideal konung över Goim, hände sig
att dessa begynte krig mot Bera, konungen i Sodom, Birsa, konungen i Gomorra, Sinab, konungen i Adma, Semeber, konungen i Seboim, och mot konungen i Bela, det är Soar.
De förenade sig alla och tågade till Siddimsdalen, där Salthavet nu är.
I tolv år hade de varit under Kedorlaomer, men i det trettonde året hade de avfallit.
Så kom nu i det fjortonde året Kedorlaomer med de konungar som voro på hans sida; och de slogo rafaéerna i Asterot-Karnaim, suséerna i Ham, eméerna i Save-Kirjataim
och horéerna på deras berg Seir och drevo dem ända till El-Paran vid öknen.
Sedan vände de om och kommo till En-Mispat, det är Kades, och härjade amalekiternas hela land; de slogo ock amoréerna som bodde i Hasason-Tamar.
Då drogo konungen i Sodom, konungen i Gomorra, konungen i Adma, konungen i Seboim och konungen i Bela, det är Soar, ut och ställde upp sig i Siddimsdalen till strid mot dem --
mot Kedorlaomer, konungen i Elam, Tideal, konungen över Goim, Amrafel, konungen i Sinear, och Arjok, konungen i Ellasar, fyra konungar mot de fem.
Men Siddimsdalen var full av jordbecksgropar.
Och konungarna i Sodom och Gomorra måste fly och föllo då i dessa, och de som kommo undan flydde till bergsbygden.
Så togo de allt gods som fanns i Sodom och Gomorra, och alla livsmedel där, och tågade bort;
de togo ock med sig Lot, Abrams brorson, och hans ägodelar, när de tågade bort; ty denne bodde i Sodom.
Men en av de räddade kom och berättade detta för Abram, hebréen; denne bodde vid den terebintlund som tillhörde amoréen Mamre, Eskols och Aners broder, och dessa voro i förbund med Abram.
Då nu Abram hörde att hans frände var fången, lät han sina mest beprövade tjänare, sådana som voro födda i hans hus, tre hundra aderton män, rycka ut, och förföljde fienderna ända till Dan.
Och han delade sitt folk och överföll dem så om natten med sina tjänare och slog dem, och förföljde dem sedan ända till Hoba, norr om Damaskus,
och tog tillbaka allt godset; sin frände Lot och hans ägodelar tog han ock tillbaka, ävensom kvinnorna och det övriga folket.
Då han nu var på återvägen, sedan han hade slagit Kedorlaomer och de konungar som voro på hans sida, gick konungen i Sodom honom till mötes i Savedalen, det är Konungsdalen.
Och Melki-Sedek, konungen i Salem, lät bära ut bröd och vin; denne var präst åt Gud den Högste.
Och han välsignade honom och sade: »Välsignad vare Abram av Gud den Högste, himmelens och jordens skapare!
Och välsignad vare Gud den Högste, som har givit dina ovänner i din hand!»
Och Abram gav honom tionde av allt.
Och konungen i Sodom sade till Abram: »Giv mig folket; godset må du behålla för dig själv.»
Men Abram svarade konungen i Sodom: »Jag lyfter min hand upp till HERREN, till Gud den Högste, himmelens och jordens skapare, och betygar
att jag icke vill taga ens en tråd eller en skorem, än mindre något annat som tillhör dig.
Du skall icke kunna säga: 'Jag har riktat Abram.'
Jag vill intet hava; det är nog med vad mina män hava förtärt och den del som tillkommer mina följeslagare.
Aner, Eskol och Mamre, de må få sin del.»
En tid härefter kom HERRENS ord i en syn till Abram; han sade: »Frukta icke, Abram, jag är din sköld, din lön skall bliva mycket stor.»
Men Abram sade: »Herre, HERRE, vad vill du då giva mig?
Jag går ju barnlös bort, och arvinge till mitt hus bliver en man från Damaskus, Elieser.»
Och Abram sade ytterligare: »Mig har du icke givit någon livsfrukt; en av mitt husfolk skall bliva min arvinge.»
Men se, HERRENS ord kom till honom; han sade: »Nej, denne skall icke bliva din arvinge, utan en som utgår från ditt eget liv skall bliva din arvinge.»
Och han förde honom ut och sade: »Skåda upp till himmelen, och räkna stjärnorna, om du kan räkna dem.»
Och han sade till honom: »Så skall din säd bliva.»
Och han trodde på HERREN; och han räknade honom det till rättfärdighet.
Och han sade till honom: »Jag är HERREN, som har fört dig ut från det kaldeiska Ur för att giva dig detta land till besittning.»
Han svarade: »Herre, HERRE, varav skall jag veta att jag skall besitta det?»
Då sade han till honom: »Tag åt mig en treårig kviga, en treårig get och en treårig vädur, därtill en turturduva och en ung duva.»
Och han tog åt honom alla dessa djur och styckade dem mitt itu och lade styckena mitt emot varandra; dock styckade han icke fåglarna.
Och rovfåglarna slogo ned på de döda kropparna, men Abram drev bort dem.
När nu solen var nära att gå ned och en tung sömn hade fallit på Abram, se, då kom en förskräckelse över honom och ett stort mörker.
Och han sade till Abram: »Det skall du veta, att din säd skall komma att leva såsom främlingar i ett land som icke tillhör dem, och de skola där vara trälar, och man skall förtrycka dem; så skall ske i fyra hundra år.»
Men det folk vars trälar de bliva skall jag ock döma.
Sedan skola de draga ut med stora ägodelar.
Men du själv skall gå till dina fäder i frid och bliva begraven i en god ålder.
Och i det fjärde släktet skall din säd komma hit tillbaka.
Ty ännu hava icke amoréerna fyllt sin missgärnings mått.»
Då nu solen hade gått ned och det hade blivit alldeles mörkt, syntes en rykande ugn med flammande låga, som for fram mellan styckena.
På den dagen slöt HERREN ett förbund med Abram och sade: »Åt din säd skall jag giva detta land, från Egyptens flod ända till den stora floden, till floden Frat:
kainéernas, kenaséernas, kadmonéernas,
hetiternas, perisséernas, rafaéernas,
amoréernas, kananéernas, girgaséernas och jebuséernas land.»
Och Sarai, Abrams hustru, hade icke fött barn åt honom.
Men hon hade en egyptisk tjänstekvinna, som hette Hagar;
och Sarai sade till Abram: »Se, HERREN har gjort mig ofruktsam, så att jag icke föder barn; gå in till min tjänstekvinna, kanhända skall jag få avkomma genom henne.»
Abram lyssnade till Sarais ord;
och Sarai, Abrams hustru, tog sin egyptiska tjänstekvinna Hagar och gav henne till hustru åt sin man Abram, sedan denne hade bott tio år i Kanaans land.
Och han gick in till Hagar, och hon blev havande.
När hon nu såg att hon var havande, ringaktade hon sin fru.
Då sade Sarai till Abram: »Den orätt mig sker komme över dig.
Jag själv lade min tjänstekvinna i din famn, men då hon nu ser att hon är havande, ringaktar hon mig.
HERREN döme mellan mig och dig.»
Abram sade till Sarai: »Din tjänstekvinna är ju i din hand, gör med henne vad du finner för gott.»
När då Sarai tuktade henne, flydde hon bort ifrån henne.
Men HERRENS ängel kom emot henne vid en vattenkälla i öknen, den källa som ligger vid vägen till Sur.
Och han sade: »Hagar, Sarais tjänstekvinna, varifrån kommer du, och vart går du?»
Hon svarade: »Jag är stadd på flykt ifrån min fru Sarai.»
Då sade HERRENS ängel till henne: »Vänd tillbaka till din fru, och ödmjuka dig under henne.»
Och HERRENS ängel sade till henne: »Jag skall göra din säd mycket talrik, så att man icke skall kunna räkna den för dess myckenhets skull.»
Ytterligare sade HERRENS ängel till henne: »Se, du är havande och skall föda en son; honom skall du giva namnet Ismael, därför att HERREN har hört ditt lidande.
Och han skall bliva lik en vildåsna; hans hand skall vara emot var man, och var mans hand emot honom; och han skall ligga i strid med alla sina bröder.»
Och hon gav HERREN, som hade talat med henne, ett namn, i det hon sade: »Du är Seendets Gud.»
Hon tänkte nämligen: »Har jag då verkligen här fått se en skymt av honom som ser mig ?»
Därav kallades brunnen Beer-Lahai-Roi; den ligger mellan Kades och Bered.
Och Hagar födde åt Abram en son; och Abram gav den son som Hagar hade fött åt honom namnet Ismael.
Och Abram var åttiosex år gammal, när Hagar födde Ismael åt Abram.
När Abram var nittionio år gammal, uppenbarade sig HERREN för honom och sade till honom: »Jag är Gud den Allsmäktige.
Vandra inför mig och var ostrafflig.
Jag vill göra ett förbund mellan mig och dig, och jag skall föröka dig övermåttan.»
Då föll Abram ned på sitt ansikte, och Gud talade så med honom:
»Se, det förbund som jag å min sida gör med dig är detta, att du skall bliva en fader till många folk.
Därför skall du icke mer heta Abram, utan Abraham skall vara ditt namn, ty jag skall låta dig bliva en fader till många folk.
Och jag skall göra dig övermåttan fruktsam och låta folkslag komma av dig, och konungar skola utgå från dig.
Och jag skall upprätta ett förbund mellan mig och dig och din säd efter dig, från släkte till släkte, ett evigt förbund, så att jag skall vara din Gud och din säds efter dig;
och jag skall giva dig och din säd efter dig det land där du nu bor såsom främling, hela Kanaans land, till evärdlig besittning, och jag skall vara deras Gud.
Och Gud sade ytterligare till Abraham: »Du åter skall hålla mitt förbund, du och din säd efter dig, från släkte till släkte.»
Och detta är det förbund mellan mig och eder och din säd efter dig, som I skolen hålla: allt mankön bland eder skall omskäras;
på eder förhud skolen I omskäras, och detta skall vara tecknet till förbundet mellan mig och eder.
Släkte efter släkte skall vart gossebarn bland eder omskäras, när det är åtta dagar gammalt, jämväl den hemfödde tjänaren och den som är köpt för penningar från något främmande folk, och som icke är av din säd.
Omskäras skall både din hemfödde tjänare och den som du har köpt för penningar; och så skall mitt förbund vara på edert kött betygat såsom ett evigt förbund.
Men en oomskuren av mankön, en vilkens förhud icke har blivit omskuren, han skall utrotas ur sin släkt; han har brutit mitt förbund.»
Och Gud sade åter till Abraham: »Din hustru Sarai skall du icke mer kalla Sarai, utan Sara skall vara hennes namn.
Och jag skall välsigna henne och skall också med henne giva dig en son; ja, jag skall välsigna henne, och folkslag skola komma av henne, konungar över folk skola härstamma från henne.»
Då föll Abraham ned på sitt ansikte och log, ty han sade vid sig själv: »Skulle barn födas åt en man som är hundra år gammal?
Och skulle Sara föda barn, hon som är nittio år gammal?»
Och Abraham sade till Gud: »Måtte allenast Ismael få leva inför dig!»
Då sade Gud: »Nej, din hustru Sara skall föda dig en son, och du skall giva honom namnet Isak; och med honom skall jag upprätta mitt förbund, ett evigt förbund, som skall gälla hans säd efter honom.
Men angående Ismael har jag ock hört din bön; se, jag skall välsigna honom och göra honom fruktsam och föröka honom övermåttan.
Tolv hövdingar skall han få till söner, och jag skall göra honom till ett stort folk.
Men mitt förbund skall jag upprätta med Isak, honom som Sara skall föda åt dig vid denna tid nästa år.»
Då Gud nu hade talat ut med Abraham, for han upp från honom.
Och Abraham tog sin son Ismael och alla sina tjänare, de hemfödda och de som voro köpta för penningar, allt mankön bland Abrahams husfolk, och omskar på denna samma dag deras förhud, såsom Gud hade tillsagt honom.
Och Abraham var nittionio år gammal, när hans förhud blev omskuren.
Och hans son Ismael var tretton år gammal, när hans förhud blev omskuren.
På denna samma dag omskuros Abraham och hans son Ismael;
och alla män i hans hus, de hemfödda tjänarna och de som voro köpta för penningar ifrån främmande folk, blevo omskurna tillika med honom.
Och HERREN uppenbarade sig för honom vid Mamres terebintlund, där han satt vid ingången till sitt tält, då det var som hetast på dagen.
När han lyfte upp sina ögon, fick han se tre män stå framför sig.
Och då han såg dem, skyndade han emot dem från tältets ingång och bugade sig ned till jorden
och sade: »Herre, har jag funnit nåd för dina ögon, så gå icke förbi din tjänare.
Låt mig hämta litet vatten, så att I kunnen två edra fötter; och vilen eder under trädet.
Jag vill ock hämta ett stycke bröd, så att I kunnen vederkvicka eder, innan I gån vidare, eftersom I nu haven tagit vägen förbi eder tjänare.»
De sade: »Gör såsom du har sagt.»
Och Abraham skyndade in i tältet till Sara och sade: »Skynda dig och tag tre sea-mått fint mjöl, knåda det och baka kakor.»
Men själv hastade Abraham bort till boskapen och tog en god ungkalv och gav den åt sin tjänare, och denne skyndade sig att tillreda den.
Och han tog gräddmjölk och söt mjölk och kalven, som han hade låtit tillreda, och satte fram för dem; och han stod själv hos dem under trädet, medan de åto.
Och de sade till honom: »Var är din hustru Sara?»
Han svarade: »Därinne i tältet.»
Då sade han: »Jag skall komma tillbaka till dig nästa år vid denna tid, och se, då skall din hustru Sara hava en son.»
Detta hörde Sara, där hon stod i ingången till tältet, som var bakom honom.
Men Abraham och Sara voro gamla och komna till hög ålder, och Sara hade icke mer, såsom kvinnor pläga hava.
Därför log Sara vid sig själv och tänkte: »Skulle jag väl nu på min ålderdom giva mig till lusta, nu då också min herre är gammal?»
Men HERREN sade till Abraham: »Varför log Sara och tänkte: 'Skulle jag verkligen föda barn, så gammal som jag är?'
Är då något så underbart, att HERREN icke skulle förmå det?
På den bestämda tiden skall jag komma tillbaka till dig, vid denna tid nästa år, och då skall Sara hava en son.»
Då nekade Sara och sade: »Jag log icke»; ty hon blev förskräckt.
Men han sade: »Jo, du log.»
Och männen stodo upp för att gå därifrån och vände sina blickar ned mot Sodom, och Abraham gick med för att ledsaga dem.
Och HERREN sade: »Kan jag väl dölja för Abraham vad jag tänker göra?
Av Abraham skall ju bliva ett stort och mäktigt folk, och i honom skola alla folk på jorden varda välsignade.
Ty därtill har jag utvalt honom, för att han skall bjuda sina barn och sitt hus efter sig att hålla HERRENS väg och öva rättfärdighet och rätt, på det att HERREN må låta det komma över Abraham, som han har lovat honom.»
Och HERREN sade: »Ropet från Sodom och Gomorra är stort, och deras synd är mycket svår;
därför vill jag gå ditned och se om de verkligen i allt hava gjort efter det rop som har kommit till mig; om så icke är, vill jag veta det.»
Och männen begåvo sig därifrån och gingo mot Sodom; men Abraham stod ännu kvar inför HERREN.
Och Abraham trädde närmare och sade: »Vill du då förgöra den rättfärdige tillika med den ogudaktige?
Kanhända finnas femtio rättfärdiga i staden; vill du då förgöra den och icke skona orten för de femtio rättfärdigas skull som finnas där?
Bort det, att du skulle så göra och döda den rättfärdige tillika med den ogudaktige, så att det skulle gå den rättfärdige likasom den ogudaktige; bort det ifrån dig!
Skulle han som är hela jordens domare icke göra vad rätt är?»
HERREN sade: »Om jag i Sodom finner femtio rättfärdiga inom staden, så vill jag skona orten för deras skull.»
Men Abraham svarade och sade: »Se, jag har dristat mig att tala till Herren, fastän jag är stoft och aska.»
Kanhända skall det fattas fem i de femtio rättfärdiga; vill du då för de fems skull fördärva hela staden?»
Han sade: »Om jag där finner fyrtiofem; så skall jag icke fördärva den.»
Men han fortfor att tala till honom och sade: »Kanhända skola fyrtio finnas där.»
Han svarade: »Jag skall då icke göra det, för de fyrtios skull.»
Då sade han: »Herre, vredgas icke över att jag ännu talar något.
Kanhända skola trettio finnas där.»
Han svarade: »Om jag där finner trettio, så skall jag icke göra det.»
Men han sade: »Se, jag har dristat mig att tala till Herren.
Kanhända skola tjugu finnas där.»
Han svarade: »Jag skall då icke fördärva den, för de tjugus skull.»
Då sade han: »Herre, vredgas icke över att jag talar allenast ännu en gång.
Kanhända skola tio finnas där.»
Han svarade: »Jag skall då icke fördärva den, för de tios skull.»
Och HERREN gick bort, sedan han hade talat ut med Abraham; och Abraham vände tillbaka hem.
Och de två änglarna kommo om aftonen till Sodom, och Lot satt då i Sodoms port.
När Lot fick se dem, stod han upp och gick emot dem och föll ned till jorden på sitt ansikte
och sade: »I herrar, tagen härbärge i eder tjänares hus och stannen där över natten, och tvån edra fötter; sedan kunnen I i morgon bittida fortsätta eder färd.»
De svarade: »Nej, vi vilja stanna på gatan över natten.»
Men han bad dem så enträget, att de togo härbärge hos honom och kommo in i hans hus.
Och han tillredde en måltid åt dem och bakade osyrat bröd, och de åto.
Men innan de hade lagt sig, omringades huset av männen i staden, Sodoms män, både unga och gamla, allt folket, så många de voro.
Dessa kallade på Lot och sade till honom: »Var äro de män som hava kommit till dig i natt?
För dem ut till oss, så att vi få känna dem.»
Då gick Lot ut till dem i porten och stängde dörren efter sig
och sade: »Mina bröder, gören icke så illa.
Se, jag har två döttrar, som ännu icke veta av någon man.
Dem vill jag föra ut till eder, så kunnen I göra med dem vad I finnen för gott.
Gören allenast icke något mot dessa män, eftersom de nu hava gått in under skuggan av mitt tak.»
Men de svarade: »Bort med dig!»
Och de sade ytterligare: »Denne, en ensam man, har kommit hit och bor här såsom främling, och han vill dock ständigt upphäva sig som domare.
Men nu skola vi göra dig mer ont än dem.»
Och de trängde med våld in på mannen Lot och stormade fram för att spränga dörren.
Då räckte männen ut sina händer och togo Lot in till sig i huset och stängde dörren.
Och de män som stodo utanför husets port slogo de med blindhet, både små och stora, så att de förgäves sökte finna porten.
Och männen sade till Lot: »Har du någon mer här, någon måg, eller några söner eller döttrar, eller någon annan som tillhör dig i staden, så för dem bort ifrån detta ställe.
Ty vi skola fördärva detta ställe; ropet från dem har blivit så stort inför HERREN, att HERREN har utsänt oss till att fördärva dem.»
Då gick Lot ut och talade till sina mågar, som skulle få hans döttrar, och sade: »Stån upp och gån bort ifrån detta ställe; ty HERREN skall fördärva staden.»
Men hans mågar menade att han skämtade.
När nu morgonrodnaden gick upp, manade änglarna på Lot och sade: »Stå upp och tag med dig din hustru och dina båda döttrar, som du har hos dig, på det att du icke må förgås genom stadens missgärning.»
Och då han ännu dröjde, togo männen honom vid handen jämte hans hustru och hans båda döttrar, ty HERREN ville skona honom; och de förde honom ut, och när de voro utanför staden, släppte de honom.
Och medan de förde dem ut, sade den ene: »Fly för ditt livs skull; se dig icke tillbaka, och dröj ingenstädes på Slätten.
Fly undan till bergen, så att du icke förgås.»
Men Lot sade till dem: »Ack nej, Herre.
Se, din tjänare har ju funnit nåd för dina ögon, och stor är den barmhärtighet som du gör med mig, då du vill rädda mitt liv; men jag förmår icke fly undan till bergen; jag rädes att olyckan hinner mig, så att jag omkommer.
Se, staden därborta ligger helt nära, och det är lätt att fly dit, och den är liten; låt mig fly undan dit -- den är ju så liten -- på det att jag må bliva vid liv.»
Då svarade han honom: »Välan, jag skall ock häri göra dig till viljes; jag skall icke omstörta den stad som du talar om.
Men skynda att fly undan dit; ty jag kan intet göra, förrän du har kommit dit.»
Därav fick staden namnet Soar .
Då nu solen hade gått upp över jorden och Lot hade kommit till Soar,
lät HERREN svavel och eld regna från himmelen, från HERREN, över Sodom och Gomorra;
och han omstörtade dessa städer med hela Slätten och alla dem som bodde i städerna och det som växte på marken.
Och Lots hustru, som följde efter honom, såg sig tillbaka; då blev hon en saltstod.
Och när Abraham bittida följande morgon gick till den plats där han hade stått inför HERREN,
och blickade ned över Sodom och Gomorra och över hela Slättlandet, då fick han se en rök stiga upp från landet, lik röken från en smältugn.
Så skedde då, att när Gud fördärvade städerna på Slätten, tänkte han på Abraham och lät Lot komma undan omstörtningen, då han omstörtade städerna där Lot hade bott.
Och Lot drog upp från Soar till bergsbygden och bodde där med sina båda döttrar, ty han fruktade för att bo kvar i Soar; och han bodde med sina båda döttrar i en grotta.
Då sade den äldre till den yngre: »Vår fader är gammal, och ingen man finnes i landet, som kan gå in till oss efter all världens sedvänja.
Kom, låt oss giva vår fader vin att dricka och lägga oss hos honom, för att vi må skaffa oss livsfrukt genom vår fader.»
Så gåvo de sin fader vin att dricka den natten, och den äldre gick in och lade sig hos sin fader, och han märkte icke när hon lade sig, ej heller när hon stod upp.
Dagen därefter sade den äldre till den yngre: »Se, jag låg i natt hos min fader; låt oss också denna natt giva honom vin att dricka, och gå du in och lägg dig hos honom, för att vi må skaffa oss livsfrukt genom vår fader.»
Så gåvo de också den natten sin fader vin att dricka; och den yngre gick och lade sig hos honom, och han märkte icke när hon lade sig, ej heller när hon stod upp.
Så blevo Lots båda döttrar havande genom sin fader.
Och den äldre födde en son, och hon gav honom namnet Moab; från honom härstamma moabiterna ända till denna dag.
Den yngre födde ock en son, och hon gav honom namnet Ben-Ammi; från honom härstamma Ammons barn ända till denna dag.
Och Abraham bröt upp därifrån och drog till Sydlandet; där uppehöll han sig mellan Kades och Sur, och någon tid bodde han i Gerar.
Och Abraham sade om sin hustru Sara att hon var hans syster.
Då sände Abimelek, konungen i Gerar, och lät hämta Sara till sig.
Men Gud kom till Abimelek i en dröm om natten och sade till honom: »Se, du måste dö för den kvinnas skull som du har tagit till dig, fast hon är en annan mans äkta hustru.»
Men Abimelek hade icke kommit vid henne.
Och han svarade: »Herre, vill du då dräpa också rättfärdiga människor?
Sade han icke själv till mig: 'Hon är min syster'?
Och likaså sade hon: 'Han är min broder.'
I mitt hjärtas oskuld och med rena händer har jag gjort detta.»
Då sade Gud till honom i drömmen: »Ja, jag vet att du har gjort detta i ditt hjärtas oskuld, och jag har själv hindrat dig från att synda mot mig; därför har jag icke tillstatt dig att komma vid henne.
Men giv nu mannen hans hustru tillbaka; ty han är en profet.
Och han må bedja för dig, så att du får leva.
Men om du icke giver henne tillbaka, så vet att du skall döden dö, du själv och alla som tillhöra dig.
Då stod Abimelek upp bittida om morgonen och kallade till sig alla sina tjänare och berättade allt detta för dem; och männen blevo mycket förskräckta.
Sedan kallade Abimelek Abraham till sig och sade till honom: »Vad har du gjort mot oss!
Vari har jag försyndat mig mot dig, eftersom du har velat komma mig och mitt rike att begå en så stor synd?
På otillbörligt sätt har du handlat mot mig.»
Och Abimelek sade ytterligare till Abraham: »Vad var din mening, när du gjorde detta?»
Abraham svarade: »Jag tänkte: 'På denna ort fruktar man nog icke Gud; de skola dräpa mig för min hustrus skull.'
Hon är också verkligen min syster, min faders dotter, fastän icke min moders dotter; och så blev hon min hustru.
Men när Gud sände mig ut på vandring bort ifrån min faders hus, sade jag till henne: 'Bevisa mig din kärlek därmed att du säger om mig, varthelst vi komma, att jag är din broder.'»
Då tog Abimelek får och fäkreatur, tjänare och tjänarinnor och gav dem åt Abraham.
Han gav honom ock hans hustru Sara tillbaka.
Och Abimelek sade: »Se, mitt land ligger öppet för dig; du må bo var du finner för gott.»
Och till Sara sade han: »Se, jag giver åt din broder tusen siklar silver; det skall för dig vara en försoningsgåva inför allt ditt folk.
Så har du inför alla fått upprättelse.»
Och Abraham bad till Gud, och Gud botade Abimelek och hans hustru och hans tjänstekvinnor, så att de åter kunde föda barn.
HERREN hade nämligen gjort alla kvinnor i Abimeleks hus ofruktsamma, för Saras, Abrahams hustrus, skull.
Och HERREN såg till Sara, såsom han hade lovat, och HERREN gjorde med Sara såsom han hade sagt.
Sara blev havande och födde åt Abraham en son på hans ålderdom, vid den bestämda tid som Gud hade sagt honom.
Och Abraham gav den son som var född åt honom, den som Sara hade fött åt honom, namnet Isak.
Och Abraham omskar sin son Isak, när denne var åtta dagar gammal, såsom Gud hade bjudit honom.
Och Abraham var hundra år gammal, när hans son Isak föddes åt honom.
Och Sara sade: »Gud har berett mig ett löje; var och en som får höra detta skall le mot mig.»
Och hon sade: »Vem skulle hava sagt Abraham att Sara skulle giva barn di?
Och nu har jag fött honom en son på hans ålderdom!»
Och barnet växte upp och blev avvant; och den dag då Isak avvandes gjorde Abraham ett stort gästabud.
Då fick Sara se Hagars, den egyptiska kvinnans, son, som denna hade fött åt Abraham, leka och skämta;
och hon sade till Abraham: »Driv ut denna tjänstekvinna och hennes son, ty denna tjänstekvinnas son skall icke ärva med min son Isak.»
Det talet misshagade Abraham mycket för hans sons skull.
Men Gud sade till Abraham: »Du må icke för gossens och för din tjänstekvinnas skull låta detta misshaga dig.
Lyssna till Sara i allt vad hon säger dig; ty genom Isak är det som säd skall uppkallas efter dig.
Men också tjänstekvinnans son skall jag göra till ett folk, därför att han är din säd.»
Bittida följande morgon tog Abraham bröd och en lägel med vatten och gav det åt Hagar; han lade det på hennes rygg och gav henne barnet med och lät henne gå.
Och hon begav sig åstad och irrade omkring i Beer-Sebas öken.
Men när vattnet i lägeln hade tagit slut, kastade hon barnet ifrån sig under en buske
och gick bort och satte sig ett stycke därifrån, på ett bågskotts avstånd, ty hon tänkte: »Jag förmår icke se på, huru barnet dör.»
Och där hon nu satt, på något avstånd, brast hon ut i gråt.
Då hörde Gud gossens röst, och Guds ängel ropade till Hagar från himmelen och sade till henne: »Vad fattas dig, Hagar?
Frukta icke; ty Gud har hört gossens röst, där han ligger.
Gå och lyft upp gossen, och tag honom vid handen; jag skall göra honom till ett stort folk.»
Och Gud öppnade hennes ögon, så att hon blev varse en vattenbrunn.
Och hon gick dit och fyllde sin lägel med vatten och gav gossen att dricka.
Och Gud var med gossen, och han växte upp och bodde i öknen och blev med tiden en bågskytt.
Han bodde i öknen Paran; och hans moder tog en hustru åt honom från Egyptens land.
Vid den tiden kom Abimelek med Pikol, sin härhövitsman, och talade med Abraham och sade: »Gud är med dig i allt vad du gör.
Så lova mig nu här med ed vid Gud att du icke skall göra dig skyldig till något svek mot mig eller mina barn och efterkommande, utan att du skall bevisa mig och det land där du nu bor såsom främling samma godhet som jag har bevisat dig.»
Abraham sade: »Det vill jag lova dig.»
Dock gjorde Abraham Abimelek förebråelser angående en vattenbrunn som Abimeleks tjänare hade tagit ifrån honom.
Men Abimelek svarade: »Jag vet icke vem som har gjort detta; själv har du ingenting sagt mig, och jag har icke hört något därom förrän i dag.»
Då tog Abraham får och fäkreatur och gav åt Abimelek; och de slöto förbund med varandra.
Men Abraham ställde sju lamm av hjorden avsides.
Då sade Abimelek till Abraham: »Vad betyda de sju lammen som du har ställt där avsides?»
Han svarade: »Dessa sju lamm skall du taga emot av mig, för att detta må vara mig till ett vittnesbörd därom att det är jag som har grävt denna brunn.»
Därav kallades det stället Beer-Seba , eftersom de båda där gingo eden.
När de så hade slutit förbund vid Beer-Seba, stodo Abimelek och hans härhövitsman Pikol upp och vände tillbaka till filistéernas land.
Och Abraham planterade en tamarisk vid Beer-Seba och åkallade där HERRENS, den evige Gudens, namn.
Och Abraham bodde i filistéernas land en lång tid.
En tid härefter hände sig att Gud satte Abraham på prov.
Han sade till honom: »Abraham!»
Han svarade: »Här är jag.»
Då sade han: »Tag din son Isak, din ende son, som du har kär, och gå bort till Moria land, och offra honom där såsom brännoffer, på ett berg som jag skall säga dig.»
Bittida följande morgon lastade Abraham sin åsna och tog med sig två sina tjänare och sin son Isak; och sedan han hade huggit sönder ved till brännoffer, bröt han upp och begav sig på väg till den plats som Gud hade sagt honom.
När nu Abraham på tredje dagen lyfte upp sina ögon och fick se platsen på avstånd,
sade han till sina tjänare: »Stannen I här med åsnan; jag och gossen vilja gå ditbort.
När vi hava tillbett, skola vi komma tillbaka till eder.»
Och Abraham tog veden till brännoffret och lade den på sin son Isak, men själv tog han elden och kniven, och de gingo så båda tillsammans.
Då talade Isak till sin fader Abraham och sade: »Min fader!»
Han svarade: »Vad vill du, min son?»
Han sade: »Se, här är elden och veden, men var är fåret till brännoffret?»
Abraham svarade: »Gud utser nog åt sig fåret till brännoffret, min son.»
Så gingo de båda tillsammans.
När de nu hade kommit till den plats som Gud hade sagt Abraham, byggde han där ett altare och lade veden därpå, sedan band han sin son Isak och lade honom på altaret ovanpå veden.
Och Abraham räckte ut sin hand och tog kniven för att slakta sin son.
Då ropade HERRENS ängel till honom från himmelen och sade: »Abraham!
Abraham!»
Han svarade: »Här är jag.»
Då sade han: »Låt icke din hand komma vid gossen, och gör honom intet; ty nu vet jag att du fruktar Gud, nu då du icke har undanhållit mig din ende son.»
När då Abraham lyfte upp sina ögon, fick han bakom sig se en vädur, som hade fastnat med sina horn i ett snår; och Abraham gick dit och tog väduren och offrade den till brännoffer i sin sons ställe.
Och Abraham gav den platsen namnet HERREN utser ; nu för tiden heter den Berget där HERREN låter se sig .
Och HERRENS ängel ropade för andra gången till Abraham från himmelen
och sade: »Jag svär vid mig själv, säger HERREN: Eftersom du har gjort detta och icke undanhållit mig din ende son
därför skall jag rikligen välsigna dig och göra din säd talrik såsom stjärnorna på himmelen och såsom sanden på havets strand; och din säd skall intaga sina fienders portar.
Och i din säd skola alla folk på jorden välsigna sig, därför att du lyssnade till mina ord.»
Sedan vände Abraham tillbaka till sina tjänare; och de stodo upp och gingo tillsammans till Beer-Seba.
Och Abraham bodde i Beer-Seba.
En tid härefter blev så berättat för Abraham: »Se, Milka har ock fött barn åt din broder Nahor.»
Barnen voro Us, hans förstfödde, och Bus, dennes broder, och Kemuel, Arams fader,
vidare Kesed, Haso, Pildas, Jidlaf och Betuel.
Men Betuel födde Rebecka.
Dessa åtta föddes av Milka åt Nahor, Abrahams broder.
Och hans bihustru, som hette Reuma, födde ock barn, nämligen Teba, Gaham, Tahas och Maaka.
Och Sara blev ett hundra tjugusju år gammal; så gammal blev Sara.
Och Sara dog i Kirjat-Arba, det är Hebron, i Kanaans land.
Och Abraham kom och höll dödsklagan efter Sara och begrät henne.
Därefter stod Abraham upp och gick bort ifrån den döda och talade så till Hets barn:
»Jag är en främling och gäst hos eder.
Låten mig nu få en egen grav hos eder, så att jag kan föra min döda dit och begrava henne.»
Då svarade Hets barn Abraham och sade till honom:
»Hör oss, herre.
Du är en Guds hövding bland oss; begrav din döda i den förnämligaste av våra gravar.
Ingen av oss skall vägra att giva dig sin grav till att där begrava din döda.»
Men Abraham stod upp och bugade sig för landets folk, Hets barn;
och han talade med dem och sade: »Om I tillstädjen att jag för ut min döda och begraver henne, så hören mig och läggen eder ut för mig hos Efron, Sohars son,
så att han giver mig den grotta i Makpela, som tillhör honom, och som ligger vid ändan av hans åker.
Mot full betalning i eder krets må han giva mig den till egen grav.»
Men Efron satt där bland Hets barn.
Och Efron, hetiten, svarade Abraham i närvaro av Hets barn, alla som bodde inom hans stadsport; han sade:
»Icke så, min herre.
Hör mig: Jag skänker dig åkern; grottan som finnes där skänker jag dig ock; jag skänker dig den inför mina landsmäns ögon; begrav där din döda.»
Men Abraham bugade sig för landets folk;
och han talade till Efron i närvaro av landets folk och sade: »Värdes dock höra mig.
Jag vill betala åkerns värde; tag emot det av mig, och låt mig där begrava min döda.»
Då svarade Efron Abraham och sade till honom:
»Min herre, hör mig.
Ett jordstycke till ett värde av fyra hundra siklar silver, vad betyder det mellan mig och dig?
Begrav du din döda.»
Och Abraham förstod Efron och vägde upp åt honom den summa som Efron hade uppgivit i närvaro av Hets barn, fyra hundra siklar silver, sådant silver som var gångbart i handel.
Så skedde det att Efrons åker i Makpela, gent emot Mamre, själva åkern med grottan som fanns där och alla träd på åkern, så långt dess område sträckte sig runt omkring, blev överlåten åt Abraham till egendom
inför Hets barns ögon, inför alla som bodde inom hans stadsport.
Därefter begrov Abraham sin hustru Sara i grottan på åkern i Makpela, gent emot Mamre, det är Hebron, i Kanaans land.
Åkern med grottan som fanns där blev så av Hets barn överlåten åt Abraham till egen grav.
Abraham var nu gammal och kommen till hög ålder, och HERREN hade välsignat Abraham i alla stycken.
Då sade han till sin äldste hustjänare, den som förestod all hans egendom: »Lägg din hand under min länd;
jag vill av dig taga en ed vid HERREN, himmelens Gud och jordens Gud, att du icke till hustru åt min son skall taga en dotter till någon av kananéerna bland vilka jag bor,
utan att du skall gå till mitt eget land och till min släkt och där taga hustru åt min son Isak.»
Tjänaren sade till honom: »Men om så händer, att kvinnan icke vill följa mig hit till landet, måste jag då föra din son tillbaka till det land som du har kommit ifrån?»
Abraham svarade honom: »Tag dig till vara för att föra min son dit tillbaka.
HERREN, himmelens Gud, som har fört mig bort ifrån min faders hus och ifrån mitt fädernesland, han som har talat till mig och svurit och sagt: 'Åt din säd skall jag giva detta land', han skall sända sin ängel framför dig, så att du därifrån skall kunna få en hustru åt min son.
Men om kvinnan icke vill följa dig, så är du fri ifrån denna din ed till mig.
Allenast må du icke föra min son dit tillbaka.»
Då lade tjänaren sin hand under sin herre Abrahams länd och lovade honom detta med ed.
Och tjänaren tog tio av sin herres kameler och drog åstad med allahanda dyrbara gåvor från sin herre; han stod upp och drog åstad till Nahors stad i Aram-Naharaim.
Där lät han kamelerna lägra sig utanför staden, vid en vattenbrunn; och det led mot aftonen, den tid då kvinnorna plägade komma ut för att hämta vatten.
Och han sade: »HERRE, min herre Abrahams Gud, låt mig i dag få ett lyckosamt möte, och gör nåd med min herre Abraham.
Se, jag står här vid vattenkällan, och stadsbornas döttrar komma hitut för att hämta vatten.
Om jag nu säger till en flicka: 'Håll hit din kruka, och låt mig få dricka' och hon då svarar: 'Drick; dina kameler vill jag ock vattna', må hon då vara den som du har utsett åt din tjänare Isak, så skall jag därav veta att du har gjort nåd med min herre.»
Och se, innan han hade slutat att tala, kom Rebecka ditut, en dotter till Betuel, som var son till Milka, Abrahams broder Nahors hustru; och hon bar sin kruka på axeln.
Och flickan var mycket fager att skåda, en jungfru som ingen man hade känt.
Hon gick nu ned till källan och fyllde sin kruka och steg så upp igen.
Då skyndade tjänaren emot henne och sade: »Låt mig få dricka litet vatten ur din kruka.»
Hon svarade: »Drick, min herre» och lyfte strax ned krukan på sin hand och gav honom att dricka.
Och sedan hon hade givit honom att dricka, sade hon: »Jag vill ock ösa upp vatten åt dina kameler, till dess att de alla hava fått dricka.»
Och hon tömde strax sin kruka i vattenhon och skyndade åter till brunnen för att hämta vatten och öste så upp åt alla hans kameler.
Men mannen såg på henne under tystnad och undrade om HERREN hade gjort hans resa lyckosam eller icke.
Och när alla kamelerna hade druckit, tog mannen fram en näsring av guld, en halv sikel i vikt, och två armband av guld, tio siklar i vikt,
och frågade: »Vems dotter är du?
Säg mig det.
Och säg mig om vi kunna få natthärbärge i din faders hus?»
Hon svarade honom: »Jag är dotter till Betuel, Milkas son, som av henne föddes åt Nahor.»
Och hon sade ytterligare till honom: »Vi hava rikligt med både halm och foder; natthärbärge kan du ock få.»
Då böjde mannen sig ned och tillbad HERREN
och sade: »Lovad vare HERREN, min herre Abrahams Gud, som icke har tagit sin nåd och trofasthet ifrån min herre!
Mig har HERREN ledsagat på vägen, hem till min herres fränder.»
Och flickan skyndade åstad och berättade allt detta i sin moders hus.
Men Rebecka hade en broder som hette Laban.
Och Laban skyndade åstad till mannen därute vid källan.
När han nämligen såg näsringen och armbanden som hans syster bar, och när han hörde huru hans syster Rebecka berättade: 'Så och så talade mannen till mig', då begav han sig ut till mannen, där denne stod hos kamelerna vid källan.
Och han sade: »Kom in, du HERRENS välsignade; varför står du härute?
Jag har berett plats i huset, och rum finnes för kamelerna.»
Så kom då mannen in i huset; och man lastade av kamelerna, och tog fram halm och foder åt kamelerna, och vatten till att två hans och hans följeslagares fötter.
Och man satte fram mat för honom; men han sade: »Jag vill icke äta, förrän jag har framfört mitt ärende.»
Laban svarade: »Så tala då.»
Då sade han: »Jag är Abrahams tjänare.
Och HERREN har rikligen välsignat min herre, så att han har blivit en mäktig man; han har givit honom får och fäkreatur, silver och guld, tjänare och tjänarinnor, kameler och åsnor.
Och Sara, min herres hustru, har fött åt min herre en son på sin ålderdom, och åt denne har han givit allt vad han äger.
Och min herre har tagit en ed av mig och sagt: 'Till hustru åt min son skall du icke taga en dotter till någon av kananéerna i vilkas land jag bor,
utan du skall gå till min faders hus och till min släkt och där taga hustru åt min son.'
Då sade jag till min herre: 'Men om nu kvinnan icke vill följa med mig?'
Han svarade mig: 'HERREN, inför vilken jag har vandrat, skall sända sin ängel med dig och göra din resa lyckosam, så att du åt min son får en hustru av min släkt och av min faders hus;
i sådant fall skall du vara löst från din ed till mig, när du har kommit till min släkt.
Också om de icke giva henne åt dig, skall du vara fri ifrån eden till mig.'
Så kom jag i dag till källan, och jag sade: HERRE, min herre Abrahams Gud, om du vill låta den resa på vilken jag är stadd bliva lyckosam,
må det då ske, när jag nu står här vid vattenkällan, att om en ung kvinna kommer ut för att hämta vatten och jag säger till henne: 'Låt mig få dricka litet vatten ur din kruka'
och hon då svarar mig: 'Drick du; åt dina kameler vill jag ock ösa upp vatten' -- må hon då vara den kvinna som HERREN har utsett åt min herres son.
Och innan jag hade slutat att så tala för mig själv, se, då kom Rebecka ut med sin kruka på axeln och gick ned till källan för att hämta vatten.
Då sade jag till henne: 'Låt mig få dricka.'
Och strax lyfte hon ned sin kruka från axeln och sade: 'Drick; dina kameler vill jag ock vattna.'
Så drack jag, och hon vattnade också kamelerna.
Och jag frågade henne och sade: 'Vems dotter är du?'
Hon svarade: 'Jag är dotter till Betuel, Nahors son, som föddes åt honom av Milka.'
Då satte jag ringen i hennes näsa och armbanden på hennes armar.
Och jag böjde mig ned och tillbad HERREN och lovade HERREN, min herre Abrahams Gud, som hade ledsagat mig på den rätta vägen, så att jag åt hans son skulle få min herres frändes dotter.
Om I nu viljen visa min herre kärlek och trofasthet, så sägen mig det; varom icke, så sägen mig ock det, för att jag då må vända mig åt annat håll, till höger eller till vänster.»
Då svarade Laban och Betuel och sade: »Från HERREN har detta utgått; vi kunna i den saken intet säga till dig, varken ont eller gott.
Se, där står Rebecka inför dig, tag henne och drag åstad; må hon bliva hustru åt din herres son, såsom HERREN har sagt.»
När Abrahams tjänare hörde deras ord, föll han ned på jorden och tillbad HERREN.
Sedan tog tjänaren fram smycken av silver och guld, så ock kläder, och gav detta åt Rebecka.
Jämväl åt hennes broder och hennes moder gav han dyrbara skänker.
Och de åto och drucko, han och hans följeslagare, och stannade sedan där över natten.
Men om morgonen, när de hade stått upp, sade han: »Låten mig nu fara till min herre.»
Då sade hennes broder och hennes moder: »Låt flickan stanna hos oss några dagar, tio eller så; sedan må du fara.»
Men han svarade dem: »Uppehållen mig icke, eftersom HERREN har gjort min resa lyckosam.
Låten mig fara; jag vill resa hem till min herre.»
Då sade de: »Vi vilja kalla hit flickan och fråga henne själv.»
Och de kallade Rebecka till sig och sade till henne: »Vill du resa med denne man?»
Hon svarade: »Ja.»
Då bestämde de att deras syster Rebecka jämte sin amma skulle fara med Abrahams tjänare och dennes män.
Och de välsignade Rebecka och sade till henne: »Av dig, du vår syster, komme tusen gånger tio tusen, och må dina avkomlingar intaga sina fienders portar.»
Och Rebecka och hennes tärnor stodo upp och satte sig på kamelerna och följde med mannen; så tog tjänaren Rebecka med sig och for sin väg.
Men Isak var på väg hem från Beer-Lahai-Roi, ty han bodde i Sydlandet.
Och mot aftonen hade Isak gått ut på fältet i sorgsna tankar.
När han då lyfte upp sina ögon, fick han se kameler komma.
Då nu också Rebecka lyfte upp sina ögon och fick se Isak, steg hon med hast ned från kamelen;
och hon frågade tjänaren: »Vem är den mannen som kommer emot oss där på fältet?»
Tjänaren svarade: »Det är min herre.»
Då tog hon sin slöja och höljde sig i den.
Och tjänaren förtäljde för Isak huru han hade uträttat allt.
Och Isak förde henne in i sin moder Saras tält; och han tog Rebecka till sig, och hon blev hans hustru, och han hade henne kär.
Så blev Isak tröstad i sorgen efter sin moder.
Och Abraham tog sig ännu en hustru, och hon hette Ketura.
Hon födde åt honom Simran, Joksan, Medan, Midjan, Jisbak och Sua.
Och Joksan födde Saba och Dedan, och Dedans söner voro assuréerna, letuséerna och leumméerna.
Och Midjans söner voro Efa, Efer, Hanok, Abida och Eldaa.
Alla dessa voro Keturas söner.
Och Abraham gav allt vad han ägde åt Isak.
Men åt sönerna till sina bihustrur gav Abraham skänker och skilde dem, medan han själv ännu levde, från sin son Isak och lät dem draga österut, bort till Österlandet.
Och detta är antalet av Abrahams levnadsår: ett hundra sjuttiofem år;
därefter gav Abraham upp andan och dog i en god ålder, gammal och mätt på livet, och blev samlad till sina fäder.
Och hans söner Isak och Ismael begrovo honom i grottan i Makpela, på hetiten Efrons, Sohars sons, åker gent emot Mamre,
den åker som Abraham hade köpt av Hets barn; där blev Abraham begraven, såväl som hans hustru Sara.
Och efter Abrahams död välsignade Gud hans son Isak.
Och Isak bodde vid Beer-Lahai-Roi.
Och detta är berättelsen om Ismaels släkt, Abrahams sons, som föddes åt Abraham av Hagar, Saras egyptiska tjänstekvinna.
Dessa äro namnen på Ismaels söner, med deras namn, efter deras ättföljd: Nebajot, Ismaels förstfödde, vidare Kedar, Adbeel, Mibsam,
Misma, Duma och Massa,
Hadad och Tema, Jetur, Nafis och Kedma.
Dessa voro Ismaels söner och dessa deras namn, i deras byar och tältläger, tolv hövdingar efter deras stammar.
Och detta är antalet av Ismaels levnadsår: ett hundra trettiosju år; därefter gav han upp andan och dog och blev samlad till sina fäder.
Och de hade sina boningsplatser från Havila ända till Sur, som ligger gent emot Egypten, fram emot Assyrien.
Han kom i strid med alla sina bröder.
Och detta är berättelsen om Isaks, Abrahams sons, släkt.
Abraham födde Isak;
och Isak var fyrtio år gammal, när han till hustru åt sig tog Rebecka, som var dotter till araméen Betuel från Paddan-Aram och syster till araméen Laban.
Och Isak bad till HERREN för sin hustru Rebecka, ty hon var ofruktsam; och HERREN bönhörde honom, så att hans hustru Rebecka blev havande.
Men barnen stötte varandra i hennes liv; då sade hon: »Om det skulle gå så, varför skulle jag då vara till?»
Och hon gick bort för att fråga HERREN.
Och HERREN svarade henne: »Två folk finnas i ditt liv, två folkstammar skola ur ditt sköte söndras från varandra; den ena stammen skall vara den andra övermäktig, och den äldre skall tjäna den yngre.»
När sedan tiden var inne att hon skulle föda, se, då funnos tvillingar i hennes liv.
Den som först kom fram var rödlätt och över hela kroppen såsom en hårmantel; och de gåvo honom namnet Esau.
Därefter kom hans broder fram, och denne höll med sin hand i Esaus häl; och han fick namnet Jakob.
Men Isak var sextio år gammal, när de föddes.
Och barnen växte upp, och Esau blev en skicklig jägare, som höll sig ute på marken; Jakob åter blev en fromsint man, som bodde i tält.
Och Isak hade Esau kärast, ty han hade smak för villebråd; men Rebecka hade Jakob kärast.
En gång, då Jakob höll på att koka något till soppa, kom Esau hem från marken, uppgiven av hunger.
Och Esau sade till Jakob: »Låt mig få till livs av det röda, det röda du har där; ty jag är uppgiven av hunger.»
Därav fick han namnet Edom .
Men Jakob sade: »Sälj då nu åt mig din förstfödslorätt.»
Esau svarade: »Jag är ju döden nära; vartill gagnar mig då min förstfödslorätt?»
Jakob sade: »Så giv mig nu din ed därpå.»
Och han gav honom sin ed och sålde så sin förstfödslorätt till Jakob.
Men Jakob gav Esau bröd och linssoppa; och han åt och drack och stod sedan upp och gick sin väg.
Så ringa aktade Esau sin förstfödslorätt.
Men en hungersnöd uppstod i landet, en ny hungersnöd, efter den som hade varit förut, i Abrahams tid.
Då begav sig Isak till Abimelek, filistéernas konung, i Gerar.
Och HERREN uppenbarade sig för honom och sade: »Drag icke ned till Egypten; bo kvar i det land som jag skall säga dig.
Stanna såsom främling här i landet; jag skall vara med dig och välsigna dig, ty åt dig och din säd skall jag giva alla dessa länder, och skall hålla den ed som jag har svurit din fader Abraham.
Jag skall göra din säd talrik såsom stjärnorna på himmelen, och jag skall giva åt din säd alla dessa länder; och i din säd skola alla folk på jorden välsigna sig,
därför att Abraham har lyssnat till mina ord och hållit vad jag har bjudit honom hålla, mina bud, mina stadgar och mina lagar.»
Så stannade Isak kvar i Gerar.
Och när männen på orten frågade honom om hans hustru, sade han: »Hon är min syster.»
Han fruktade nämligen för att säga att hon var hans hustru, ty han tänkte: »Männen här på orten kunde då dräpa mig för Rebeckas skull, eftersom hon är så fager att skåda.»
Men när han hade varit där en längre tid, hände sig en gång, då Abimelek, filistéernas konung, blickade ut genom fönstret, att han fick se Isak kärligt skämta med sin hustru Rebecka.
Då kallade Abimelek Isak till sig och sade: »Hon är ju din hustru; huru har du då kunnat säga: 'Hon är min syster'?»
Isak svarade honom: »Jag fruktade att jag annars skulle bliva dödad för hennes skull.»
Då sade Abimelek: »Vad har du gjort mot oss!
Huru lätt kunde det icke hava skett att någon av folket hade lägrat din hustru?
Och så hade du dragit skuld över oss.»
Sedan bjöd Abimelek allt folket och sade: »Den som kommer vid denne man eller vid hans hustru, han skall straffas med döden.»
Och Isak sådde där i landet och fick det året hundrafalt, ty HERREN välsignade honom.
Och han blev en mäktig man; hans makt blev större och större, så att han till slut var mycket mäktig.
Han ägde så många får och fäkreatur och så många tjänare, att filistéerna begynte avundas honom.
Och alla de brunnar som hans faders tjänare hade grävt i hans fader Abrahams tid, dem hade filistéerna kastat igen och fyllt med grus.
Och Abimelek sade till Isak: »Drag bort ifrån oss; ty du har blivit oss alltför mäktig.»
Då drog Isak bort därifrån och slog upp sitt läger i Gerars dal och bodde där.
Och Isak lät åter gräva ut de vattenbrunnar som hade blivit grävda i hans fader Abrahams tid, men som filistéerna efter Abrahams död hade kastat igen; och han gav dem åter de namn som hans fader hade givit dem.
Och Isaks tjänare grävde i dalen och funno där en brunn med rinnande vatten.
Men herdarna i Gerar begynte tvista med Isaks herdar och sade: »Vattnet är vårt.»
Då gav han den brunnen namnet Esek , eftersom de hade kivat med honom.
Därefter grävde de en annan brunn, men om den kommo de ock i tvist; då gav han den namnet Sitna .
Sedan begav han sig därifrån till en annan plats och grävde åter en brunn; om den tvistade de icke.
Därför gav han denna namnet Rehobot , i det han sade: »Nu har ju HERREN givit oss utrymme, så att vi kunna föröka oss i landet.»
Sedan drog han därifrån upp till Beer-Seba.
Och HERREN uppenbarade sig för honom den natten och sade: »Jag är Abrahams, din faders, Gud.
Frukta icke, ty jag är med dig, och jag skall välsigna dig och göra din säd talrik, för min tjänare Abrahams skull.»
Då byggde han där ett altare och åkallade HERRENS namn och slog där upp sitt tält.
Och Isaks tjänare grävde där en brunn.
Och Abimelek begav sig till honom från Gerar med Ahussat, sin vän, och Pikol, sin härhövitsman.
Men Isak sade till dem: »Varför kommen I till mig, I som haten mig och haven drivit mig ifrån eder?»
De svarade: »Vi hava tydligt sett att HERREN är med dig; därför tänkte vi: 'Låt oss giva varandra en ed, vi och du, så att vi sluta ett förbund med dig,
att du icke skall göra oss något ont, likasom vi å vår sida icke hava kommit vid dig, och likasom vi icke hava gjort dig annat än gott och hava låtit dig fara i frid.'
Du är nu HERRENS välsignade.»
Då gjorde han ett gästabud för dem, och de åto och drucko.
Bittida följande morgon svuro de varandra eden; sedan lät Isak dem gå, och de foro ifrån honom i frid.
Samma dag kommo Isaks tjänare och berättade för honom om den brunn som de hade grävt och sade till honom: »Vi hava funnit vatten.»
Och han kallade den Sibea.
Därav heter staden Beer-Seba ännu i dag.
När Esau var fyrtio år gammal, tog han till hustrur Judit, dotter till hetiten Beeri, och Basemat, dotter till hetiten Elon.
Men dessa blevo en hjärtesorg för Isak och Rebecka.
När Isak hade blivit gammal och hans ögon voro skumma, så att han icke kunde se, kallade han till sig Esau, sin äldste son, och sade till honom: »Min son!»
Han svarade honom: »Vad vill du?»
Då sade han: »Se, jag är gammal och vet icke när jag skall dö.
Så tag nu dina jaktredskap, ditt koger och din båge, och gå ut i marken och jaga villebråd åt mig;
red sedan till åt mig en smaklig rätt, en sådan som jag tycker om, och bär in den till mig till att äta, på det att min själ må välsigna dig, förrän jag dör.»
Men Rebecka hörde huru Isak talade till sin son Esau.
Och medan Esau gick ut i marken för att jaga villebråd till att föra hem,
sade Rebecka till sin son Jakob: »Se, jag har hört din fader tala så till din broder Esau:
'Hämta mig villebråd och red till åt mig en smaklig rätt, på det att jag må äta och sedan välsigna dig inför HERREN, förrän jag dör.'
Så hör nu vad jag säger, min son, och gör vad jag bjuder dig.
Gå bort till hjorden och hämta mig därifrån två goda killingar, så vill jag av dem tillreda en smaklig rätt åt din fader, en sådan som han tycker om.
Och du skall bära in den till din fader till att äta, på det att han må välsigna dig, förrän han dör.»
Men Jakob sade till sin moder Rebecka: »Min broder Esau är ju luden, och jag är slät.
Kanhända tager min fader på mig, och jag bliver då av honom hållen för en bespottare och skaffar mig förbannelse i stället för välsignelse.»
Då sade hans moder till honom: »Den förbannelsen komme över mig, min son; hör nu allenast vad jag säger, och gå och hämta dem åt mig.»
Då gick han och hämtade dem och bar dem till sin moder; och hans moder tillredde en smaklig rätt, en sådan som hans fader tyckte om.
Och Rebecka tog Esaus, sin äldre sons, högtidskläder, som hon hade hos sig i huset, och satte dem på Jakob, sin yngre son.
Och med skinnen av killingarna beklädde hon hans händer och den släta delen av hans hals.
Sedan lämnade hon åt sin son Jakob den smakliga rätten och brödet som hon hade tillrett.
Och han gick in till sin fader och sade: »Min fader!»
Han svarade: »Vad vill du?
Vem är du, min son?»
Då sade Jakob till sin fader: »Jag är Esau, din förstfödde.
Jag har gjort såsom du tillsade mig; sätt dig upp och ät av mitt villebråd, på det att din själ må välsigna mig.»
Men Isak sade till sin son: »Huru har du så snart kunnat finna något, min son?»
Han svarade: »HERREN, din Gud, skickade det i min väg.»
Då sade Isak till Jakob: »Kom hit, min son, och låt mig taga på dig och känna om du är min son Esau eller icke.»
Och Jakob gick fram till sin fader Isak; och när denne hade tagit på honom, sade han: »Rösten är Jakobs röst, men händerna äro Esaus händer.»
Och han kände icke igen honom, ty hans händer voro ludna såsom hans broder Esaus händer; och han välsignade honom.
Men han frågade: »Är du verkligen min son Esau?»
Han svarade: »Ja.»
Då sade han: »Bär hit maten åt mig och låt mig äta av min sons villebråd, på det att min själ må välsigna dig.»
Och han bar fram den till honom, och han åt; och han räckte honom vin, och han drack.
Därefter sade hans fader Isak till honom: »Kom hit och kyss mig, min son.»
När han då gick fram och kysste honom, kände han lukten av hans kläder och välsignade honom; han sade: »Se, av min son utgår doft, lik doften av en mark, som HERREN har välsignat.
Så give dig Gud av himmelens dagg och av jordens fetma och säd och vin i rikligt mått.
Folk tjäne dig, och folkslag falle ned för dig.
Bliv en herre över dina bröder, och må din moders söner falla ned för dig.
Förbannad vare den som förbannar dig, och välsignad vare den som välsignar dig!»
Men när Isak hade givit Jakob sin välsignelse och Jakob just hade gått ut från sin fader Isak, kom hans broder Esau hem från jakten.
Därefter tillredde också han en smaklig rätt och bar in den till sin fader och sade till sin fader: »Må min fader stå upp och äta av sin sons villebråd, på det att din själ må välsigna mig.»
Hans fader Isak frågade honom: »Vem är du?»
Han svarade: »Jag är Esau, din förstfödde son.»
Då blev Isak övermåttan häpen och sade: »Vem var då den jägaren som bar in till mig sitt villebråd, så att jag åt av allt, förrän du kom, och sedan välsignade honom?
Välsignad skall han ock förbliva.»
När Esau hörde sin faders ord, brast han ut i högljudd och bitter klagan och sade till sin fader: »Välsigna också mig, min fader.»
Men han svarade: »Din broder har kommit med svek och tagit din välsignelse.»
Då sade han: »Han heter ju Jakob, och han har nu också två gånger bedragit mig.
Min förstfödslorätt har han tagit, och se, nu har han ock tagit min välsignelse.»
Och han frågade: »Har du då ingen välsignelse kvar för mig?»
Isak svarade och sade till Esau: »Se, jag har satt honom till en herre över dig, och alla hans bröder har jag givit honom till tjänare, och med säd och vin har jag begåvat honom; vad skall jag då nu göra för dig, min son?»
Esau sade till sin fader: »Har du då allenast den enda välsignelsen, min fader?
Välsigna också mig, min fader.»
Och Esau brast ut i gråt.
Då svarade hans fader Isak och sade till honom: »Se, fjärran ifrån jordens fetma skall din boning vara och utan dagg från himmelen ovanefter.
Av ditt svärd skall du leva, och du skall tjäna din broder.
Men det skall ske, när du samlar din kraft, att du river hans ok från din hals.»
Och Esau blev hätsk mot Jakob för den välsignelses skull som hans fader hade givit honom.
Och Esau sade vid sig själv: »Snart skola de dagar komma, då vi få sörja vår fader; då skall jag dräpa min broder Jakob.»
När man nu berättade för Rebecka vad hennes äldre son Esau hade sagt, sände hon och lät kalla till sig sin yngre son Jakob och sade till honom: »Se, din broder Esau vill hämnas på dig och dräpa dig.
Så hör nu vad jag säger, min son: stå upp och fly till min broder Laban i Haran,
och stanna någon tid hos honom, till dess din broders förbittring har upphört,
ja, till dess din broders vrede mot dig har upphört och han förgäter vad du har gjort mot honom.
Då skall jag sända åstad och hämta dig därifrån.
Varför skall jag mista eder båda på samma gång?»
Och Rebecka sade till Isak: »Jag är led vid livet för Hets döttrars skull.
Om Jakob tager hustru bland Hets döttrar, en sådan som dessa, någon bland landets döttrar, varför skulle jag då leva?»
Då kallade Isak till sig Jakob och välsignade honom; och han bjöd honom och sade till honom: »Tag dig icke till hustru någon av Kanaans döttrar,
utan stå upp och begiv dig till Paddan-Aram, till Betuels, din morfaders, hus, och tag dig en hustru därifrån, någon av Labans, din morbroders, döttrar.
Och må Gud den Allsmäktige välsigna dig och göra dig fruktsam och föröka dig, så att skaror av folk komma av dig;
må han giva åt dig Abrahams välsignelse, åt dig och din säd med dig, så att du får taga i besittning det land som Gud har givit åt Abraham, och där du nu bor såsom främling.»
Så sände Isak åstad Jakob, och denne begav sig till Paddan-Aram, till araméen Laban, Betuels son, som var broder till Rebecka, Jakobs och Esaus moder.
När nu Esau såg att Isak hade välsignat Jakob och sänt honom till Paddan-Aram för att därifrån taga sig hustru -- ty han hade välsignat honom och bjudit honom och sagt: »Du skall icke taga till hustru någon av Kanaans döttrar» --
och när han såg att Jakob hade lytt sin fader och moder och begivit sig till Paddan-Aram,
då märkte Esau att Kanaans döttrar misshagade hans fader Isak;
och Esau gick bort till Ismael och tog Mahalat, Abrahams son Ismaels dotter, Nebajots syster, till hustru åt sig, utöver de hustrur han förut hade.
Men Jakob begav sig från Beer-Seba på väg till Haran.
Och han kom då till den heliga platsen och stannade där över natten, ty solen hade gått ned; och han tog en av stenarna på platsen för att hava den till huvudgärd och lade sig att sova där.
Då hade han en dröm.
Han såg en stege vara rest på jorden, och dess övre ände räckte upp till himmelen, och Guds änglar stego upp och ned på den.
Och se, HERREN stod framför honom och sade: »Jag är HERREN, Abrahams, din faders, Gud och Isaks Gud.
Det land där du ligger skall jag giva åt dig och din säd.
Och din säd skall bliva såsom stoftet på jorden, och du skall utbreda dig åt väster och öster och norr och söder, och alla släkter på jorden skola varda välsignade i dig och i din säd.
Och se, jag är med dig och skall bevara dig, varthelst du går, och jag skall föra dig tillbaka till detta land; ty jag skall icke övergiva dig, till dess jag har gjort vad jag har lovat dig.»
När Jakob vaknade upp ur sömnen sade han: »HERREN är sannerligen på denna plats, och jag visste det icke!»
Och han betogs av fruktan och sade: »Detta måste vara en helig plats, här bor förvisso Gud, och här är himmelens port.»
Och bittida om morgonen stod Jakob upp och tog stenen som han hade haft till huvudgärd och reste den till en stod och göt olja därovanpå.
Och han gav den platsen namnet Betel; förut hade staden hetat Lus.
Och Jakob gjorde ett löfte och sade: »Om Gud är med mig och bevarar mig under den resa som jag nu är stadd på och giver mig bröd till att äta och kläder till att kläda mig med,
så att jag kommer i frid tillbaka till min faders hus, då skall HERREN vara min Gud;
och denna sten som jag har rest till en stod skall bliva ett Guds hus, och av allt vad du giver mig skall jag giva dig tionde.»
Och Jakob begav sig åstad på väg till Österlandet.
Där fick han se en brunn på fältet, och vid den lågo tre fårhjordar, ty ur denna brunn plägade man vattna hjordarna.
Och stenen som låg över brunnens öppning var stor;
därför plägade man låta alla hjordarna samlas dit och vältrade så stenen från brunnens öppning och vattnade fåren; sedan lade man stenen tillbaka på sin plats över brunnens öppning.
Och Jakob sade till männen: »Mina bröder, varifrån ären I?»
De svarade: »Vi äro från Haran.»
Då sade han till dem: »Kännen I Laban, Nahors son?»
De svarade: »Ja.»
Han frågade dem vidare: »Står det väl till med honom?»
De svarade: »Ja; och se, där kommer hans dotter Rakel med fåren.»
Han sade: »Det är ju ännu full dag; ännu är det icke tid att samla boskapen.
Vattnen fåren, och fören dem åter i bet.»
Men de svarade: »Vi kunna icke göra det, förrän alla hjordarna hava blivit samlade och man har vältrat stenen från brunnens öppning; då vattna vi fåren.»
Medan han ännu talade med dem, hade Rakel kommit dit med sin faders får; ty hon plägade vakta dem.
När Jakob fick se sin morbroder Labans dotter Rakel komma med Labans, hans morbroders, får, gick han fram och vältrade stenen från brunnens öppning och vattnade sin morbroder Labans får.
Och Jakob kysste Rakel och brast ut i gråt.
Och Jakob omtalade för Rakel att han var hennes faders frände, och att han var Rebeckas son; och hon skyndade åstad och omtalade det för sin fader.
Då nu Laban fick höras talas om sin systerson Jakob, skyndade han emot honom och tog honom i famn och kysste honom och förde honom in i sitt hus; och han förtäljde för Laban allt som hade hänt honom.
Och Laban sade till honom: »Ja, du är mitt kött och ben.»
Och han stannade hos honom en månads tid.
Och Laban sade till Jakob: »Du är ju min frände.
Skulle du då tjäna mig för intet?
Säg mig vad du vill hava i lön?»
Nu hade Laban två döttrar; den äldre hette Lea, och den yngre hette Rakel.
Och Leas ögon voro matta, men Rakel hade en skön gestalt och var skön att skåda.
Och Jakob hade fattat kärlek till Rakel; därför sade han: »Jag vill tjäna dig i sju år för Rakel, din yngre dotter.»
Laban svarade: »Det är bättre att jag giver henne åt dig, än att jag skulle giva henne åt någon annan; bliv kvar hos mig.»
Så tjänade Jakob för Rakel i sju år, och det tycktes honom vara allenast några dagar; så kär hade han henne.
Därefter sade Jakob till Laban: »Giv mig min hustru, ty min tid är nu förlupen; låt mig gå in till henne.»
Då bjöd Laban tillhopa allt folket på orten och gjorde ett gästabud.
Men när aftonen kom, tog han sin dotter Lea och förde henne till honom, och han gick in till henne.
Och Laban gav sin tjänstekvinna Silpa åt sin dotter Lea till tjänstekvinna.
Om morgonen fick Jakob se att det var Lea.
Då sade han till Laban: »Vad har du gjort mot mig?
Var det icke för Rakel jag tjänade hos dig?
Varför har du så bedragit mig?»
Laban svarade: »Det är icke sed på vår ort att man giver bort den yngre före den äldre.
Låt nu dennas bröllopsvecka gå till ända, så vilja vi giva dig också den andra, mot det att du gör tjänst hos mig i ännu ytterligare sju år.»
Och Jakob samtyckte härtill och lät hennes bröllopsvecka gå till ända.
Sedan gav han honom sin dotter Rakel till hustru.
Och Laban gav sin tjänstekvinna Bilha åt sin dotter Rakel till tjänstekvinna.
Så gick han in också till Rakel, och han hade Rakel kärare än Lea.
Sedan tjänade han hos honom i ännu ytterligare sju år.
Men då HERREN såg att Lea var försmådd, gjorde han henne fruktsam, medan Rakel var ofruktsam.
Och Lea blev havande och födde en son, och hon gav honom namnet Ruben, ty hon tänkte: »HERREN har sett till mitt lidande ; ja, nu skall min man hava mig kär.»
Och hon blev åter havande och födde en son.
Då sade hon: »HERREN har hört att jag har varit försmådd, därför har han givit mig också denne.»
Och hon gav honom namnet Simeon.
Och åter blev hon havande och födde en son.
Då sade hon: »Nu skall väl ändå min man hålla sig till mig; jag har ju fött honom tre söner.»
Därav fick denne namnet Levi.
Åter blev hon havande och födde en son.
Då sade hon: »Nu vill jag tacka HERREN.»
Därför gav hon honom namnet Juda.
Sedan upphörde hon att föda.
Då nu Rakel såg att hon icke födde barn åt Jakob, avundades hon sin syster och sade till Jakob: »Skaffa mig barn, eljest dör jag.»
Då upptändes Jakobs vrede mot Rakel, och han svarade: »Håller du då mig för Gud?
Det är ju han som förmenar dig livsfrukt.»
Hon sade: »Se, där är min tjänarinna Bilha; gå in till henne, för att hon må föda barn i mitt sköte, så att genom henne också jag får avkomma.»
Så gav hon honom sin tjänstekvinna Bilha till hustru, och Jakob gick in till henne.
Och Bilha blev havande och födde åt Jakob en son.
Då sade Rakel: »Gud har skaffat rätt åt mig; han har hört min röst och givit mig en son.»
Därför gav hon honom namnet Dan.
Åter blev Bilha, Rakels tjänstekvinna, havande, och hon födde åt Jakob en andre son.
Då sade Rakel: »Strider om Gud har jag stritt med min syster och har vunnit seger.»
Och hon gav honom namnet Naftali.
Då Lea nu såg att hon hade upphört att föda, tog hon sin tjänstekvinna Silpa och gav henne åt Jakob till hustru.
Och Silpa, Leas tjänstekvinna, födde åt Jakob en son.
Då sade Lea: »Till lycka !»
Och hon gav honom namnet Gad.
Och Silpa, Leas tjänstekvinna, födde åt Jakob en andre son.
Då sade Lea: »Till sällhet för mig!
Ja, jungfrur skola prisa mig säll.»
Och hon gav honom namnet Aser.
Men Ruben gick ut en gång vid tiden för veteskörden och fann då kärleksäpplen på marken och bar dem till sin moder Lea.
Då sade Rakel till Lea: »Giv mig några av din sons kärleksäpplen.»
Men hon svarade henne: »Är det icke nog att du har tagit min man?
Vill du ock taga min sons kärleksäpplen?»
Rakel sade: »Må han då i natt ligga hos dig, om jag får din sons kärleksäpplen.»
När nu Jakob om aftonen kom hem från marken, gick Lea honom till mötes och sade: »Till mig skall du gå in; ty jag har givit min sons kärleksäpplen såsom lön för dig.»
Så låg han hos henne den natten.
Och Gud hörde Lea, så att hon blev havande, och hon födde åt Jakob en femte son.
Då sade Lea: »Gud har givit mig min lön , för det att jag gav min tjänstekvinna åt min man.»
Och hon gav honom namnet Isaskar.
Åter blev Lea havande, och hon födde åt Jakob en sjätte son.
Då sade Lea: »Gud har givit mig en god gåva .
Nu skall min man förbliva boende hos mig, ty jag har fött honom sex söner.»
Och hon gav honom namnet Sebulon.
Därefter födde hon en dotter och gav henne namnet Dina.
Men Gud tänkte på Rakel; Gud hörde henne och gjorde henne fruktsam.
Hon blev havande och födde en son.
Då sade hon: »Gud har tagit bort min smälek.»
Och hon gav honom namnet Josef, i det hon sade: »HERREN give mig ännu en son.»
Då nu Rakel hade fött Josef, sade Jakob till Laban: »Låt mig fara; jag vill draga hem till min ort och till mitt land.
Giv mig mina hustrur och mina barn, som jag har tjänat dig för, och låt mig draga hem; du vet ju själv huru jag har tjänat dig.»
Laban svarade honom: »Låt mig finna nåd för dina ögon; jag vet genom hemliga tecken att HERREN för din skull har välsignat mig.»
Och han sade ytterligare: »Bestäm vad du vill hava i lön av mig, så skall jag giva dig det.»
Han svarade honom: »Du vet själv huru jag har tjänat dig, och vad det har blivit av din boskap under min vård.
Ty helt litet var det som du hade, förrän jag kom, men det har förökat sig och blivit mycket, ty HERREN har välsignat dig, varhelst jag har gått fram.
Men när skall jag nu också få göra något för mitt eget hus?»
Han svarade: »Vad skall jag giva dig?»
Och Jakob sade: »Du skall icke alls giva mig något.
Om du vill göra mot mig såsom jag nu säger, så skall jag fortfara att vara herde för din hjord och vakta den.
Jag vill i dag gå igenom hela din hjord och avskilja ur den alla spräckliga och brokiga såväl som alla svarta djur bland fåren, så ock vad som är brokigt och spräckligt bland getterna; sådant må sedan bliva min lön.
Och när du framdeles kommer för att med egna ögon se vad som har blivit min lön, då skall min rättfärdighet vara mitt vittne; alla getter hos mig, som icke äro spräckliga eller brokiga, och alla får hos mig, som icke äro svarta, de skola räknas såsom stulna.»
Då sade Laban: »Välan, blive det såsom du har sagt.»
Och samma dag avskilde han de strimmiga och brokiga bockarna och alla spräckliga och brokiga getter -- alla djur som något vitt fanns på -- och alla svarta djur bland fåren; och detta lämnade han i sina söners vård.
Och han lät ett avstånd av tre dagsresor vara mellan sig och Jakob.
Och Jakob fick Labans övriga hjord att vakta.
Men Jakob tog sig friska käppar av poppel, mandelträd och lönn och skalade på dem vita ränder, i det han blottade det vita på käpparna.
Sedan lade han käpparna, som han hade skalat, i rännorna eller vattenhoarna dit hjordarna kommo för att dricka, så att djuren hade dem framför sig; och de hade just sin parningstid, när de nu kommo för att dricka.
Och djuren parade sig vid käpparna, och så blev djurens avföda strimmig, spräcklig och brokig.
Därefter avskilde Jakob lammen och ordnade djuren så, att de vände huvudena mot det som var strimmigt och mot allt som var svart i Labans hjord; så skaffade han sig egna hjordar, som han icke lät komma ihop med Labans hjord.
Och så ofta de kraftigare djuren skulle para sig, lade Jakob käpparna framför djurens ögon i rännorna, så att de parade sig vid käpparna.
Men när det var de svagare djuren, lade han icke dit dem.
Härigenom tillföllo de svaga Laban och de kraftiga Jakob.
Så blev mannen övermåttan rik; han fick mycken småboskap, därtill ock tjänarinnor och tjänare, kameler och åsnor.
Men han fick höra huru Labans söner talade så: »Jakob har tagit allt vad vår fader ägde; av det vår fader ägde är det som han har skaffat sig all denna rikedom.»
Jakob märkte också att Laban icke såg på honom med samma ögon som förut.
Och HERREN sade till Jakob: »Vänd tillbaka till dina fäders land och till din släkt; jag skall vara med dig.»
Då sände Jakob och lät kalla Rakel och Lea ut på marken till sin hjord;
och han sade till dem: »Jag märker att eder fader icke ser på mig med samma ögon som förut, nu då min faders Gud har varit med mig.
Och I veten själva att jag har tjänat eder fader av alla mina krafter;
men eder fader har handlat svikligt mot mig och tio gånger förändrat min lön.
Dock har Gud icke tillstatt honom att göra mig något ont.
När han sade: 'De spräckliga skola vara din lön', då fick hela hjorden spräcklig avföda; och när han sade: 'De strimmiga skola vara din lön', då fick hela jorden strimmig avföda.
Så tog Gud eder faders boskap och gav den åt mig.
Ty när parningstiden kom, lyfte jag upp mina ögon och fick se i drömmen att hannarna som betäckte småboskapen voro strimmiga, spräckliga och fläckiga.
Och Guds ängel sade till mig i drömmen: 'Jakob!'
Jag svarade: 'Här är jag.'
Då sade han: 'Lyft upp dina ögon och se huru alla hannar som betäcka småboskapen äro strimmiga, spräckliga och fläckiga.
Jag har ju sett allt vad Laban gör mot dig.
Jag är den Gud som du såg i Betel, där du smorde en stod, och där du gjorde mig ett löfte.
Stå nu upp och drag ut ur detta land, och vänd tillbaka till ditt fädernesland.'»
Då svarade Rakel och Lea och sade till honom: »Hava vi numera någon lott eller arvedel i vår faders hus?
Blevo vi icke av honom aktade såsom främlingar, när han sålde oss?
Sedan har han ju ock förtärt vad han fick i betalning för oss.
Ja, all den rikedom som Gud har avhänt vår fader tillhör oss och våra barn.
Så gör nu allt vad Gud har sagt dig.»
Då stod Jakob upp och satte sina barn och sina hustrur på kamelerna
och förde bort med sig all boskap och alla ägodelar som han hade förvärvat, den boskap han ägde, och som han hade förvärvat i Paddan-Aram, och begav sig på väg till sin fader Isak i Kanaans land.
Men Laban hade gått bort för att klippa sina får; då stal Rakel sin faders husgudar,
och Jakob stal sig undan från araméen Laban, så att han icke lät denne märka att han ämnade fly.
Så flydde han med allt sitt; han bröt upp och gick över floden och ställde sin färd mot Gileads berg.
Men på tredje dagen fick Laban veta att Jakob hade flytt.
Då tog han med sig sina fränder och satte efter honom sju dagsresor och hann upp honom på Gileads berg.
Men Gud kom till araméen Laban i en dröm om natten och sade till honom: »Tag dig till vara för att tala något mot Jakob, vad det vara må.»
Och Laban hann upp Jakob.
Denne hade då slagit upp sitt tält på berget, och Laban med sina fränder hade ock sitt tält uppslaget på Gileads berg.
Då sade Laban till Jakob: »Vad är detta för ett tilltag, att du har stulit dig undan från mig och fört bort mina döttrar, likasom vore de tagna med svärd?
Varför dolde du din flykt och stal dig undan från mig?
Därigenom att du icke lät mig veta något därom hindrades jag att ledsaga dig till vägs med jubel och sång, med pukor och harpor.
Du förunnade mig icke ens att kyssa mina barnbarn och mina döttrar.
Du har handlat dåraktigt.
Det stode nu i min makt att göra eder ont; men eder faders Gud sade till mig i natt: 'Tag dig till vara för att tala något mot Jakob, vad det vara må.'
Och då du nu äntligen ville fara, eftersom du längtade så mycket till din faders hus, varför skulle du stjäla mina gudar?»
Då svarade Jakob och sade till Laban: »Jag fruktade för dig, ty jag tänkte att du skulle med våld taga dina döttrar ifrån mig.
Men den som du finner dina gudar hos, han skall icke få behålla livet.
I våra fränders närvaro må du se efter, om något är ditt av det jag har i min ägo, och i så fall taga det.»
Ty Jakob visste icke att Rakel hade stulit dem.
Då gick Laban in i Jakobs tält, därefter i Leas tält och i de båda tjänstekvinnornas tält, men fann intet.
Och när han hade kommit ut ur Leas tält, gick han in i Rakels tält.
Men Rakel hade tagit husgudarna och lagt dem i kamelsadeln och satt sig därovanpå.
Och Laban sökte igenom hela tältet, men fann dem icke.
Och hon sade till sin fader: »Vredgas icke, min herre, över att jag ej kan stiga upp för dig, ty det är med mig på kvinnors vis.»
Så sökte han efter husgudarna, men fann dem icke.
Då blev Jakob vred och for ut mot Laban; Jakob tog till orda och sade till Laban: »Vari har jag då förbrutit mig eller syndat, eftersom du så häftigt förföljer mig?
Nu har du genomsökt allt mitt bohag; vad har du där funnit av bohagsting som tillhöra dig?
Lägg det fram här inför mina fränder och dina fränder, så att de få döma mellan oss båda.
I tjugu år har jag nu varit hos dig; dina tackor och dina getter hava icke fött i otid, och av vädurarna i din hjord har jag icke ätit.
Intet ihjälrivet djur förde jag till dig; jag måste själv ersätta det; du utkrävde det av mig, evad det var stulet om dagen eller stulet om natten.
Sådan var min lott: om dagen förtärdes jag av hetta och om natten av köld, och sömnen flydde mina ögon.
I tjugu år har jag nu varit i ditt hus; jag har tjänat dig i fjorton år för dina båda döttrar och i sex år för din boskap, men du har tio gånger förändrat min lön.
Om icke min faders Gud hade varit med mig, Abrahams Gud, han som ock Isak fruktar, så hade du nu säkert låtit mig fara med tomma händer.
Men Gud såg mitt lidande och min möda, och han fällde domen i natt.»
Då svarade Laban och sade till Jakob: »Döttrarna äro mina döttrar, och barnen äro mina barn, och hjordarna äro mina hjordar, och allt det du ser är mitt; vad skulle jag då nu kunna göra mot dessa mina döttrar eller mot barnen som de hava fött?
Så kom nu och låt oss sluta ett förbund med varandra, och må det vara ett vittne mellan mig och dig.»
Då tog Jakob en sten och reste den till en stod.
Och Jakob sade till sina fränder: »Samlen tillhopa stenar.»
Och de togo stenar och gjorde ett röse och höllo måltid där på röset.
Och Laban kallade det Jegar-Sahaduta , men Jakob kallade det Galed .
Och Laban sade: »Detta röse vare i dag vittne mellan mig och dig.»
Därav fick det namnet Galed;
men det kallades ock Mispa , ty han sade: »HERREN vare väktare mellan mig och dig, när vi icke mer se varandra.
Om du behandlar mina döttrar illa eller tager andra hustrur jämte mina döttrar, så vet, att om ock ingen människa är tillstädes, så är dock Gud vittne mellan mig och dig.»
Och Laban sade ytterligare till Jakob: »Se, detta röse och stoden som jag har rest mellan mig och dig --
detta röse vare ett vittne, och stoden vare ett vittne, att jag icke skall draga till dig förbi detta röse, och att icke heller du skall draga till mig förbi detta röse och denna stod, med ont uppsåt.
Abrahams Gud och Nahors Gud, han som var deras faders Gud, han vare domare mellan oss.»
Och Jakob svor eden vid honom som hans fader Isak fruktade.
Och Jakob offrade ett slaktoffer på berget och inbjöd sina fränder att hålla måltid med sig.
Och de åto och stannade sedan på berget över natten.
Men om morgonen stod Laban bittida upp, och sedan han hade kysst sina barnbarn och sina döttrar och välsignat dem, for han sin väg hem igen.
Men när Jakob drog sin väg fram, mötte honom Guds änglar;
och då Jakob såg dem, sade han: »Detta är Guds skara.»
Och han gav den platsen namnet Mahanaim .
Och Jakob sände budbärare framför sig till sin broder Esau i Seirs land, på Edoms mark;
och han bjöd dem och sade: »Så skolen I säga till min herre Esau: Din tjänare Jakob låter säga: Jag har vistats borta hos Laban och dröjt kvar där ända till nu;
och jag har fått oxar, åsnor, får, tjänare och tjänarinnor.
Och jag har nu velat sända bud för att låta min herre veta detta, på det att jag må finna nåd för dina ögon.»
När sedan budbärarna kommo tillbaka till Jakob, sade de: »Vi träffade din broder Esau, som redan drager emot dig med fyra hundra man.»
Då blev Jakob mycket förskräckt och betogs av ångest; och han delade sitt folk och fåren och fäkreaturen och kamelerna i två skaror.
Ty han tänkte: »Om Esau överfaller den ena skaran och slår den, så kan dock den andra skaran undkomma.»
Och Jakob sade: »Min fader Abrahams Gud och min fader Isaks Gud, HERRE, du som sade till mig: 'Vänd tillbaka till ditt land och till din släkt, så skall jag göra dig gott',
jag är för ringa till all den nåd och all den trofasthet som du har bevisat din tjänare; ty jag hade icke mer än min stav, när jag gick över denna Jordan, och nu har jag förökats till två skaror.
Rädda mig undan min broder Esaus hand, ty jag fruktar att han kommer och förgör mig, utan att ens skona mödrar och barn.
Du har själv sagt: 'Jag skall göra dig mycket gott och låta din säd bliva såsom havets sand, som man icke kan räkna för dess myckenhets skull.'»
Och han stannade där den natten.
Och av det han hade förvärvat tog han ut till skänker åt sin broder Esau
två hundra getter och tjugu bockar, två hundra tackor och tjugu vädurar,
trettio kamelston som gåvo di, jämte deras föl, därtill fyrtio kor och tio tjurar samt tjugu åsninnor med tio föl.
Och han lämnade detta i sina tjänares vård, var hjord för sig, och sade till sina tjänare: »Gån framför mig och låten ett mellanrum vara mellan hjordarna.»
Och han bjöd den förste och sade: »När min broder Esau möter dig och frågar dig: 'Vem tillhör du, och vart går du, och vem tillhöra djuren som du driver framför dig?',
då skall du svara: 'De tillhöra din tjänare Jakob; de äro skänker som han sänder till min herre Esau, och själv kommer han här efter oss.'»
Och han bjöd likaledes den andre och den tredje och alla de övriga som drevo hjordarna: »Såsom jag nu har sagt eder skolen I säga till Esau, när I kommen fram till honom.
Och I skolen vidare säga: 'Också din tjänare Jakob kommer här efter oss.'»
Ty han tänkte: »Jag vill blidka honom med de skänker som gå före mig; sedan vill jag själv komma inför hans ansikte; kanhända tager han då nådigt emot mig.»
Så kommo nu skänkerna före honom, medan han själv den natten stannade i lägret.
Men under natten stod han upp och tog sina båda hustrur och sina båda tjänstekvinnor och sina elva söner och gick över Jabboks vad.
Han tog dem och förde dem över bäcken och förde tillika över vad han eljest ägde.
Och Jakob blev ensam kvar.
Då brottades en man med honom, till dess morgonrodnaden gick upp.
Och när denne såg att han icke kunde övervinna Jakob, gav han honom ett slag på höftleden, så att höften gick ur led, under det han brottades med honom.
Och mannen sade: »Släpp mig, ty morgonrodnaden går upp.»
Men han svarade: »Jag släpper dig icke, med mindre du välsignar mig.»
Då sade han till honom: »Vad är ditt namn?»
Han svarade: »Jakob.»
Han sade: »Du skall icke mer heta Jakob, utan Israel, ty du har kämpat med Gud och med människor och vunnit seger.»
Då frågade Jakob och sade: »Låt mig veta ditt namn.»
Han svarade: »Varför frågar du efter mitt namn?»
Och han välsignade honom där.
Men Jakob gav platsen namnet Peniel , »ty», sade han, »jag har sett Gud ansikte mot ansikte, och dock har mitt liv blivit räddat».
Och när han hade kommit förbi Penuel, såg han solen gå upp; men han haltade på höften.
Fördenskull äta Israels barn ännu i dag icke höftsenan som ligger på höftleden, därför nämligen, att han gav Jakob ett slag på höftleden, på höftsenan.
Och Jakob lyfte upp sina ögon och fick se Esau komma med fyra hundra man.
Då fördelade han sina barn på Lea och Rakel och de båda tjänstekvinnorna.
Och han lät tjänstekvinnorna med deras barn gå främst, Lea med hennes barn därnäst, och Rakel med Josef sist.
Och själv gick han framför dem och bugade sig sju gånger ned till jorden, till dess han kom fram till sin broder.
Men Esau skyndade emot honom och tog honom i famn och föll honom om halsen och kysste honom; och de gräto.
Och när han lyfte upp sina ögon och fick se kvinnorna och barnen, sade han: »Vilka äro dessa som du har med dig?»
Han svarade: »Det är barnen som Gud har beskärt din tjänare.»
Och tjänstekvinnorna gingo fram med sina barn och bugade sig.
Därefter gick ock Lea fram med sina barn, och de bugade sig.
Slutligen gingo Josef och Rakel fram och bugade sig.
Sedan frågade han: »Vad ville du med hela den skara som jag mötte?»
Han svarade: »Jag ville finna nåd för min herres ögon.»
Men Esau sade: »Jag har nog; behåll du vad du har, min broder.»
Jakob svarade: »Ack nej; om jag har funnit nåd för dina ögon, så tag emot skänkerna av mig, eftersom jag har fått se ditt ansikte, likasom såge jag ett gudaväsens ansikte, då du nu så gunstigt har tagit emot mig.
Tag hälsningsskänkerna som jag har skickat emot dig; ty Gud har varit mig nådig, och jag har allt fullt upp.»
Och han bad honom så enträget, att han tog emot dem.
Och Esau sade: »Låt oss bryta upp och draga vidare; jag vill gå framför dig.»
Men han svarade honom: »Min herre ser själv att barnen äro späda, och att jag har med mig får och kor som giva di; driver man dessa för starkt en enda dag, så dör hela hjorden.
Må därför min herre draga åstad före sin tjänare, så vill jag komma efter i sakta mak, i den mån boskapen, som drives framför mig, och barnen orka följa med, till dess jag kommer till min herre i Seir.»
Då sade Esau: »Så vill jag åtminstone lämna kvar hos dig en del av mitt folk.»
Men han svarade: »Varför så?
Må jag allenast finna nåd för min herres ögon.»
Så vände Esau om, samma dag, och tog vägen till Seir.
Men Jakob bröt upp och drog till Suckot och byggde sig där ett hus.
Och åt sin boskap gjorde han lövhyddor ; därav fick platsen namnet Suckot.
Och Jakob kom på sin färd ifrån Paddan-Aram välbehållen till Sikems stad i Kanaans land och slog upp sitt läger utanför staden.
Och det jordstycke där han hade slagit upp sitt tält köpte han av Hamors, Sikems faders, barn för hundra kesitor.
Och han reste där ett altare och kallade det El-Elohe-Israel .
Men Dina, den dotter som Lea hade fött åt Jakob, gick ut för att besöka landets döttrar.
Och Sikem, som var son till hivéen Hamor, hövdingen i landet, fick se henne, och han tog henne till sig och lägrade henne och kränkte henne.
Och hans hjärta fäste sig vid Dina, Jakobs dotter, och flickan blev honom kär, och han talade vänligt med flickan.
Och Sikem sade till sin fader Hamor: »Skaffa mig denna flicka till hustru.»
Och Jakob hade fått höra att hans dotter Dina hade blivit skändad.
Men eftersom hans söner voro med hans boskap ute på marken, teg Jakob, till dess de kommo hem.
Så gick nu Hamor, Sikems fader, ut till Jakob för att tala med honom.
Men när Jakobs söner kommo hem från marken, sedan de hade fått höra vad som hade hänt, blevo de förbittrade och vredgades högeligen över att han hade gjort vad som var en galenskap i Israel, i det han hade lägrat Jakobs dotter -- en otillbörlig gärning.
Då talade Hamor med dem och sade: »Min son Sikems hjärta har fäst sig vid eder syster; given henne åt honom till hustru.
Och befrynden eder med oss; given edra döttrar åt oss, och tagen I våra döttrar till hustrur,
och bosätten eder hos oss, ty landet skall ligga öppet för eder; där mån I bo och draga omkring och förvärva besittningar.»
Och Sikem sade till hennes fader och hennes bröder: »Låten mig finna nåd för edra ögon; vad I fordren av mig vill jag giva.
Begären av mig huru stor brudgåva och skänk som helst; jag vill giva vad I fordren av mig; given mig allenast flickan till hustru.»
Då svarade Jakobs söner Sikem och hans fader Hamor med listiga ord, eftersom han hade skändat deras syster Dina,
och sade till dem: »Vi kunna icke samtycka till att giva vår syster åt en man som har förhud; ty sådant hålla vi för skamligt.
Allenast på det villkoret skola vi göra eder till viljes, att I bliven såsom vi, därigenom att allt mankön bland eder omskäres.
Då skola vi giva våra döttrar åt eder och själva taga edra döttrar till hustrur; och vi skola då bo hos eder och bliva med eder ett enda folk.
Men om I icke viljen lyssna till oss och låta omskära eder, så skola vi taga vår syster och draga bort.»
Och Hamor och Sikem, Hamors son, voro till freds med vad de begärde.
Och den unge mannen dröjde icke att göra så, ty han hade fått behag till Jakobs dotter.
Och han hade större myndighet än någon annan i hans faders hus.
Så trädde då Hamor och hans son Sikem upp i sin stads port och talade till männen i staden och sade:
»Dessa män äro fredligt sinnade mot oss; må vi alltså låta dem bo i landet och draga omkring där; landet har ju utrymme nog för dem.
Vi vilja taga deras döttrar till hustrur åt oss och giva dem våra döttrar.
Men allenast på det villkoret skola männen göra oss till viljes och bo hos oss och bliva ett enda folk med oss, att allt mankön bland oss omskäres, likasom de själva äro omskurna.
Och då bliva ju deras boskap och deras egendom och alla deras dragare vår tillhörighet.
Må vi fördenskull allenast göra dem till viljes, så skola de bo kvar hos oss.»
Och folket lydde Hamor och hans son Sikem, alla de som bodde inom hans stadsport; allt mankön, så många som bodde inom hans stadsport, läto omskära sig.
Men på tredje dagen, då de voro sjuka av såren, togo Jakobs två söner Simeon och Levi, Dinas bröder, var sitt svärd och överföllo staden oförtänkt och dräpte allt mankön.
Också Hamor och hans son Sikem dräpte de med svärdsegg och togo Dina ut ur Sikems hus och gingo sin väg.
Och Jakobs söner kommo över de slagna och plundrade staden, därför att deras syster hade blivit skändad;
de togo deras får och fäkreatur och åsnor, både vad som fanns i staden och vad som fanns på fältet.
Och allt deras gods och alla deras barn och deras kvinnor förde de bort såsom byte, tillika med allt annat som fanns i husen.
Men Jakob sade till Simeon och Levi: »I haven dragit olycka över mig, då I nu haven gjort mig förhatlig för landets inbyggare, kananéerna och perisséerna.
Mitt folk är allenast en ringa hop; man skall nu församla sig mot mig och slå mig ihjäl; så skall jag med mitt hus förgöras.»
Men de svarade: »Skulle man då få behandla vår syster såsom en sköka?»
Och Gud sade till Jakob: »Stå upp, drag till Betel och stanna där, och res där ett altare åt den Gud som uppenbarade sig för dig, när du flydde för din broder Esau.»
Då sade Jakob till sitt husfolk och till alla som voro med honom: »Skaffen bort de främmande gudar som I haven bland eder, och renen eder och byten om kläder,
och låt oss så stå upp och draga till Betel; där vill jag resa ett altare åt den Gud som bönhörde mig, när jag var i nöd, och som var med mig på den väg jag vandrade.»
Då gåvo de åt Jakob alla de främmande gudar som de hade hos sig, därtill ock sina örringar; och Jakob grävde ned detta under terebinten vid Sikem.
Sedan bröto de upp; och en förskräckelse ifrån Gud kom över de kringliggande städerna, så att man icke förföljde Jakobs söner.
Och Jakob kom till Lus, det är Betel, i Kanaans land, jämte allt det folk som var med honom.
Och han byggde där ett altare och kallade platsen El-Betel , därför att Gud där hade uppenbarat sig för honom, när han flydde för sin broder.
Och Debora, Rebeckas amma, dog och blev begraven nedanför Betel, under en ek; den fick namnet Gråtoeken.
Och Gud uppenbarade sig åter för Jakob, när han hade kommit tillbaka från Paddan-Aram, och välsignade honom.
Och Gud sade till honom: »Ditt namn är Jakob; men du skall icke mer heta Jakob, utan Israel skall vara ditt namn.»
Så fick han namnet Israel.
Och Gud sade till honom: »Jag är Gud den Allsmäktige; var fruktsam och föröka dig.
Ett folk, ja, skaror av folk skola komma av dig, och konungar skola utgå från din länd.
Och det land som jag har givit åt Abraham och Isak skall jag giva åt dig; åt din säd efter dig skall jag ock giva det landet.
Och Gud for upp från honom, på den plats där han hade talat med honom.
Men Jakob reste en stod på den plats där han hade talat med honom, en stod av sten; och han offrade drickoffer därpå och göt olja över den.
Och Jakob gav åt platsen där Gud hade talat med honom namnet Betel.
Sedan bröto de upp från Betel.
Och när det ännu var ett stycke väg fram till Efrat, kom Rakel i barnsnöd, och barnsnöden blev henne svår.
Då nu hennes barnsnöd var som svårast, sade hjälpkvinnan till henne: »Frukta icke; ty också denna gång får du en son.»
Men när hon höll på att giva upp andan, ty hon skulle nu dö, gav hon honom namnet Ben-Oni ; men hans fader kallade honom Benjamin .
Så dog Rakel, och hon blev begraven vid vägen till Efrat, det är Bet-Lehem.
Och Jakob reste en vård på hennes grav; det är den som ännu i dag kallas Rakels gravvård.
Och Israel bröt upp därifrån och slog upp sitt tält på andra sidan om Herdetornet.
Och medan Israel bodde där i landet, gick Ruben åstad och lägrade Bilha, sin faders bihustru; och Israel fick höra det.
Och Jakob hade tolv söner.
Leas söner voro Ruben, Jakobs förstfödde, vidare Simeon, Levi, Juda, Isaskar och Sebulon.
Rakels söner voro Josef och Benjamin.
Bilhas, Rakels tjänstekvinnas, söner voro Dan och Naftali.
Silpas, Leas tjänstekvinnas, söner voro Gad och Aser.
Dessa voro Jakobs söner, och de föddes åt honom i Paddan-Aram.
Och Jakob kom till sin fader Isak i Mamre vid Kirjat-Arba, det är Hebron, där Abraham och Isak hade bott såsom främlingar.
Och Isak levde ett hundra åttio år;
därefter gav Isak upp andan och dog och blev samlad till sina fäder, gammal och mätt på att leva.
Och hans söner Esau och Jakob begrovo honom.
Detta är berättelsen om Esaus, det är Edoms, släkt.
Esau hade tagit sina hustrur bland Kanaans döttrar: Ada, hetiten Elons dotter, och Oholibama, dotter till Ana och sondotter till hivéen Sibeon,
så ock Basemat, Ismaels dotter, Nebajots syster.
Och Ada födde Elifas åt Esau, men Basemat födde Reguel.
Och Oholibama födde Jeus, Jaelam och Kora.
Dessa voro Esaus söner, vilka föddes åt honom i Kanaans land.
Och Esau tog sina hustrur, sina söner och döttrar och allt sitt husfolk, sin boskap och alla sina dragare och all annan egendom som han hade förvärvat i Kanaans land och drog till ett annat land och skilde sig så från sin broder Jakob.
Ty deras ägodelar voro så stora att de icke kunde bo tillsammans; landet där de uppehöllo sig räckte icke till åt dem, för deras boskapshjordars skull.
Och Esau bosatte sig i Seirs bergsbygd.
Esau, det är densamme som Edom.
Och detta är berättelsen om Esaus släkt, hans som var stamfader för edoméerna, i Seirs bergsbygd.
Dessa äro namnen på Esaus söner: Elifas, son till Ada, Esaus hustru, och Reguel, son till Basemat, Esaus hustru.
Men Elifas' söner voro Teman, Omar, Sefo, Gaetam och Kenas.
Och Timna, som var Elifas', Esaus sons, bihustru, födde Amalek åt Elifas.
Dessa voro söner till Ada, Esaus hustru.
Men Reguels söner voro dessa: Nahat och Sera, Samma och Missa.
Dessa voro söner till Basemat, Esaus hustru.
Men söner till Oholibama, Esaus hustru, dotter till Ana och sondotter till Sibeon, voro dessa, som hon födde åt Esau: Jeus, Jaelam och Kora.
Dessa voro stamfurstarna bland Esaus söner: Elifas', Esaus förstföddes, söner voro dessa: fursten Teman, fursten Omar, fursten Sefo, fursten Kenas,
fursten Kora, fursten Gaetam, fursten Amalek.
Dessa voro de furstar som härstammade från Elifas, i Edoms land; dessa voro Adas söner.
Och dessa voro Reguels, Esaus sons, söner: fursten Nahat, fursten Sera, fursten Samma, fursten Missa.
Dessa voro de furstar som härstammade från Reguel, i Edoms land; dessa voro söner till Basemat, Esaus hustru.
Och dessa voro Oholibamas, Esaus hustrus, söner: fursten Jeus, fursten Jaelam, fursten Kora.
Dessa voro de furstar som härstammade från Oholibama, Anas dotter och Esaus hustru.
Dessa voro Esaus söner, och dessa deras stamfurstar.
Han är densamme som Edom.
Dessa voro horéen Seirs söner, landets förra inbyggare: Lotan, Sobal, Sibeon, Ana,
Dison, Eser och Disan.
Dessa voro horéernas, Seirs söners, stamfurstar i Edoms land.
Men Lotans söner voro Hori och Hemam; och Lotans syster var Timna.
Och dessa voro Sobals söner: Alvan, Manahat och Ebal, Sefo och Onam.
Och dessa voro Sibeons söner: Aja och Ana; det var denne Ana som fann de varma källorna i öknen, när han vaktade sin fader Sibeons åsnor.
Men dessa voro Anas barn: Dison och Oholibama, Anas dotter.
Och dessa voro Disans söner: Hemdan, Esban, Jitran och Keran.
Och dessa voro Esers söner: Bilhan, Saavan och Akan.
Dessa voro Disans söner: Us och Aran.
Dessa voro horéernas stamfurstar: fursten Lotan, fursten Sobal, fursten Sibeon, fursten Ana,
fursten Dison, fursten Eser, fursten Disan.
Dessa voro horéernas stamfurstar i Seirs land, var furste för sig.
Och dessa voro de konungar som regerade i Edoms land, innan ännu någon israelitisk konung var konung där:
Bela, Beors son, var konung i Edom, och hans stad hette Dinhaba.
När Bela dog, blev Jobab, Seras son, från Bosra, konung efter honom.
När Jobab dog, blev Husam från temanéernas land konung efter honom.
När Husam dog, blev Hadad, Bedads son, konung efter honom, han som slog midjaniterna på Moabs mark; och hans stad hette Avit.
När Hadad dog, blev Samla från Masreka konung efter honom.
När Samla dog, blev Saul från Rehobot vid floden konung efter honom.
När Saul dog, blev Baal-Hanan, Akbors son, konung efter honom.
När Baal-Hanan, Akbors son, dog, blev Hadar konung efter honom; och hans stad hette Pagu, och hans hustru hette Mehetabel, dotter till Matred, som var dotter till Me-Sahab.
Och dessa äro namnen på Esaus stamfurstar, efter deras släkter och orter, med deras namn: fursten Timna, fursten Alva, fursten Jetet,
fursten Oholibama, fursten Ela, fursten Pinon,
fursten Kenas, fursten Teman, fursten Mibsar,
fursten Magdiel, fursten Iram.
Dessa voro Edoms stamfurstar, efter deras boningsorter i det land de hade tagit i besittning -- hans som ock kallas Esau, edoméernas stamfader.
Men Jakob bosatte sig i det land där hans fader hade bott såsom främling, nämligen i Kanaans land.
Detta är berättelsen om Jakobs släkt.
När Josef var sjutton år gammal, gick han, jämte sina bröder, i vall med fåren; han följde då såsom yngling med Bilhas och Silpas, sin faders hustrurs, söner.
Och Josef bar fram till deras fader vad ont som sades om dem.
Men Israel hade Josef kärare än alla sina andra söner, eftersom han hade fött honom på sin ålderdom; och han lät göra åt honom en fotsid livklädnad.
Då nu hans bröder sågo att deras fader hade honom kärare än alla hans bröder, blevo de hätska mot honom och kunde icke tala vänligt till honom.
Därtill hade Josef en gång en dröm, som han omtalade för sina bröder; sedan hatade de honom ännu mer.
Han sade nämligen till dem: »Hören vilken dröm jag har haft.
Jag tyckte att vi bundo kärvar på fältet; och se, min kärve reste sig upp och blev stående, och edra kärvar ställde sig runt omkring och bugade sig för min kärve.»
Då sade hans bröder till honom: »Skulle du bliva vår konung, och skulle du råda över oss?»
Och de hatade honom ännu mer för hans drömmars skull och för vad han hade sagt.
Sedan hade han ännu en annan dröm som han förtäljde för sina bröder; han sade: »Hören, jag har haft ännu en dröm.
Jag tyckte att solen och månen och elva stjärnor bugade sig för mig.»
När han förtäljde detta för sin fader och sina bröder, bannade hans fader honom och sade till honom: »Vad är detta för en dröm som du har haft?
Skulle då jag och din moder och dina bröder komma och buga oss ned till jorden för dig?»
Och hans bröder avundades honom; men hans fader bevarade detta i sitt minne.
Då nu en gång hans bröder hade gått bort för att vakta sin faders får i Sikem,
sade Israel till Josef: »Se, dina bröder vakta fåren i Sikem; gör dig redo, jag vill sända dig till dem.»
Han svarade honom: »Jag är redo.»
Då sade han till honom: »Gå och se efter, om det står väl till med dina bröder, och om det står väl till med fåren, och kom tillbaka till mig med svar.»
Så sände han honom åstad från Hebrons dal, och han kom till Sikem.
Där mötte han en man, medan han gick omkring villrådig på fältet; och mannen frågade honom: »Vad söker du?»
Han svarade: »Jag söker efter mina bröder; säg mig var de vakta sin hjord.»
Mannen svarade: »De hava brutit upp härifrån; ty jag hörde dem säga: 'Låt oss gå till Dotain.'»
Då gick Josef vidare efter sina bröder och fann dem i Dotan.
När de nu på avstånd fingo se honom, innan han ännu hade hunnit fram till dem, lade de råd om att döda honom.
De sade till varandra: »Se, där kommer drömmaren.
Upp, låt oss dräpa honom och kasta honom i en brunn; sedan kunna vi säga att ett vilddjur har ätit upp honom.
Så få vi se huru det går med hans drömmar.»
Men när Ruben hörde detta, ville han rädda honom undan deras händer och sade: »Låt oss icke slå ihjäl honom.»
Ytterligare sade Ruben till dem: »Utgjuten icke blod; kasten honom i brunnen här i öknen, men bären icke hand på honom.»
Han ville nämligen rädda honom undan deras händer och föra honom tillbaka till hans fader.
Då nu Josef kom fram till sina bröder, togo de av honom hans livklädnad, den fotsida klädnaden som han hade på sig,
och grepo honom och kastade honom i brunnen; men brunnen var tom, intet vatten fanns däri.
Därefter satte de sig ned för att äta.
När de då lyfte upp sina ögon, fingo de se ett tåg av ismaeliter komma från Gilead, och deras kameler voro lastade med dragantgummi, balsam och ladanum; de voro på väg med detta ned till Egypten.
Då sade Juda till sina bröder: »Vad gagn hava vi därav att vi dräpa vår broder och dölja hans blod?»
Nej, låt oss sälja honom till ismaeliterna; må vår hand icke komma vid honom, ty han är ju vår broder, vårt eget kött.»
Och hans bröder lydde honom.
Då nu midjanitiska köpmän kommo där förbi, drogo de upp Josef ur brunnen; och de sålde Josef för tjugu siklar silver till ismaeliterna.
Dessa förde så Josef till Egypten.
När sedan Ruben kom tillbaka till brunnen, se, då fanns Josef icke i brunnen.
Då rev han sönder sina kläder
och vände tillbaka till sina bröder och sade: »Gossen är icke där, vart skall jag nu taga vägen?»
Men de togo Josefs livklädnad och slaktade en bock och doppade klädnaden i blodet;
därefter sände de den fotsida livklädnaden hem till sin fader och läto säga: »Denna har vi funnit; se efter, om det är din sons livklädnad eller icke.»
Och han kände igen den och sade: »Det är min sons livklädnad; ett vilddjur har ätit upp honom, förvisso är Josef ihjälriven.»
Och Jakob rev sönder sina kläder och svepte säcktyg om sina länder och sörjde sin son i lång tid.
Och alla hans söner och alla hans döttrar kommo för att trösta honom; men han ville icke låta trösta sig, utan sade: »Jag skall med sorg fara ned i dödsriket till min son.»
Så begrät hans fader honom.
Men medaniterna förde honom till Egypten och sålde honom till Potifar, som var hovman hos Farao och hövitsman för drabanterna.
Vid den tiden begav sig Juda åstad bort ifrån sina bröder och slöt sig till en man i Adullam, som hette Hira.
Där fick Juda se dottern till en kananeisk man som hette Sua, och han tog henne till sig och gick in till henne.
Och hon blev havande och födde en son, och han fick namnet Er.
Åter blev hon havande och födde en son och gav honom namnet Onan.
Och hon födde ännu en son, och åt denne gav hon namnet Sela; och när han föddes, var Juda i Kesib.
Och Juda tog åt Er, sin förstfödde, en hustru som hette Tamar.
Men Er, Judas förstfödde, misshagade HERREN; därför dödade HERREN honom.
Då sade Juda till Onan: »Gå in till din broders hustru, äkta henne i din broders ställe och skaffa avkomma åt din broder.»
Men eftersom Onan visste att avkomman icke skulle bliva hans egen, lät han, när han gick in till sin broders hustru, det spillas på jorden, för att icke giva avkomma åt sin broder.
Men det misshagade HERREN att han gjorde så; därför dödade han också honom.
Då sade Juda till sin sonhustru Tamar: »Stanna såsom änka i din faders hus, till dess min son Sela bliver fullvuxen.»
Han fruktade nämligen att annars också denne skulle dö, likasom hans bröder.
Så gick Tamar bort och stannade i sin faders hus.
En lång tid därefter dog Suas dotter, Judas hustru.
Och efter sorgetidens slut gick Juda med sin vän adullamiten Hira upp till Timna, för att se efter dem som klippte hans får.
När man nu berättade för Tamar att hennes svärfader gick upp till Timna för att klippa sina får,
lade hon av sig sina änkekläder och betäckte sig med en slöja och höljde in sig och satte sig vid porten till Enaim på vägen till Timna.
Ty hon såg, att fastän Sela var fullvuxen, blev hon likväl icke given åt honom till hustru.
Då nu Juda fick se henne, trodde han att hon var en sköka; hon hade ju nämligen sitt ansikte betäckt.
Och han vek av till henne, där hon satt vid vägen, och sade: »Kom, låt mig gå in till dig.»
Ty han visste icke att det var hans sonhustru.
Hon svarade: »Vad vill du giva mig för att få gå in till mig?»
Han sade: »Jag vill sända dig en killing ur min hjord.»
Hon svarade: »Ja, om du giver mig pant, till dess du sänder den.»
Han sade: »Vad skall jag då giva dig i pant?»
Hon svarade: »Din signetring, din snodd och staven som du har i din hand.»
Då gav han henne detta och gick in till henne, och hon blev havande genom honom.
Och hon stod upp och gick därifrån och lade av sin slöja och klädde sig åter i sina änkekläder.
Och Juda sände killingen med sin vän adullamiten, för att få igen panten av kvinnan; men denne fann henne icke.
Och han frågade folket där på orten och sade: »Var är tempeltärnan, hon som satt i Enaim vid vägen?»
De svarade: »Här har ingen tempeltärna varit.»
Och han kom tillbaka till Juda och sade: »Jag har icke funnit henne; därtill säger folket på orten att ingen tempeltärna har varit där.»
Då sade Juda: »Må hon då behålla det, så att vi icke draga smälek över oss.
Jag har nu sänt killingen, men du har icke funnit henne.»
Vid pass tre månader därefter blev så berättat för Juda: »Din sonhustru Tamar har bedrivit otukt, och i otukt har hon blivit havande.»
Juda sade: »Fören ut henne till att brännas.»
Men när hon fördes ut, sände hon bud till sin svärfader och lät säga: »Genom en man som är ägare till detta har jag blivit havande.»
Och hon lät säga: »Se efter, vem denna signetring, dessa snodder och denna stav tillhöra.»
Och Juda kände igen dem och sade: »Hon är i sin rätt mot mig, eftersom jag icke har givit henne åt min son Sela.»
Men han kom icke mer vid henne.
När hon nu skulle föda, se, då funnos tvillingar i hennes liv.
Och i födslostunden stack den ene fram en hand; då tog hjälpkvinnan en röd tråd och band den om hans hand och sade: »Denne kom först fram.»
Men när han därefter åter drog sin hand tillbaka, se, då kom hans broder fram; och hon sade: »Varför har du trängt dig fram?»
Och han fick namnet Peres .
Därefter kom hans broder fram, han som hade den röda tråden om sin hand, och han fick namnet Sera.
Och Josef fördes ned till Egypten; och Potifar, som var hovman hos Farao och hövitsman för drabanterna, en egyptisk man, köpte honom av ismaeliterna som hade fört honom ditned.
Och HERREN var med Josef, så att han blev en lyckosam man.
Och han vistades i sin herres, egyptierns, hus;
och hans herre såg att HERREN var med honom, ty allt vad han gjorde lät HERREN lyckas väl under hans hand.
Och Josef fann nåd för hans ögon och fick betjäna honom.
Och han satte honom över sitt hus, och allt vad han ägde lämnade han i hans vård.
Och från den stund då han hade satt honom över sitt hus och över allt vad han ägde, välsignade HERREN egyptierns hus, för Josefs skull; och HERRENS välsignelse vilade över allt vad han ägde, hemma och på marken.
Därför överlät han i Josefs vård allt vad han ägde, och sedan han hade fått honom till sin hjälp, bekymrade han sig icke om något, utom maten som han själv åt.
Men Josef hade en skön gestalt och var skön att skåda.
Och efter en tid hände sig att hans herres hustru kastade sina ögon på Josef och sade: »Ligg hos mig.»
Men han ville icke, utan sade till sin herres hustru: »Se, alltsedan min herre har tagit mig till sin hjälp, bekymrar han sig icke om något i huset, och allt vad han äger har han lämnat i min vård.
Han har i detta hus icke större makt än jag, och intet annat har han förbehållit sig än dig allena, eftersom du är hans hustru.
Huru skulle jag då kunna göra så mycket ont och synda mot Gud?»
Och fastän hon talade sådant dag efter dag till Josef, hörde han dock icke på henne och ville icke ligga hos henne eller vara med henne.
Men en dag då han kom in i huset för att förrätta sina sysslor, och ingen av husfolket var tillstädes därinne,
fattade hon honom i manteln och sade: »Ligg hos mig.»
Men han lämnade manteln i hennes hand och flydde och kom ut.
Då hon nu såg att han hade lämnat sin mantel i hennes hand och flytt ut,
ropade hon på sitt husfolk och sade till dem: »Sen här, han har fört hit till oss en hebreisk man, för att denne skulle locka oss till lättfärdighet.
Han kom in till mig och ville ligga hos mig; men jag ropade med hög röst.
Och när han hörde att jag hov upp min röst och ropade, lämnade han sin mantel kvar hos mig och flydde och kom ut.»
Och hon lät hans mantel ligga kvar hos sig, till dess hans herre kom hem;
då berättade hon för honom detsamma; hon sade: »Den hebreiske tjänaren som du har fört hit till oss kom in till mig, och ville locka mig till lättfärdighet.
Men då jag hov upp min röst och ropade, lämnade han sin mantel kvar hos mig och flydde ut.»
När nu hans herre hörde vad hans hustru berättade för honom, nämligen att hans tjänare hade betett sig mot henne på detta sätt, blev hans vrede upptänd.
Och Josefs herre tog honom och lät sätta honom i det fängelse där konungens fångar sutto fängslade; där fick han då vara i fängelse.
Men HERREN var med Josef och förskaffade honom ynnest och lät honom finna nåd hos föreståndaren för fängelset.
Och föreståndaren för fängelset lät alla fångar som sutto i fängelset stå under Josefs uppsikt; och allt vad där skulle göras, det gjordes genom honom.
Föreståndaren för fängelset tog sig alls icke av något som Josef hade om hand, eftersom HERREN var med denne; och vad han gjorde, det lät HERREN lyckas väl.
En tid härefter hände sig att den egyptiske konungens munskänk och hans bagare försyndade sig mot sin herre, konungen av Egypten.
Och Farao blev förtörnad på sina två hovmän, överste munskänken och överste bagaren,
och lät sätta dem i förvar i drabanthövitsmannens hus, i samma fängelse där Josef satt fången.
Och hövitsmannen för drabanterna anställde Josef hos dem till att betjäna dem; och de sutto där i förvar en tid.
Medan nu den egyptiske konungens munskänk och bagare sutto fångna i fängelset, hade de båda under samma natt var sin dröm, vardera med sin särskilda betydelse.
Och när Josef om morgonen kom in till dem, fick han se att de voro bedrövade.
Då frågade han Faraos hovmän, som med honom sutto i förvar i hans herres hus: »Varför sen I så sorgsna ut i dag?»
De svarade honom: »Vi hava haft en dröm, och ingen finnes, som kan uttyda den.»
Josef sade till dem: »Att giva uttydningen är ju Guds sak; förtäljen drömmen för mig.»
Då förtäljde överste munskänken sin dröm för Josef och sade till honom: »Jag drömde att ett vinträd stod framför mig;
på vinträdet voro tre rankor, och knappt hade det skjutit skott, så slogo dess blommor ut och dess klasar buro mogna druvor.
Och jag hade Faraos bägare i min hand, och jag tog druvorna och pressade ut dem i Faraos bägare och gav Farao bägaren i handen.»
Då sade Josef till honom: »Detta är uttydningen: de tre rankorna betyda tre dagar;
om tre dagar skall Farao upphöja ditt huvud och sätta dig åter på din plats, så att du får giva Farao bägaren i handen likasom förut, då du var hans munskänk.
Men tänk på mig, när det går dig väl, så att du gör barmhärtighet med mig och nämner om mig för Farao och skaffar mig ut från detta hus;
ty jag är med orätt bortförd från hebréernas land, och icke heller här har jag gjort något varför jag borde sättas i fängelse.»
Då nu överste bagaren såg att Josef hade givit en god uttydning, sade han till honom: »Också jag hade en dröm.
Jag tyckte att jag bar tre vetebrödskorgar på mitt huvud.
Och i den översta korgen funnos bakverk av alla slag, sådant som Farao plägar äta; men fåglarna åto därav ur korgen på mitt huvud.»
Då svarade Josef och sade: »Detta är uttydningen: de tre korgarna betyda tre dagar;
om tre dagar skall Farao upphöja ditt huvud och taga det av dig; han skall upphänga dig på trä, och fåglarna skola äta ditt kött.»
På tredje dagen därefter, då det var Faraos födelsedag, gjorde denne ett gästabud för alla sina tjänare.
Då upphöjde han, bland sina tjänare, såväl överste munskänkens huvud som överste bagarens.
Han insatte överste munskänken åter i hans ämbete, så att han fick giva Farao bägaren i handen;
men överste bagaren lät han upphänga, såsom Josef hade sagt dem i sin uttydning.
Men överste munskänken tänkte icke på Josef, utan glömde honom.
Två år därefter hände sig att Farao hade en dröm.
Han tyckte sig stå vid Nilfloden.
Och han såg sju kor, vackra och feta, stiga upp ur floden, och de betade i vassen.
Sedan såg han sju andra kor, fula och magra, stiga upp ur floden; och de ställde sig bredvid de förra korna på stranden av floden.
Och de fula och magra korna åto upp de sju vackra och feta korna.
Därefter vaknade Farao.
Men han somnade åter in och såg då i drömmen sju ax, frodiga och vackra, växa på samma strå.
Sedan såg han sju andra ax skjuta upp, tunna och svedda av östanvinden;
och de tunna axen uppslukade de sju frodiga och fulla axen.
Därefter vaknade Farao och fann att det var en dröm.
Då han nu om morgonen var orolig till sinnes, sände han ut och lät kalla till sig alla spåmän och alla vise i Egypten.
Och Farao förtäljde sina drömmar för dem; men ingen fanns, som kunde uttyda dem för Farao.
Då talade överste munskänken till Farao och sade: »Jag måste i dag påminna om mina synder.
När Farao en gång var förtörnad på sina tjänare, satte han mig jämte överste bagaren i fängelse i drabanthövitsmannens hus.
Då hade vi båda, jag och han, under samma natt en dröm, och våra drömmar hade var sin särskilda betydelse.
Och jämte oss var där en ung hebré, som var tjänare hos hövitsmannen för drabanterna.
För honom förtäljde vi våra drömmar, och han uttydde dem för oss; efter som var och en hade drömt gav han en uttydning.
Och såsom han uttydde för oss, så gick det.
Jag blev åter insatt på min plats, och den andre blev upphängd.»
Då sände Farao och lät kalla Josef till sig; och man skyndade att föra honom ut ur fängelset.
Och han lät raka sig och bytte om kläder och kom inför Farao.
Och Farao sade till Josef: »Jag har haft en dröm, och ingen finnes, som kan uttyda den.
Men jag har hört sägas om dig, att allenast du får höra en dröm, kan du uttyda den.»
Josef svarade Farao och sade: »I min makt står det icke; men Gud skall giva Farao ett lyckosamt svar.»
Då sade Farao till Josef: »Jag drömde att jag stod på stranden av Nilfloden.
Och jag såg sju kor stiga upp ur floden, feta och vackra, och de betade i vassen.
Sedan såg jag sju andra kor stiga upp, avfallna och mycket fula och magra; i hela Egyptens land har jag icke sett några så fula som dessa.
Och de magra och fula korna åto upp de sju första, feta korna.
Men när de hade sväljt ned dem, kunde man icke märka att de hade sväljt ned dem, utan de förblevo fula såsom förut.
Därefter vaknade jag.
Åter drömde jag och såg då sju ax, fulla och vackra, växa på samma strå.
Sedan såg jag sju andra ax skjuta upp, förtorkade, tunna och svedda av östanvinden;
och de tunna axen uppslukade de sju vackra axen.
Detta omtalade jag för spåmännen; men ingen fanns, som kunde förklara det för mig.»
Då sade Josef till Farao: »Faraos drömmar hava en och samma betydelse; vad Gud ämnar göra, det har han förkunnat för Farao.
De sju vackra korna betyda sju år, de sju vackra axen betyda ock sju år; drömmarna hava en och samma betydelse.
Och de sju magra och fula korna som stego upp efter dessa betyda sju år, så ock de sju tomma axen, de som voro svedda av östanvinden; sju hungerår skola nämligen komma.
Detta menade jag, när jag sade till Farao: Vad Gud ämnar göra, det har han låtit Farao veta.
Se, sju år skola komma med stor ymnighet över hela Egyptens land.
Men efter dem skola sju hungerår inträffa, sådana, att man skall förgäta all den förra ymnigheten i Egyptens land, och hungersnöden skall förtära landet.
Och man skall icke hava något minne av den förra ymnigheten i landet, för den hungersnöds skull som sedan kommer, ty den skall bliva mycket svår.
Men att Farao har haft drömmen två gånger, det betyder att detta är av Gud bestämt, och att Gud skall låta det ske snart.
Må nu alltså Farao utse en förståndig och vis man, som han kan sätta över Egyptens land.
Må Farao göra så; må han ock förordna tillsyningsmän över landet och taga upp femtedelen av avkastningen i Egyptens land under de sju ymniga åren.
Må man under dessa kommande goda år samla in allt som kan tjäna till föda och hopföra säd under Faraos vård i städerna, för att tjäna till föda, och må man sedan förvara den,
så att dessa födoämnen finnas att tillgå för landet under de sju hungerår som skola komma över Egyptens land.
Så skall landet icke behöva förgås genom hungersnöden.»
Det talet behagade Farao och alla hans tjänare.
Och Farao sade till sina tjänare: »Kunna vi finna någon i vilken Guds Ande så är som i denne?»
Och Farao sade till Josef: »Eftersom Gud har kungjort för dig allt detta, finnes ingen som är så förståndig och vis som du.
Du skall förestå mitt hus, och efter dina befallningar skall allt mitt folk rätta sig; allenast däri att tronen förbliver min vill jag vara förmer än du.»
Ytterligare sade Farao till Josef: »Jag sätter dig nu över hela Egyptens land.»
Och Farao tog ringen av sin hand och satte den på Josefs hand och lät kläda honom i kläder av fint linne och hängde den gyllene kedjan om hans hals.
Och han lät honom åka i vagnen närmast efter sin egen, och man utropade framför honom »abrek ».
Och han satte honom över hela Egyptens land.
Och Farao sade till Josef: »Jag är Farao; utan din vilja skall ingen i hela Egyptens land lyfta hand eller fot.»
Och Farao gav Josef namnet Safenat-Panea och gav honom till hustru Asenat, dotter till Poti-Fera, prästen i On.
Och Josef begav sig ut och besåg Egyptens land.
Josef var trettio år gammal, när han stod inför Farao, konungen i Egypten.
Och Josef gick ut ifrån Farao och färdades omkring i hela Egyptens land.
Och landet gav under de sju ymniga åren avkastning i överflöd
och under dessa sju år som kommo i Egyptens land samlade han in allt som kunde tjäna till föda och lade upp det i städerna.
I var särskild stad lade han upp de födoämnen som man hämtade ifrån fälten däromkring.
Så hopförde Josef säd i stor myckenhet, såsom sanden i havet, till dess man måste upphöra att hålla räkning på den, eftersom det var omöjligt att hålla räkning på den.
Och åt Josef föddes två söner, innan något hungerår kom; de föddes åt honom av Asenat, dotter till Poti-Fera, prästen i On.
Och Josef gav åt den förstfödde namnet Manasse , »ty», sade han, »Gud har låtit mig förgäta all min olycka och hela min faders hus.»
Och åt den andre gav han namnet Efraim , »ty», sade han, »Gud har gjort mig fruktsam i mitt lidandes land».
Men de sju ymniga åren som först hade kommit i Egyptens land gingo till ända;
sedan begynte de sju hungeråren, såsom Josef hade förutsagt.
Och hungersnöd uppstod i alla andra länder; men i Egyptens land fanns bröd överallt.
Och när hela Egyptens land begynte hungra och folket ropade till Farao efter bröd, sade Farao till alla egyptier: »Gån till Josef, och gören vad han säger eder.»
När nu alltså hungersnöd var över hela landet, öppnade Josef alla förrådshus och sålde säd åt egyptierna.
Men hungersnöden blev allt större i Egyptens land;
och från alla länder kom man till Josef i Egypten för att köpa säd, ty hungersnöden blev allt större i alla länder.
Men när Jakob förnam att säd fanns i Egypten, sade han till sina söner: »Varför stån I så rådlösa?»
Och han sade vidare: »Se, jag har hört att i Egypten finnes säd; faren ditned och köpen därifrån säd åt oss, för att vi må leva och icke dö.»
Då foro tio av Josefs bröder ned för att köpa säd i Egypten.
Men Benjamin, Josefs broder, blev icke av Jakob sänd åstad med sina bröder, ty han fruktade att någon olycka kunde hända honom.
Så kommo då, bland de andra, också Israels söner för att köpa säd; ty hungersnöd rådde i Kanaans land.
Och Josef var den som hade att befalla i landet; det var han som sålde säd åt allt folket i landet.
Då nu Josefs bröder kommo dit, föllo de ned till jorden på sitt ansikte inför honom.
När då Josef fick se sina bröder, kände han igen dem; men han ställde sig främmande mot dem och tilltalade dem hårt och frågade dem: »Varifrån kommen I?»
De svarade: »Från Kanaans land, för att köpa säd till föda åt oss.»
Och fastän Josef kände igen sina bröder, kände de icke igen honom.
Men Josef tänkte på de drömmar som han hade drömt om dem.
Och han sade till dem: »I ären spejare, I haven kommit för att se efter, var landet är utan skydd.»
De svarade honom: »Nej, herre, dina tjänare hava kommit för att köpa säd till föda åt sig.
Vi äro alla söner till en och samma man; vi äro redliga män, dina tjänare äro inga spejare.»
Men han sade till dem: »Jo, I haven kommit för att se efter, var landet är utan skydd.»
De svarade: »Vi, dina tjänare, äro tolv bröder, söner till en och samma man i Kanaans land; men den yngste är nu hemma hos vår fader, och en är icke mer till.»
Josef sade till dem: »Det är såsom jag sade eder: I ären spejare.
Och på detta sätt vill jag pröva eder: så sant Farao lever, I skolen icke slippa härifrån, med mindre eder yngste broder kommer hit.
En av eder må fara och hämta hit eder broder.
Men I andra skolen stanna såsom fångar, för att jag så må pröva om I haven talat sanning.
Ty om så icke är, då ären I spejare, så sant Farao lever.»
Därefter lät han hålla dem allasammans i fängelse under tre dagar.
Men på tredje dagen sade Josef till dem: »Om I viljen leva, så gören på detta sätt, ty jag fruktar Gud:
ären I redliga män, så må en av eder, I bröder, stanna såsom fånge i huset där I haven suttit fängslade; men I andra mån fara eder väg, och föra hem med eder den säd som I haven köpt till hjälp mot hungersnöden hemma hos eder.
Fören sedan eder yngste broder hit till mig; om så edra ord visa sig vara sanna, skolen I slippa att dö.»
Och de måste göra så.
Men de sade till varandra: »Förvisso hava vi dragit skuld över oss genom det som vi gjorde mot vår broder; ty vi sågo hans själs ångest, när han bad oss om misskund, och vi ville dock icke lyssna till honom.
Därför hava vi själva kommit i denna ångest.»
Ruben svarade dem: »Sade jag icke till eder: 'Försynden eder icke på gossen'?
Men I lyssnaden icke till mig; se, därför utkräves nu hans blod.»
Men de visste icke att Josef förstod detta, ty han talade med dem genom tolk.
Och han vände sig bort ifrån dem och grät.
Sedan vände han sig åter till dem och talade med dem; och han tog Simeon ut ur deras krets och lät fängsla honom inför deras ögon.
Och Josef bjöd att man skulle fylla deras säckar med säd, och lägga vars och ens penningar tillbaka i hans säck, och giva dem kost för resan.
Och man gjorde så med dem.
Och de lastade säden på sina åsnor och foro därifrån.
Men när vid ett viloställe en av dem öppnade sin säck för att giva foder åt sin åsna, fick han se sina penningar ligga överst i säcken.
Då sade han till sina bröder: »Mina penningar hava blivit lagda hit tillbaka; se, de äro här i min säck.»
Då blevo de utom sig av häpnad och sågo förskräckta på varandra och sade: »Vad har Gud gjort mot oss!»
När de kommo hem till sin fader Jakob i Kanaans land, berättade de för honom allt vad som hade hänt dem och sade:
»Mannen som var herre där i landet tilltalade oss hårt och behandlade oss såsom om vi ville bespeja landet.
Men vi sade till honom: 'Vi äro redliga män och inga spejare;
vi äro tolv bröder, samma faders söner; en är icke mer till, och den yngste är nu hemma hos vår fader i Kanaans land.'
Men mannen som var herre i landet svarade oss: 'Därav skall jag veta att I ären redliga män: lämnen kvar hos mig en av eder, I bröder; tagen så vad I haven köpt till hjälp mot hungersnöden hemma hos eder, och faren eder väg.
Sedan mån I föra eder yngste broder hit till mig, så kan jag veta att I icke ären spejare, utan redliga män.
Då skall jag giva eder broder tillbaka åt eder, och I skolen fritt få draga omkring i landet.
När de sedan tömde sina säckar, fann var och en sin penningpung i sin säck.
Och då de och deras fader fingo se penningpungarna, blevo de förskräckta.
Och Jakob, deras fader, sade till dem: »I gören mig barnlös; Josef är borta, Simeon är borta, Benjamin viljen I ock taga ifrån mig; över mig kommer allt detta.»
Då svarade Ruben sin fader och sade: »Mina båda söner må du döda, om jag icke för honom åter till dig.
Anförtro honom åt mig, jag skall föra honom tillbaka till dig.»
Men han svarade: »Min son får icke fara ditned med eder.
Hans broder är ju död, och han är allena kvar; om nu någon olycka hände honom på den resa I viljen företaga, så skullen I bringa mina grå hår med sorg ned i dödsriket.»
Men hungersnöden var svår i landet.
Och när de hade förtärt den säd som de hade hämtat från Egypten, sade deras fader till dem: »Faren tillbaka och köpen litet säd till föda åt oss.»
Men Juda svarade honom och sade: »Mannen betygade högtidligt och sade till oss: 'I fån icke komma inför mitt ansikte, med mindre eder broder är med eder.'
Om du nu låter vår broder följa med oss, så skola vi fara ned och köpa säd till föda åt dig.
Men om du icke låter honom följa med oss, så vilja vi icke fara, ty mannen sade till oss: 'I fån icke komma inför mitt ansikte, med mindre eder broder är med eder.'
Då sade Israel: »Varför gjorden I så illa mot mig och berättaden för mannen att I haden ännu en broder?»
De svarade: »Mannen frågade noga om oss och vår släkt; han sade: 'Lever eder fader ännu?
Haven I någon broder?'
Då omtalade vi för honom huru det förhöll sig.
Kunde vi veta att han skulle säga: 'Fören eder broder hitned'?»
Och Juda sade till sin fader Israel: »Låt ynglingen följa med mig, så vilja vi stå upp och begiva oss åstad, för att vi må leva och icke dö, vi själva och du och våra kvinnor och barn.
Jag vill ansvara för honom; av min hand må du utkräva honom.
Om jag icke för honom åter till dig och ställer honom inför ditt ansikte, så vill jag vara en syndare inför dig i all min tid.
Sannerligen, om vi icke hade dröjt så länge, så skulle vi redan hava varit tillbaka för andra gången.»
Då svarade deras fader Israel dem: »Måste det så vara, så gören nu på detta sätt: tagen av landets bästa frukt i edra säckar och fören det till mannen såsom skänk, litet balsam och litet honung, dragantgummi och ladanum, pistacienötter och mandlar.
Och tagen dubbla summan penningar med eder, så att I fören tillbaka dit med eder de penningar som I haven fått igen överst i edra säckar.
Kanhända var det ett misstag.
Tagen ock eder broder med eder, och stån upp och faren tillbaka till mannen.
Men Gud den Allsmäktige låte eder finna barmhärtighet inför mannen, så att han tillstädjer eder andre broder och Benjamin att återvända med eder.
Men skall jag bliva barnlös, så må det då ske.»
Då togo männen de nämnda skänkerna och togo med sig dubbla summan penningar, därtill ock Benjamin, och stodo upp och foro ned till Egypten och trädde inför Josef.
Då nu Josef såg att Benjamin var med dem, sade han till sin hovmästare: »För dessa män in i mitt hus; och låt slakta och tillreda en måltid, ty männen skola äta middag med mig.»
Och mannen gjorde såsom Josef hade sagt och förde männen in i Josefs hus.
Och männen blevo förskräckta, när de fördes in i Josefs hus; de sade: »Det är på grund av penningarna vi föras hitin, de penningar som förra gången kommo tillbaka i våra säckar; ty han vill nu störta sig på oss och överfalla oss och göra oss själva till trälar och taga ifrån oss våra åsnor.»
Och de trädde fram till Josefs hovmästare och talade med honom vid ingången till huset
och sade: »Hör oss, herre.
När vi förra gången voro härnere för att köpa säd till föda åt oss
och sedan kommo till ett viloställe och öppnade våra säckar, då fann var och en av oss sina penningar överst i sin säck, penningarna till deras fulla vikt; dem hava vi nu fört tillbaka med oss.
Och vi hava tagit andra penningar med oss för att köpa säd till föda åt oss.
Vi veta icke vem som hade lagt penningarna i våra säckar.»
Då svarade han: »Varen vid gott mod, frukten icke; det är eder Gud och eder faders Gud som har låtit eder finna en skatt i edra säckar; edra penningar har jag fått.»
Sedan hämtade han Simeon ut till dem.
Och han förde männen in i Josefs hus och gav dem vatten till att två sina fötter och gav foder åt deras åsnor.
Och de ställde i ordning sina skänker, till dess Josef skulle komma hem om middagen; ty de hade fått höra att de skulle äta där.
När sedan Josef hade kommit hem, förde de skänkerna, som de hade med sig, in till honom i huset och föllo ned för honom till jorden.
Och han hälsade dem och frågade: »Står det väl till med eder fader, den gamle, som I taladen om?
Lever han ännu?»
De svarade: »Ja, det står väl till med vår fader, din tjänare; han lever ännu.»
Och de bugade sig och föllo ned för honom.
Och när han lyfte upp sina ögon och fick se sin broder Benjamin, sin moders son, frågade han: »Är detta eder yngste broder, den som I taladen om med mig?»
Därpå sade han: »Gud vare dig nådig, min son.»
Men Josef bröt av sitt tal, ty hans hjärta upprördes av kärlek till brodern, och han sökte tillfälle att gråta ut och gick in i sin kammare och grät där.
Därefter, sedan han hade tvagit sitt ansikte, gick han åter ut och betvang sig och sade: »Sätten fram mat.»
Och de satte fram särskilt för honom och särskilt för dem och särskilt för de egyptier som åto tillsammans med honom; ty egyptierna få icke äta tillsammans med hebréerna; sådant är nämligen en styggelse för egyptierna.
Och de fingo sina platser mitt emot honom, den förstfödde främst såsom den förstfödde, sedan de yngre, var och en efter sin ålder; och männen sågo med förundran på varandra.
Och han lät bära till dem av rätterna på sitt bord, och Benjamin fick fem gånger så mycket som var och en av de andra.
Och de drucko sig glada med honom.
Därefter bjöd han sin hovmästare och sade: »Fyll männens säckar med säd, så mycket de kunna rymma, och lägg vars och ens penningar överst i hans säck.
Och min bägare, silverbägaren, skall du lägga överst i den yngstes säck, tillika med penningarna för hans säd.»
Och han gjorde såsom Josef hade sagt.
Om morgonen, då det blev dager, fingo männen fara med sina åsnor.
Men när de hade kommit ett litet stycke utom staden, sade Josef till sin hovmästare: »Stå upp och sätt efter männen; och när du hinner upp dem, så säg till dem: 'Varför haven I lönat gott med ont?
Det är ju just den bägaren som min herre dricker ur, och som han plägar spå med.
Det är en ond gärning I haven gjort.'»
När han nu hann upp dem, sade han detta till dem.
Då svarade de honom: »Varför talar min herre så?
Bort det, att dina tjänare skulle göra sådant!
De penningar som vi funno överst i våra säckar hava vi ju fört tillbaka till dig från Kanaans land.
Huru skulle vi då kunna vilja stjäla silver eller guld ur din herres hus?
Den bland dina tjänare, som den finnes hos, han må dö; därtill vilja vi andra bliva min herres trälar.»
Han svarade: »Ja, vare det såsom I haven sagt; den som den finnes hos, han skall bliva min träl.
Men I andra skolen vara utan skuld.»
Och de skyndade sig att lyfta ned var och en sin säck på jorden, och öppnade var och en sin säck.
Och han begynte att söka hos den äldste och slutade hos den yngste; och bägaren fanns i Benjamins säck.
Då revo de sönder sina kläder och lastade åter var och en sin åsna och vände tillbaka till staden.
Och Juda och hans bröder gingo in i Josefs hus, där denne ännu var kvar; och de föllo ned till jorden för honom.
Då sade Josef till dem: »Vad haven I gjort!
Förstoden I icke att en man sådan som jag kan spå?»
Juda svarade: Vad skola vi säga till min herre, vad skola vi tala, och huru skola vi rättfärdiga oss?
Gud har funnit dina tjänares missgärning.
Se, vi äro min herres trälar, vi andra såväl som den som bägaren har blivit funnen hos.»
Men han sade: »Bort det, att jag skulle så göra!
Den som bägaren har blivit funnen hos, han skall bliva min träl.
Men I andra mån i frid fara hem till eder fader.»
Då trädde Juda fram till honom och sade: »Hör mig, herre; låt din tjänare tala ett ord inför min herre, och må din vrede icke upptändas mot din tjänare; ty du är såsom Farao.
Min herre frågade sina tjänare och sade: 'Haven I eder fader eller någon broder ännu därhemma?'
Och vi svarade min herre: 'Vi hava en åldrig fader och en son till honom, en som är född på hans ålderdom och ännu är ung; men en broder till denne är död, så att han allena är kvar efter sin moder, och hans fader har honom kär.'
Då sade du till dina tjänare: 'Fören honom hitned till mig, så att jag kan låta mitt öga vila på honom.'
Och vi svarade min herre: 'Ynglingen kan icke lämna sin fader, ty om han lämnade sin fader, så skulle denne dö.'
Men du sade till dina tjänare: 'Om eder yngste broder icke följer med eder hitned, så fån I icke mer komma inför mitt ansikte.'
När vi därefter hade kommit hem till din tjänare, min fader, berättade vi för honom vad min herre hade sagt.
Och när sedan vår fader sade: 'Faren tillbaka och köpen litet säd till föda åt oss',
svarade vi: 'Vi kunna icke fara ditned; allenast på det villkoret vilja vi fara, att vår yngste broder följer med oss; ty vi få icke komma inför mannens ansikte om vår yngste broder icke är med oss.
Men din tjänare, min fader, sade till oss: 'I veten själva att min hustru har fött åt mig två söner,
och den ene gick bort ifrån mig, och jag sade: förvisso är han ihjälriven.
Och jag har icke sett honom sedan den tiden.
Om I nu tagen också denne ifrån mig och någon olycka händer honom, så skolen I bringa mina grå hår med jämmer ned i dödsriket.'
Om jag alltså kommer hem till din tjänare, min fader, utan att vi hava med oss ynglingen, som vår faders hjärta är så fäst vid,
då bliver det hans död, när han ser att ynglingen icke är med; och dina tjänare skulle så bringa din tjänares, vår faders, grå hår med sorg ned i dödsriket.
Ty jag, din tjänare, har lovat min fader att ansvara för ynglingen och har sagt, att om jag icke för denne till honom igen, så vill jag vara en syndare inför min fader i all min tid.
Låt nu därför din tjänare stanna kvar hos min herre såsom träl, i ynglingens ställe, men låt ynglingen fara hem med sina bröder.
Ty huru skulle jag kunna fara hem till min fader utan att hava ynglingen med mig?
Jag förmår icke se den jämmer som då skulle komma över min fader.»
Då kunde Josef icke längre betvinga sig inför alla dem som stodo omkring honom.
Han ropade: »Må alla gå ut härifrån.»
Och ingen fick stanna inne hos Josef, när han gav sig till känna för sina bröder.
Och han brast ut i högljudd gråt, så att egyptierna hörde det; också Faraos husfolk hörde det.
Och Josef sade till sina bröder: »Jag är Josef.
Lever min fader ännu?»
Men hans bröder kunde icke svara honom, så förskräckta blevo de för honom.
Då sade Josef till sina bröder: »Kommen hitfram till mig.»
Och när de kommo fram, sade han: »Jag är Josef, eder broder, som I sålden till Egypten.
Men varen nu icke bedrövade och grämen eder icke däröver att I haven sålt mig hit: ty för att bevara människors liv har Gud sänt mig hit före eder.
I två år har nu hungersnöd varit i landet, och ännu återstå fem år under vilka man varken skall plöja eller skörda.
Men Gud sände mig hit före eder, för att I skullen bliva kvar på jorden och behållas vid liv, ja, till räddning för många.
Så haven nu icke I sänt mig hit, utan Gud; och han har gjort mig till Faraos högste rådgivare och till en herre över hela hans hus och till en furste över hela Egyptens land.
Skynden eder nu och faren hem till min fader, och sägen till honom: 'Så säger din son Josef: Gud har satt mig till en herre över hela Egypten; kom ned till mig, dröj icke.
Du skall få bo i landet Gosen och vara mig nära, du med dina barn och barnbarn, dina får och fäkreatur och allt vad som tillhör dig.
Jag vill där försörja dig -- ty ännu återstå fem hungerår -- så att varken du eller ditt hus eller någon som hör dig till skall lida nöd.
I sen ju med egna ögon, också min broder Benjamin ser med egna ögon, att det är jag, som med egen mun talar till eder.
Berätten nu för min fader om all min härlighet i Egypten och om allt vad I haven sett, och skynden eder att föra min fader hitned.»
Så föll han sin broder Benjamin om halsen och grät, och Benjamin grät vid hans hals.
Och han kysste alla sina bröder och grät i deras armar.
Sedan samtalade hans bröder med honom.
När nu det ryktet spordes i Faraos hus, att Josefs bröder hade kommit, behagade detta Farao och hans tjänare väl.
Och Farao sade till Josef: »Säg till dina bröder: 'Detta skolen I göra: lasten edra djur och faren hem till Kanaans land;
hämten så eder fader och edert folk och kommen hit till mig, så skall jag giva eder det bästa som finnes i Egyptens land, och I skolen få äta av landets fetma.'
Alltså bjuder jag dig nu att säga: 'Detta skolen I göra: tagen eder vagnar i Egyptens land för edra späda barn och edra hustrur, och hämten eder fader och kommen hit.
Och bekymren eder icke om edert bohag; ty det bästa som finnes i hela Egyptens land skall höra eder till.'»
Israels söner gjorde så, och Josef gav dem vagnar, efter Faraos befallning, och gav dem kost för resan.
Och han gav åt dem alla var sin högtidsdräkt, men åt Benjamin gav han tre hundra siklar silver och fem högtidsdräkter.
Och till sin fader sände han likaledes gåvor: tio åsnor, lastade med det bästa Egypten hade, och tio åsninnor, lastade med säd och bröd och andra livsmedel åt hans fader för resan.
Därefter lät han sina bröder fara, och de begåvo sig åstad; och han sade till dem: »Kiven icke på vägen.»
Så foro de upp från Egypten och kommo till sin fader Jakob i Kanaans land;
och de berättade för honom och sade: »Josef lever ännu, och han är en furste över hela Egyptens land.»
Då greps hans hjärta av vanmakt, ty han kunde icke tro dem.
Men när de omtalade för honom allt vad Josef hade sagt till dem, och när han såg vagnarna som Josef hade sänt för att hämta honom, då fick deras fader Jakobs ande åter liv.
Och Israel sade: »Det är nog; min son Josef lever ännu.
Jag vill fara och se honom, förrän jag dör.»
Och Israel bröt upp med allt vad honom tillhörde.
Och när han kom till Beer-Seba, offrade han slaktoffer åt sin fader Isaks Gud.
Och Gud talade till Israel i en syn om natten; han sade: »Jakob!
Jakob!»
Han svarade: »Här är jag.»
Då sade han: »Jag är Gud, din faders Gud; frukta icke för att draga ned till Egypten, ty där skall jag göra dig till ett stort folk.
Jag skall själv draga ned med dig till Egypten, jag skall ock föra dig åter upp därifrån; och Josefs hand skall tillsluta dina ögon.»
Och Jakob bröt upp från Beer-Seba; och Israels söner satte sin fader Jakob och sina späda barn och sina hustrur på vagnarna som Farao hade sänt för att hämta honom.
Och de togo sin boskap och de ägodelar som de hade förvärvat i Kanaans land och kommo så till Egypten, Jakob och alla hans avkomlingar med honom.
Sina söner och sonsöner, sina döttrar och sondöttrar, alla sina avkomlingar, förde han med sig till Egypten.
Dessa äro namnen på Israels barn som kommo till Egypten: Jakob och hans söner.
Jakobs förstfödde var Ruben,
och Rubens söner voro Hanok, Pallu, Hesron och Karmi.
Simeons söner voro Jemuel, Jamin, Ohad, Jakin, Sohar och Saul, den kananeiska kvinnans son.
Levis söner voro Gerson, Kehat och Merari.
Judas söner voro Er, Onan, Sela, Peres och Sera -- men Er och Onan dogo i Kanaans land -- och Peres' söner voro Hesron och Hamul.
Isaskars söner voro Tola, Puva, Job och Simron.
Sebulons söner voro Sered, Elon och Jaleel.
Dessa voro Leas söner, de som hon födde åt Jakob i Paddan-Aram; tillika födde hon åt honom dottern Dina.
Söner och döttrar utgjorde tillsammans trettiotre personer.
Gads söner voro Sifjon och Haggi, Suni och Esbon, Eri och Arodi och Areli.
Asers söner voro Jimna, Jisva, Jisvi och Beria; och deras syster var Sera; men Berias söner voro Heber och Malkiel.
Dessa voro söner till Silpa, som Laban hade givit åt sin dotter Lea, och dessa födde hon åt Jakob, sexton personer.
Rakels, Jakobs hustrus, söner voro Josef och Benjamin.
Och de söner som föddes åt Josef i Egyptens land voro Manasse och Efraim; de föddes åt honom av Asenat, dotter till Poti-Fera, prästen i On.
Och Benjamins söner voro Bela, Beker och Asbel, Gera och Naaman, Ehi och Ros, Muppim och Huppim och Ard.
Dessa voro Rakels söner, de som föddes åt Jakob, tillsammans fjorton personer.
Dans söner voro Husim.
Naftalis söner voro Jaseel, Guni, Jeser och Sillem.
Dessa voro söner till Bilha, som Laban hade givit åt sin dotter Rakel, och dessa födde hon åt Jakob, tillsammans sju personer.
De som kommo med Jakob till Egypten, de som hade utgått från hans länd, utgjorde alla tillsammans sextiosex personer, förutom Jakobs sonhustrur.
Och Josefs söner, vilka föddes åt honom i Egypten, voro två.
De personer av Jakobs hus, som kommo till Egypten, utgjorde tillsammans sjuttio.
Och han sände Juda framför sig till Josef, för att denne skulle visa honom vägen till Gosen.
Så kommo de till landet Gosen.
Och Josef lät spänna för sin vagn och for upp till Gosen för att möta sin fader Israel.
Och när han kom fram till honom, föll han honom om halsen och grät länge vid hans hals.
Och Israel sade till Josef: »Nu vill jag gärna dö, sedan jag har sett ditt ansikte och sett att du ännu lever.»
Därefter sade Josef till sina bröder och sin faders folk: »Jag vill fara upp och berätta för Farao och säga till honom: 'Mina bröder och min faders folk, som hittills hava bott i Kanaans land, hava kommit till mig.
Och dessa män äro fårherdar, ty de hava idkat boskapsskötsel; och sina får och fäkreatur och allt vad de äga hava de fört med sig.'
När sedan Farao kallar eder till sig och frågar: 'Vad är edert yrke?',
skolen I svara: 'Vi, dina tjänare, hava idkat boskapsskötsel från vår ungdom ända till nu, vi såväl som våra fäder.'
Så skolen I få bo i landet Gosen; ty alla fårherdar äro en styggelse för egyptierna.»
Och Josef kom och berättade för Farao och sade: »Min fader och mina bröder hava kommit från Kanaans land med sina får och fäkreatur och allt vad de äga; och de äro nu i landet Gosen.»
Och han hade bland sina bröder tagit ut fem män; dem ställde han fram inför Farao.
Då frågade Farao hans bröder: »Vad är edert yrke?»
De svarade Farao: »Dina tjänare äro fårherdar, såsom ock våra fäder hava varit.»
Och de sade ytterligare till Farao: »Vi hava kommit för att bo någon tid här i landet; ty dina tjänare hade intet bete för sina får, eftersom hungersnöden är så svår i Kanaans land.
Så låt nu dina tjänare bo i landet Gosen.»
Då sade Farao till Josef: »Din fader och dina bröder hava alltså nu kommit till dig.
Egyptens land ligger öppet för dig; i den bästa delen av landet må du låta din fader och dina bröder bo.
Må de bo i landet Gosen, och ifall du vet om några bland dem att de äro dugande män, så sätt dessa till uppsyningsmän över min boskap.»
Sedan hämtade Josef sin fader Jakob och förde honom fram inför Farao, och Jakob hälsade Farao.
Men Farao frågade Jakob: »Huru hög är din ålder?»
Jakob svarade Farao: »Min vandringstid har varat ett hundra trettio år.
Få och onda hava mina levnadsår varit, de nå icke upp till antalet av mina fäders levnadsår under deras vandringstid.»
Och Jakob tog avsked av Farao och gick ut ifrån honom.
Men Josef lät sin fader och sina bröder bo i Egyptens land och gav dem besittning där, i den bästa delen av landet, i landet Rameses, såsom Farao hade bjudit.
Och Josef försörjde sin fader och sina bröder och hela sin faders hus, och gav var och en underhåll efter antalet av hans barn.
Men ingenstädes i landet fanns bröd, ty hungersnöden var mycket svår, så att Egyptens land och Kanaans land försmäktade av hunger.
Och för den säd som folket köpte samlade Josef till sig alla penningar som funnos i Egyptens land och i Kanaans land; och Josef lät föra penningarna in i Faraos hus.
Men när penningarna togo slut i Egyptens land och i Kanaans land, kommo alla egyptier till Josef och sade: »Giv oss bröd; icke vill du väl att vi skola dö i din åsyn?
Vi hava ju inga penningar mer.»
Josef svarade: »Fören hit eder boskap, så skall jag giva eder bröd i utbyte mot eder boskap, om I icke mer haven några penningar.»
Då förde de sin boskap till Josef, och Josef gav dem bröd i utbyte mot deras hästar, får, fäkreatur och åsnor.
Så underhöll han dem det året och gav dem bröd i utbyte mot all deras boskap.
Så gick detta år till ända.
Men det följande året kommo de åter till honom och sade till honom: »Vi vilja icke dölja det för min herre: penningarna äro slut, och den boskap vi ägde har kommit i min herres ägo; intet annat finnes nu kvar att giva åt min herre än våra kroppar och vår jord.
Icke vill du att vi skola förgås inför dina ögon, vi med vår åkerjord?
Köp oss och vår jord för bröd, så vilja vi med vår jord bliva Faraos trälar; giv oss allenast utsäde, för att vi må leva och icke dö, och för att jorden icke må läggas öde.»
Då köpte Josef all jord i Egypten åt Farao; ty egyptierna sålde var och en sin åker, eftersom hungersnöden så svårt tryckte dem.
Så blev jorden Faraos egendom.
Och folket förflyttade han till städerna, från den ena ändan av Egyptens område till den andra.
Allenast prästernas jord köpte han icke, ty prästerna hade sitt bestämda underhåll av Farao, och de levde av det bestämda underhåll som Farao gav dem; därför behövde de icke sälja sin jord.
Och Josef sade till folket: »Se, jag har nu köpt eder och eder jord åt Farao.
Där haven I utsäde; besån nu jorden.
Och när grödan kommer in, skolen I giva en femtedel åt Farao; men fyra femtedelar skolen I själva hava till utsäde på åkern och till föda för eder och dem som I haven i edra hus och till föda för edra barn.»
De svarade: »Du har behållit oss vid liv; låt oss finna nåd för min herres ögon, så vilja vi vara Faraos trälar.»
Så gjorde Josef det till en stadga, som ännu i dag gäller för Egyptens jord, att man skulle giva femtedelen åt Farao.
Allenast prästernas jord blev icke Faraos egendom.
Så bodde nu Israel i Egyptens land, i landet Gosen; och de fingo sina besittningar där och voro fruktsamma och förökade sig storligen.
Och Jakob levde sjutton år i Egyptens land, så att hans levnadsålder blev ett hundra fyrtiosju år.
Då nu tiden närmade sig att Israel skulle dö, kallade han till sig sin son Josef och sade till honom: »Om jag har funnit nåd för dina ögon, så lägg din hand under min länd och lova att visa mig din kärlek och trofasthet därmed att du icke begraver mig i Egypten;
fastmer, när jag har gått till vila hos mina fäder, skall du föra mig från Egypten och begrava mig i deras grav.»
Han svarade: »Jag skall göra såsom du har sagt.»
Men han sade: »Giv mig din ed därpå.»
Och han gav honom sin ed.
Då tillbad Israel, böjd mot sängens huvudgärd.
En tid härefter blev det sagt till Josef: »Din fader är nu sjuk.»
Då tog han med sig sina båda söner, Manasse och Efraim.
Och man berättade för Jakob och sade: »Din son Josef har nu kommit till dig.»
Då tog Israel styrka till sig och satte sig upp i sängen.
Och Jakob sade till Josef: »Gud den Allsmäktige uppenbarade sig för mig i Lus i Kanaans land och välsignade mig
och sade till mig: 'Se, jag skall göra dig fruktsam och föröka dig och låta skaror av folk komma av dig, och skall giva åt din säd efter dig detta land till evärdlig besittning.'
Dina båda söner, som äro födda åt dig i Egyptens land, innan jag kom hit till dig i Egypten, de skola nu vara mina: Efraim och Manasse skola vara mina, likasom Ruben och Simeon.
Men de barn som du har fött efter dem skola vara dina; de skola bära sina bröders namn i dessas arvedel.
Se, när jag kom från Paddan, dog Rakel ifrån mig i Kanaans land, under resan, då det ännu var ett stycke väg fram till Efrat; och jag begrov henne där vid vägen till Efrat.»
Stället heter nu Bet-Lehem.
Då nu Israel fick se Josefs söner, sade han: »Vilka äro dessa?»
Josef svarade sin fader: »Det är mina söner, som Gud har givit mig här.»
Då sade han: »För dem hit till mig, på det att jag må välsigna dem.»
Och Israels ögon voro skumma av ålder, så att han icke kunde se.
Så förde han dem då fram till honom, och han kysste dem och tog dem i famn.
Och Israel sade till Josef: »Jag hade icke tänkt att jag skulle få se ditt ansikte, men nu har Gud låtit mig se till och med avkomlingar av dig.»
Och Josef förde dem bort ifrån hans knän och föll ned till jorden på sitt ansikte.
Sedan tog Josef dem båda vid handen, Efraim i sin högra hand, till vänster framför Israel, och Manasse i sin vänstra hand, till höger framför Israel, och förde dem så fram till honom.
Men Israel räckte ut sin högra hand och lade den på Efraims huvud, fastän han var den yngre, och sin vänstra hand på Manasses huvud; han lade alltså sina händer korsvis, ty Manasse var den förstfödde.
Och han välsignade Josef och sade: »Den Gud inför vilken mina fäder, Abraham och Isak, hava vandrat, den Gud som har varit min herde från min födelse ända till denna dag,
den ängel som har förlossat mig från allt ont, han välsigne dessa barn; och må de uppkallas efter mitt och mina fäders, Abrahams och Isaks, namn, och må de föröka sig och bliva talrika på jorden.»
Men när Josef såg att hans fader lade sin högra hand på Efraims huvud, misshagade detta honom, och han fattade sin faders hand och ville flytta den från Efraims huvud på Manasses huvud.
Och Josef sade till sin fader: »Icke så, min fader; denne är den förstfödde, lägg din högra hand på hans huvud.»
Men hans fader ville icke; han sade: »Jag vet det, min son, jag vet det; också av honom skall ett folk komma, också han skall bliva stor; men hans yngre broder skall dock bliva större än han, och hans avkomma skall bliva ett talrikt folk.»
Så välsignade han dem på den dagen och sade: »Med ditt namn skall Israel välsigna, så att man skall säga: Gud göre dig lik Efraim och Manasse.»
Så satte han Efraim framför Manasse.
Och Israel sade till Josef: »Se, jag dör; men Gud skall vara med eder och föra eder tillbaka till edra fäders land.
Och utöver vad jag giver dina bröder giver jag dig en särskild höjdsträcka som jag med mitt svärd och min båge har tagit från amoréerna.»
Och Jakob kallade sina söner till sig och sade: Församlen eder, på det att jag må förkunna eder vad som skall hända eder i kommande dagar:
Kommen tillhopa och hören, I Jakobs söner; hören på eder fader Israel.
Ruben, min förstfödde är du, min kraft och min styrkas förstling, främst i myndighet och främst i makt.
Du sjuder över såsom vatten, du skall icke bliva den främste, ty du besteg din faders läger; då gjorde du vad skändligt var.
Ja, min bädd besteg han!
Simeon och Levi äro bröder; deras vapen äro våldets verktyg.
Min själ inlåte sig ej i deras råd, min ära tage ingen del i deras samkväm; ty i sin vrede dräpte de män, och i sitt överdåd stympade de oxar.
Förbannad vare deras vrede, som är så våldsam, och deras grymhet, som är så hård!
Jag skall förströ dem i Jakob, jag skall förskingra dem i Israel.
Dig, Juda, dig skola dina bröder prisa ; din hand skall vara på dina fienders nacke, för dig skola din faders söner buga sig.
Ett ungt lejon är Juda; från rivet byte har du dragit ditupp, min son.
Han har lagt sig ned, han vilar såsom ett lejon, såsom en lejoninna -- vem vågar oroa honom?
Spiran skall icke vika ifrån Juda, icke härskarstaven ifrån hans fötter, till dess han kommer till Silo och folken bliva honom hörsamma.
Han binder vid vinträdet sin åsna, vid ädla rankan sin åsninnas fåle.
Han tvår sina kläder i vin, sin mantel i druvors blod.
Hans ögon äro dunkla av vin och hans tänder vita av mjölk.
Sebulon skall bo vid havets strand, vid stranden, där skeppen ligga; sin sida skall han vända mot Sidon.
Isaskar är en stark åsna, som ligger i ro i sin inhägnad.
Och han såg att viloplatsen var god, och att landet var ljuvligt; då böjde han sin rygg under bördor och blev en arbetspliktig tjänare.
Dan skall skaffa rätt åt sitt folk, han såväl som någon av Israels stammar.
Dan skall vara en orm på vägen, en huggorm på stigen, en som biter hästen i foten, så att ryttaren faller baklänges av.
HERRE, jag bidar efter din frälsning!
Gad skall trängas av skaror , men själv skall han tränga dem på hälarna.
Från Aser kommer fetma, honom till mat; konungsliga läckerheter har han att giva.
Naftali är en snabb hind; han har sköna ord att giva.
Ett ungt fruktträd är Josef, ett ungt fruktträd vid källan; dess grenar nå upp över muren.
Bågskyttar oroa honom, de skjuta på honom och ansätta honom;
dock förbliver hans båge fast, och hans händer och armar spänstiga, genom dens händer, som är den Starke i Jakob, genom honom som är herden, Israels klippa,
genom din faders Gud -- han skall hjälpa dig. genom den Allsmäktige -- han skall välsigna dig med välsignelser från himmelen därovan, välsignelser från djupet som utbreder sig därnere, välsignelser från bröst och sköte.
Din faders välsignelser nå högt, högre än mina förfäders välsignelser, de nå upp till de eviga höjdernas härlighet.
De skola komma över Josefs huvud, över dens hjässa, som är en furste bland sina bröder.
Benjamin är en glupande ulv; om morgonen förtär han rov, och om aftonen utskiftar han byte.»
Alla dessa äro Israels stammar, tolv till antalet, och detta är vad deras fader talade till dem, när han välsignade dem; åt var och en av dem gav han sin särskilda välsignelse.
Och han bjöd dem och sade till dem: »Jag skall nu samlas till mitt folk; begraven mig bredvid mina fäder, i grottan på hetiten Efrons åker,
i den grotta som ligger på åkern i Makpela, gent emot Mamre, i Kanaans land, den åker som Abraham köpte till egen grav av hetiten Efron,
där de hava begravit Abraham och hans hustru Sara, där de ock hava begravit Isak och hans hustru Rebecka, och där jag själv har begravit Lea,
på den åkern som jämte grottan där köptes av Hets barn.»
När Jakob hade givit sina söner denna befallning, drog han sina fötter upp i sängen; och han gav upp andan och blev samlad till sina fäder.
Då föll Josef ned över sin faders ansikte och grät över honom och kysste honom.
Och Josef bjöd läkarna som han hade i sin tjänst att de skulle balsamera hans fader; och läkarna balsamerade Israel.
Därtill åtgingo fyrtio dagar; så många dagar åtgå nämligen för balsamering.
Och egyptierna begräto honom i sjuttio dagar.
Men när gråtodagarna efter honom voro förbi, talade Josef till Faraos husfolk och sade: »Om jag har funnit nåd för edra ögon, så framfören till Farao dessa mina ord:
Min fader har tagit en ed av mig och sagt: 'När jag är död, begrav mig då i den grav som jag har låtit gräva åt mig i Kanaans land.'
Så låt mig nu fara ditupp och begrava min fader; sedan skall jag komma tillbaka igen.»
Farao svarade: »Far ditupp och begrav din fader, efter den ed som han har tagit av dig.»
Då for Josef upp för att begrava sin fader, och med honom foro alla Faraos tjänare, de äldste i hans hus och alla de äldste i Egyptens land,
därtill allt Josefs husfolk och hans bröder och hans faders husfolk; allenast sina kvinnor och barn, och sina får och fäkreatur lämnade de kvar i landet Gosen.
Och med honom foro ditupp både vagnar och ryttare; och det var en mycket stor skara.
När de nu kommo till Goren-Haatad, på andra sidan Jordan, höllo de där en mycket stor och högtidlig dödsklagan, och han anställde en sorgefest efter sin fader i sju dagar.
Och när landets inbyggare, kananéerna, sågo sorgefesten i Goren-Haatad, sade de: »Det är en högtidlig sorgefest som egyptierna här hålla.»
Därav fick stället namnet Abel-Misraim; det ligger på andra sidan Jordan.
Och hans söner gjorde med honom såsom han hade bjudit dem:
hans söner förde honom till Kanaans land och begrovo honom i grottan på åkern i Makpela, den åker som Abraham hade köpt till egen grav av hetiten Efron, gent emot Mamre.
Och sedan Josef hade begravit sin fader, vände han tillbaka till Egypten med sina bröder och alla dem som hade farit upp med honom för att begrava hans fader.
Men när Josefs bröder sågo att deras fader var död, tänkte de: »Kanhända skall Josef nu bliva hätsk mot oss och vedergälla oss allt det onda som vi hava gjort mot honom.»
Därför sände de bud till Josef och läto säga: »Din fader bjöd oss så före sin död:
'Så skolen I säga till Josef: Käre, förlåt dina bröder vad de hava brutit och syndat, i det att de hava handlat så illa mot dig.'
Förlåt alltså nu din faders Guds tjänare vad de hava brutit.»
Och Josef grät, när de läto säga detta till honom.
Sedan kommo ock hans bröder själva och föllo ned för honom och sade: »Se, vi vilja vara tjänare åt dig.»
Men Josef sade till dem: »Frukten icke.
Hållen I då mig för Gud?
I tänkten ont mot mig, men Gud har tänkt det till godo, för att låta det ske, som nu har skett, och så behålla mycket folk vid liv.
Frukten därför nu icke; jag skall försörja eder och edra kvinnor och barn.»
Och han tröstade dem och talade vänligt med dem.
Och Josef bodde kvar i Egypten med sin faders hus; och Josef blev ett hundra tio år gammal.
Och Josef fick se Efraims barn till tredje led; också av Makir, Manasses son, föddes barn i Josefs sköte.
Och Josef sade till sina bröder: »Jag dör, men Gud skall förvisso se till eder, och föra eder upp från detta land till det land som han med ed har lovat åt Abraham, Isak och Jakob.»
Och Josef tog en ed av Israels barn och sade: »När nu Gud ser till eder, fören då mina ben härifrån.»
Och Josef dog, när han var ett hundra tio år gammal.
Och man balsamerade honom, och han lades i en kista, i Egypten.
Och dessa äro namnen på Israels söner, som kommo till Egypten; med Jakob kommo de, var och en med sitt hus:
Ruben, Simeon, Levi och Juda,
Isaskar, Sebulon och Benjamin,
Dan och Naftali, Gad och Aser.
Tillsammans utgjorde de som hade utgått från Jakobs länd sjuttio personer; men Josef var redan förut i Egypten.
Och Josef dog och alla hans bröder och hela det släktet.
Men Israels barn voro fruktsamma och växte till och förökade sig och blevo övermåttan talrika, så att landet blev uppfyllt av dem.
Då uppstod en ny konung över Egypten, en som icke visste av Josef.
Och denne sade till sitt folk: »Se, Israels barns folk är oss för stort och mäktigt.
Välan, låt oss då gå klokt till väga med dem; eljest kunde de ännu mer föröka sig; och om ett krig komme på, kunde de förena sig med våra fiender och begynna krig mot oss och sedan draga bort ur landet.»
Alltså satte man arbetsfogdar över dem och förtryckte dem med trälarbeten.
Och de måste bygga åt Farao förrådsstäder, Pitom och Raamses.
Men ju mer man förtryckte dem, dess mer förökade de sig, och dess mer utbredde de sig, så att man begynte gruva sig för Israels barn.
Därför pålade egyptierna Israels barn ytterligare tvångsarbeten
och förbittrade deras liv med hårt arbete på murbruk och tegel och med alla slags arbeten på marken korteligen, med tvångsarbeten av alla slag, som de läto dem utföra
Och konungen i Egypten talade till de hebreiska kvinnor -- den ena hette Sifra, den andra Pua -- som hjälpte barnaföderskorna,
han sade: »När I förlösen de hebreiska kvinnorna, så sen efter, då de föda: om det är ett gossebarn, så döden det; är det ett flickebarn, så må det leva.»
Men hjälpkvinnorna fruktade Gud och gjorde icke såsom konungen i Egypten hade sagt till dem, utan läto barnen leva.
Då kallade konungen i Egypten hjälpkvinnorna till sig och sade till dem: »Varför gören I så och låten barnen leva?»
Hjälpkvinnorna svarade Farao: »De hebreiska kvinnorna äro icke såsom de egyptiska.
De äro kraftigare; förrän hjälpkvinnan kommer till dem, hava de fött.»
Och Gud lät det gå väl för hjälpkvinnorna; och folket förökade sig och blev mycket talrikt.
Eftersom hjälpkvinnorna fruktade Gud, lät han deras hus förkovras.
Då bjöd Farao allt sitt folk och sade: »Alla nyfödda gossebarn- skolen I kasta i Nilfloden, men all flickebarn mån I låta leva.»
Och en man av Levis hus gick åstad och tog till hustru Levis dotter.
Och hustrun blev havande och födde en son.
Och hon såg att det var ett vackert barn och dolde honom i tre månader.
Men när hon icke längre kunde dölja honom, tog hon en kista av rör, beströk den med jordbeck och tjära och lade barnet däri och satte den så i vassen vid stranden av Nilfloden.
Och hans syster ställde sig ett stycke därifrån, för att se huru det skulle gå med honom.
Och Faraos dotter kom ned till floden för att bada, och hennes tärnor gingo utmed floden.
När hon nu fick se kistan i vassen, sände hon sin tjänarinna dit och lät hämta den till sig.
Och när hon öppnade den, fick hon se barnet och såg att det var en gosse, och han grät.
Då ömkade hon sig över honom och sade: »Detta är ett av de hebreiska barnen.»
Men hans syster frågade Faraos dotter: »Vill du att jag skall gå och kalla hit till dig en hebreisk amma som kan amma upp barnet åt dig?»
Faraos dotter svarade henne: »Ja, gå.»
Då gick flickan och kallade dit barnets moder.
Och Faraos dotter sade till henne: »Tag detta barn med dig, och amma upp det åt mig, så vill jag giva dig lön därför.»
Och kvinnan tog barnet och ammade upp det.
När sedan gossen hade vuxit upp; förde hon honom till Faraos dotter, och denna upptog honom såsom sin son och gav honom namnet Mose , »ty», sade hon, »ur vattnet har jag dragit upp honom».
På den tiden hände sig att Mose, sedan han hade blivit stor, gick ut till sina bröder och såg på deras trälarbete.
Och han fick se att en egyptisk man slog en hebreisk man, en av hans bröder.
då vände han sig åt alla sidor, och när han såg att ingen annan människa fanns där, slog han ihjäl egyptiern och gömde honom i sanden.
Dagen därefter gick han åter ut och fick då se två hebreiska män träta med varandra.
Då sade han till den som gjorde orätt: »Skall du slå din landsman?»
Han svarade: »Vem har satt dig till hövding och domare över oss?
Vill du dräpa mig, såsom du dräpte egyptiern?»
Då blev Mose förskräckt och tänkte: »Så har då saken blivit känd.»
Också fick Farao höra om denna sak och ville dräpa Mose.
Men Mose flydde bort undan Farao; och han stannade i Midjans land; där satte han sig vid en brunn.
Och prästen i Midjan hade sju döttrar.
Dessa kommo nu för att hämta upp vatten och skulle fylla hoarna för att vattna sin faders får.
Då kommo herdarna och ville driva bort dem; men Mose stod upp och hjälpte dem och vattnade deras får.
När de sedan kommo hem till sin fader Reguel, sade han: »Varför kommen I så snart hem i dag?»
De svarade: »En egyptisk man hjälpte oss mot herdarna; därtill hämtade han upp vatten åt oss och vattnade fåren.»
Då sade han till sina döttrar: »Var är han då?
Varför läten I mannen bliva kvar där?
Inbjuden honom att komma och äta med oss».
Och Mose beslöt sig för att stanna hos mannen, och denne gav åt Mose sin dotter Sippora till hustru.
Hon födde en son, och han gav honom namnet Gersom, »ty», sade han, »jag är en främling i ett land som icke är mitt».
Så förflöt en lång tid, och därunder dog konungen i Egypten.
Men Israels barn suckade över sin träldom och klagade; och deras rop över träldomen steg upp till Gud.
Och Gud hörde deras jämmer, och Gud tänkte på sitt förbund med Abraham, Isak och Jakob.
Och Gud såg till Israels barn, och Gud lät sig vårda om dem.
Och Mose vaktade fåren åt sin svärfader Jetro, prästen i Midjan.
Och han drev en gång fåren bortom öknen och kom så till Guds berg Horeb.
Där uppenbarade sig HERRENS ängel för honom i en eldslåga som slog upp ur en buske.
Han såg att busken brann av elden, och att busken dock icke blev förtärd.
Då tänkte Mose: »Jag vill gå ditbort och betrakta den underbara synen och se varför busken icke brinner upp.»
När då HERREN såg att han gick åstad för att se, ropade Gud till honom ur busken och sade: »Mose!
Mose!»
Han svarade: »Här är jag.»
Då sade han: »Träd icke hit; drag dina skor av dina fötter, ty platsen där du står är helig mark.»
Och han sade ytterligare: »Jag är din faders Gud, Abrahams Gud, Isaks Gud och Jakobs Gud.»
Då skylde Mose sitt ansikte, ty han fruktade för att se på Gud.
Och HERREN sade: »Jag har nogsamt sett mitt folks betryck i Egypten, och jag har hört huru de ropa över sina plågare; jag vet vad de måste lida.
Därför har jag stigit ned för att rädda dem ur egyptiernas våld och föra dem från det landet upp till ett gott och rymligt land, ett land som flyter av mjölk och honung, det land där kananéer, hetiter, amoréer, perisséer, hivéer och jebuséer bo.
Fördenskull, eftersom Israels barns rop har kommit till mig, och jag därjämte har sett huru egyptierna förtrycka dem,
därför må du nu gå åstad, jag vill sända dig till Farao; och du skall föra mitt folk, Israels barn, ut ur Egypten»
Men Mose sade till Gud: »Vem är jag, att jag skulle gå till Farao, och att jag skulle föra Israels barn ut ur Egypten?»
Han svarade: »Jag vill vara med dig.
Och detta skall för dig vara tecknet på att det är jag som har sänt dig: när du har fört folket ut ur Egypten, skolen I hålla gudstjänst på detta berg.»
Då sade Mose till Gud: »När jag nu kommer till Israels barn och säger till dem: 'Edra fäders Gud har sänt mig till eder', och de fråga mig; 'Vad är hans namn?', vad skall jag då svara dem?»
Gud sade till Mose: »Jag är den jag är.»
Och han sade vidare: »Så skall du säga till Israels barn: 'Jag är' har sänt mig till eder.
Och Gud sade ytterligare till Mose: »Så skall du säga till Israels barn: HERREN, edra fäders Gud, Abrahams Gud, Isaks Gud och Jakobs Gud, har sänt mig till eder.
Detta skall vara mitt namn evinnerligen, och så skall man nämna mig från släkte till släkte.
Gå nu åstad och församla de äldste i Israel, och säg till dem: HERREN, edra fäders Gud, Abrahams, Isaks och Jakobs Gud, har uppenbarat sig för mig, och han har sagt: 'Jag har sett till eder och har sett det som vederfares eder Egypten;
därför är nu mitt ord: jag vill föra eder bort ifrån betrycket i Egypten upp till kananéernas, hetiternas, amoréernas, perisséernas, hivéernas och jebuséernas land, ett land som flyter av mjölk och honung.'
Och de skola lyssna till dina ord; och du skall tillika med de äldste i Israel gå till konungen i Egypten, och I skolen säga till honom: HERREN, hebréernas Gud, har visat sig för oss, så låt oss nu gå tre dagsresor in i öknen och offra åt HERREN, vår Gud.'
Dock vet jag att konungen i Egypten icke skall tillstädja eder att gå, icke ens när han får känna min starka hand.
Men jag skall räcka ut min hand och slå Egypten med alla slags under, som jag vill göra där; sedan skall han släppa eder.
Och jag vill låta detta folk finna nåd för egyptiernas ögon, så att I, när I dragen bort, icke skolen draga bort med tomma händer;
utan var kvinna skall av sin grannkvinna och av den främmande kvinna som bor i hennes hus begära klenoder av silver och guld, så ock kläder.
Dessa skolen I sätta på edra söner och döttrar.
Så skolen I taga byte från egyptierna.»
Mose svarade och sade: »Men om de nu icke tro mig eller lyssna till mina ord, utan säga: 'HERREN har icke uppenbarat sig för dig'?»
Då sade HERREN till honom: »Vad är det du har i din hand?»
Han svarade: »En stav.»
Han sade: »Kasta den på marken.»
När han då kastade den på marken, förvandlades den till en orm; och Mose flydde för honom.
Men HERREN sade till Mose: »Räck ut din hand och tag honom i stjärten.»
Då räckte han ut sin hand och grep honom; och han förvandlades åter till en stav i hans hand.
Och HERREN sade: »Så skola de. tro att HERREN, deras fäders Gud, Abrahams Gud, Isaks Gud och Jakobs Gud, har uppenbarat sig för dig.
Och HERREN sade ytterligare till honom: »Stick din hand i barmen.»
Och han stack sin hand i barmen.
När han sedan drog ut den, se, då var handen vit såsom snö av spetälska.
Åter sade han. »Stick din hand tillbaka i barmen.»
Och han stack sin hand tillbaka i barmen.
När han sedan drog ut den igen ur barmen, se, då var den åter lik hans övriga kropp.
Och HERREN sade: »Om de icke vilja tro dig eller akta på det första tecknet, så måste de tro det andra tecknet.
Men om de icke ens tro dessa två tecken eller lyssna till dina ord, så tag av Nilflodens vatten och gjut ut det på torra landet, så skall vattnet, som du har tagit ur floden, förvandlas till blod på torra landet.»
Då sade Mose till HERREN: »Ack I Herre, jag är ingen talför man; jag har icke varit det förut, och jag är det icke heller nu, sedan du har talat till din tjänare, ty jag har ett trögt målföre och en trög tunga.
HERREN sade till honom: »Vem har givit människan munnen, eller vem gör henne stum eller döv, seende eller blind?
Är det icke jag, HERREN?
Så gå nu åstad, jag skall vara med din mun och lära dig vad du skall tala.»
Men han sade: »Ack Herre, sänd ditt budskap med vilken annan du vill.»
Då upptändes HERRENS vrede mot Mose, och han sade: »Har du icke din broder Aron, leviten?
Jag vet att han är en man som kan tala.
Och han går nu åstad för att möta dig, och när han får se dig, skall han glädjas i sitt hjärta.
Och du skall tala till honom och lägga orden i hans mun; och jag skall vara med din mun och med hans mun, och jag skall lära eder vad I skolen göra.
Och han skall tala för dig till folket; alltså skall han vara för dig såsom mun, och du skall vara för honom såsom en gud.
Och du skall taga i din hand denna stav, med vilken du skall göra dina tecken.»
Därefter vände Mose tillbaka till sin svärfader Jeter och sade till honom: »Låt mig vända tillbaka till mina bröder i Egypten, för att se om de ännu leva.»
Jetro sade till Mose: »Gå i frid.»
Och HERREN sade till Mose i Midjan: »Vänd tillbaka till Egypten, ty alla de män äro döda, som stodo efter ditt liv.»
Då tog Mose sin hustru och sina söner och satte dem på sin åsna och for tillbaka till Egyptens land; och Mose tog Guds stav i sin hand.
Och HERREN sade till Mose: »När du nu vänder tillbaka till Egypten så se till, att du inför Farao gör alla de under som jag har givit dig makt att göra.
Men jag skall förstocka hans hjärta, så att han icke släpper folket.
Och då skall du säga till Farao: Så säger HERREN: Israel är min förstfödde son,
och jag har sagt till dig: 'Släpp min son, så att han kan hålla gudstjänst åt mig.'
Men du har icke velat släppa honom.
Därför skall jag nu dräpa din förstfödde son.
Och under resan hände sig att HERREN på ett viloställe kom emot honom och ville döda honom.
Då tog Sippora en skarp sten och skar bort förhuden på sin son och berörde honom därmed nedtill och sade: »Du är mig en blodsbrudgum.»
Så lät han honom vara.
Då sade hon åter: »Ja, en blodsbrudgum till omskärelse.»
Och HERREN sade till Aron: »Gå åstad och möt Mose i öknen.»
Då gick han åstad och träffade honom på Guds berg; och han kysste honom.
Och Mose berättade för Aron allt vad HERREN hade talat, när han sände honom, och om alla de tecken som han hade bjudit honom att göra.
Sedan gingo Mose och Aron åstad och församlade alla Israels barns äldste.
Och Aron omtalade allt vad HERREN hade talat till Mose; och han gjorde tecknen inför folkets ögon.
Då trodde folket; och när de hörde att HERREN hade sett till Israels barn, och att han hade sett deras betryck, böjde de sig ned och tillbådo.
Därefter kommo Mose och Aron och sade till Farao: »Så säger HERREN, Israels Gud: Släpp mitt folk, så att de kunna hålla högtid åt mig i öknen.»
Men Farao svarade: »Vem är HERREN, eftersom jag på hans befallning skulle släppa Israel?
Jag vet icke av HERREN och vill ej heller släppa Israel.»
Då sade de: »Hebréernas Gud har visat sig för oss.
Så låt oss nu gå tre dagsresor in i öknen och offra åt HERREN, vår Gud, för att han icke må komma över oss med pest eller med svärd.»
Men konungen i Egypten svarade dem: »Mose och Aron, varför dragen I folket ifrån dess arbete?
Gån bort till edra dagsverken.
Ytterligare sade Farao: »Folket är ju redan alltför talrikt i landet, och likväl viljen I skaffa dem frihet ifrån deras dagsverken!»
Därefter bjöd Farao samma dag fogdarna och tillsyningsmännen över folket och sade:
»I skolen icke vidare såsom förut giva folket halm till att göra tegel.
Låten dem själva gå och skaffa sig halm.
Men samma antal tegel som de förut hava gjort skolen I ändå ålägga dem, utan något avdrag; ty de äro lata, därför ropa de och säga: 'Låt oss gå och offra åt vår Gud.'
Man måste lägga tungt arbete på dessa människor, så att de därigenom få något att göra och icke akta på lögnaktigt tal.»
Då gingo fogdarna och tillsyningsmännen över folket ut och sade till folket: »Så säger Farao: Jag vill icke längre giva eder halm.
Gån själva och skaffen eder halm, var I kunnen finna sådan; men i edert arbete skall intet avdrag göras.»
Då spridde sig folket över hela Egyptens land och samlade strå för att bruka det såsom halm.
Och fogdarna drevo på dem och sade: »Fullgören edert arbete, var dag det för den dagen bestämda, likasom när man gav eder halm.»
Och Israels barns tillsyningsmän, de som Faraos fogdar hade satt över dem, fingo uppbära hugg och slag, och man sade till dem: »Varför haven I icke såsom förut fullgjort edert förelagda dagsverke i tegel, varken i går eller i dag?»
Då kommo Israels barns tillsyningsmän och ropade till Farao och sade: »Varför gör du så mot dina tjänare?
Ingen halm giver man åt dina tjänare, och likväl säger man till oss: 'Skaffen fram tegel.'
Och se, dina tjänare få nu uppbära hugg och slag, fastän skulden ligger hos ditt eget folk.»
Men han svarade: »I ären lata, ja lata ären I. Därför sägen I: 'Låt oss gå och offra åt HERREN.'
Nej, gån i stället till edert arbete.
Halm skall man icke giva eder, men det bestämda antalet tegel måsten I ändå lämna.»
Då märkte Israels barns tillsyningsmän att det var illa ställt för dem, eftersom de hade fått det svaret att de icke skulle få något avdrag i det antal tegel, som de skulle lämna för var dag.
Och när de kommo ut ifrån Farao, träffade de Mose och Aron, som stodo där för att möta dem;
och de sade till dem: »Må HERREN hemsöka eder och döma eder, eftersom I haven gjort oss förhatliga för Farao och hans tjänare och satt dem svärdet i hand till att dräpa oss.
Då vände sig Mose åter till HERREN och sade: »Herre, varför har du gjort så illa mot detta folk?
Varför har du sänt mig?
Allt ifrån den tid då jag gick till Farao för att tala i ditt namn har han ju gjort illa mot detta folk, och du har ingalunda räddat ditt folk.
Men HERREN sade till Mose: »Nu skall du få se vad jag skall göra med Farao; ty genom min starka hand skall han nödgas släppa dem, ja, han skall genom min starka hand nödgas driva dem ut ur sitt land.»
Och Gud talade till Mose och sade till honom: »Jag är HERREN.
För Abraham, Isak och Jakob uppenbarade jag mig såsom 'Gud den Allsmäktige', men under mitt namn 'HERREN' var jag icke känd av dem.
Och jag upprättade ett förbund med dem och lovade att giva dem Kanaans land, det land där de bodde såsom främlingar.
Och nu har jag hört Israels barns jämmer över att egyptierna hålla dem i träldom, och jag har kommit ihåg mitt förbund.
Säg därför till Israels barn: 'Jag är HERREN, och jag skall föra eder ut från trälarbetet hos egyptierna och rädda eder från träldomen under dem, och jag skall förlossa eder med uträckt arm och genom stora straffdomar.
Och jag skall taga eder till mitt folk och vara eder Gud; och I skolen förnimma att jag är HERREN eder Gud, han som för eder ut från trälarbetet hos egyptierna.
Och jag skall föra eder till det land som jag med upplyft hand har lovat giva åt Abraham, Isak och Jakob; det skall jag giva eder till besittning.
Jag är HERREN.'»
Detta allt sade Mose till Israels barn, men de hörde icke på Mose, av otålighet och för det hårda arbetets skull.
Därefter talade HERREN till Mose och sade:
»Gå och tala med Farao, konungen i Egypten, att han släpper Israels barn ut ur sitt land.»
Men Mose talade inför HERREN och sade: »Israels barn höra ju icke på mig; huru skulle då Farao vilja höra mig -- mig som har oomskurna läppar?»
Men HERREN talade till Mose och Aron och gav dem befallning till Israels barn och till Farao, konungen i Egypten, om att Israels barn skulle föras ut ur Egyptens land.
Dessa voro huvudmännen för deras familjer.
Rubens, Israels förstföddes, söner voro Hanok och Pallu, Hesron och Karmi.
Dessa voro Rubens släkter.
Simeons söner voro Jemuel, Jamin, Ohad, Jakin, Sohar och Saul, den kananeiska kvinnans son.
Dessa voro Simeons släkter.
Och dessa voro namnen på Levis söner, efter deras ättföljd: Gerson, Kehat och Merari.
Och Levi blev ett hundra trettiosju år gammal.
Gersons söner voro Libni och Simei, efter deras släkter.
Kehats söner voro Amram, Jishar, Hebron och Ussiel.
Och Kehat blev ett hundra trettiotre år gammal.
Meraris söner voro Maheli och Musi.
Dessa voro leviternas släkter, efter deras ättföljd.
Men Amram tog sin faders syster Jokebed till hustru, och hon födde åt honom Aron och Mose.
Och Amram blev ett hundra trettiosju år gammal.
Jishars söner voro Kora, Nefeg och Sikri.
Ussiels söner voro Misael, Elsafan och Sitri.
Och Aron tog till hustru Eliseba, Amminadabs dotter, Nahesons syster, och hon födde åt honom Nadab och Abihu, Eleasar och Itamar.
Koras söner voro Assir, Elkana och Abiasaf.
Dessa voro koraiternas släkter.
Och Eleasar, Arons son, tog en av Putiels döttrar till hustru, och hon födde åt honom Pinehas.
Dessa voro huvudmännen för leviternas familjer, efter deras släkter.
Så förhöll det sig med Aron och Mose, dem till vilka HERREN sade: »Fören Israels barn ut ur Egyptens land, efter deras härskaror.
Det var dessa som talade med Farao, konungen i Egypten, om att de skulle föra Israels barn ut ur Egypten.
Så förhöll det sig med Mose och Aron,
Och när HERREN talade till Mose i Egyptens land,
talade han så till Mose: »Jag är HERREN.
Tala till Farao, konungen i Egypten, allt vad jag talar till dig.»
Men Mose sade inför HERREN: »Se, jag har oomskurna läppar; huru skulle då Farao vilja höra på mig?»
Men HERREN sade till Mose: »Se, jag har satt dig att vara såsom en gud för Farao, och din broder Aron skall vara din profet.
Du skall tala allt vad jag bjuder dig; sedan skall din broder Aron tala med Farao om att han måste släppa Israels barn ut ur sitt land.
Men jag skall förhärda Faraos hjärta och skall göra många tecken och under i Egyptens land.
Farao skall icke höra på eder; men jag skall lägga min hand på Egypten och skall föra mina härskaror, mitt folk, Israels barn, ut ur Egyptens land, genom stora straffdomar.
Och egyptierna skola förnimma att jag är HERREN, när jag räcker ut min hand över Egypten och för Israels barn ut från dem.»
Och Mose och Aron gjorde så; de gjorde såsom HERREN hade bjudit dem.
Men Mose var åttio år gammal och Aron åttiotre år gammal, när de talade med Farao.
Och HERREN talade till Mose och Aron och sade:
»När Farao talar till eder och säger: 'Låten oss se något under', då skall du säga till Aron: 'Tag din stav och kasta den inför Farao', så skall den bliva en stor orm.»
Då gingo Mose och Aron till Farao och gjorde såsom HERREN hade bjudit.
Aron kastade sin stav inför Farao och hans tjänare, och den blev en stor orm.
Då kallade också Farao till sig sina vise och trollkarlar; och dessa, de egyptiska spåmännen, gjorde ock detsamma genom sina hemliga konster:
de kastade var och en sin stav, och dessa blevo stora ormar.
Men Arons stav uppslukade deras stavar.
Dock förblev Faraos hjärta förstockat, och han hörde icke på dem, såsom HERREN hade sagt.
Därefter sade HERREN till Mose: »Faraos hjärta är tillslutet, han vill icke släppa folket.
Gå till Farao i morgon bittida -- han går nämligen då ut till vattnet -- och ställ dig i hans väg, på stranden av Nilfloden.
Och tag i din hand staven som förvandlades till en orm.
Och säg till honom: HERREN, hebréernas Gud, sände mig till dig och lät säga dig: 'Släpp mitt folk, så att de kunna hålla gudstjänst åt mig i öknen.'
Men se, du har hitintills icke velat höra.
Därför säger nu HERREN så: 'Härav skall du förnimma att jag är HERREN: se, med staven som jag håller i min hand vill jag slå på vattnet i Nilfloden, och då skall det förvandlas till blod.
Och fiskarna i floden skola dö, och floden skall bliva stinkande, så att egyptierna skola vämjas vid att dricka vatten ifrån floden.'»
Och HERREN sade till Mose: »Säg till Aron: Tag din stav, och räck ut din hand över egyptiernas vatten, över deras strömmar, kanaler och sjöar och alla andra vattensamlingar, så skola de bliva blod; över hela Egyptens land skall vara blod, både i träkärl och i stenkärl.»
Och Mose och Aron gjorde såsom HERREN hade bjudit.
Han lyfte upp staven och slog vattnet i Nilfloden inför Faraos och hans tjänares ögon; då förvandlades allt vatten floden till blod.
Och fiskarna i floden dogo, och floden blev stinkande, så att egyptierna icke kunde dricka vatten ifrån floden; och blodet var över hela Egyptens land.
Men de egyptiska spåmännen gjorde detsamma genom sina hemliga konster.
Så förblev Faraos hjärta förstockat, och han hörde icke på dem, såsom HERREN hade sagt.
Och Farao vände om och gick hem och aktade icke heller på detta.
Men i hela Egypten grävde man runt omkring Nilfloden efter vatten till att dricka; ty vattnet i floden kunde man icke dricka.
Och så förgingo sju dagar efter det att HERREN hade slagit Nilfloden.
Därefter sade HERREN till Mose: »Gå till Farao och säg till honom: Så säger HERREN: Släpp mitt folk, så att de kunna hålla gudstjänst åt mig.
Men om du icke vill släppa dem, se, då skall jag hemsöka hela ditt land med paddor.
Nilfloden skall frambringa ett vimmel av paddor, och de skola stiga upp och komma in i ditt hus och i din sovkammare och upp i din säng, och in i dina tjänares hus och bland ditt folk, och i dina bakugnar och baktråg.
Ja, på dig själv och ditt folk och alla dina tjänare skola paddorna stiga upp.»
Och HERREN sade till Mose: »Säg till Aron: Räck ut din hand med din stav över strömmarna, kanalerna och sjöarna, och låt så paddor stiga upp över Egyptens land.»
Då räckte Aron ut sin hand över Egyptens vatten, och paddor stego upp och övertäckte Egyptens land.
Men spåmännen gjorde detsamma genom sina hemliga konster och läto paddor stiga upp över Egyptens land.
Då kallade Farao Mose och Aron till sig och sade: »Bedjen till HERREN, att han tager bort paddorna från mig och mitt folk, så skall jag släppa folket, så att de kunna offra åt HERREN.»
Mose sade till Farao: »Dig vare tillstatt att förelägga mig en tid inom vilken jag, genom att bedja för dig och dina tjänare och ditt folk, skall skaffa bort paddorna från dig och dina hus, så att de finnas kvar allenast i Nilfloden.
Han svarade: »Till i morgon.»
Då sade han: »Må det ske såsom du har sagt, så att du får förnimma att ingen är såsom HERREN, vår Gud.
Paddorna skola vika bort ifrån dig och dina hus och ifrån dina tjänare och ditt folk och skola finnas kvar allenast i Nilfloden.»
Så gingo Mose och Aron ut ifrån Farao.
Och Mose ropade till HERREN om hjälp mot paddorna som han hade låtit komma över Farao.
Och HERREN gjorde såsom Mose hade begärt: paddorna dogo och försvunno ifrån husen, gårdarna och fälten.
Och man kastade dem tillsammans i högar, här en och där en; och landet uppfylldes av stank.
Men när Farao såg att han hade fått lättnad, tillslöt han sitt hjärta och hörde icke på dem, såsom HERREN hade sagt.
Därefter sade HERREN till Mose: »Säg till Aron: Räck ut din stav och slå i stoftet på jorden, så skall därav bliva mygg i hela Egyptens land.»
Och de gjorde så: Aron räckte ut sin hand med sin stav och slog i stoftet på jorden; då kom mygg på människor och boskap.
Av allt stoft på marken blev mygg i hela Egyptens land.
Och spåmännen ville göra detsamma genom sina hemliga konster och försökte skaffa fram mygg, men de kunde icke.
Och myggen kom på människor och boskap.
Då sade spåmännen till Farao: »Detta är Guds finger.»
Men Faraos hjärta förblev förstockat, och han hörde icke på dem, såsom HERREN hade sagt.
Därefter sade HERREN till Mose: »Träd i morgon bittida fram inför Farao -- han går nämligen då ut till vattnet -- och säg till honom: så säger HERREN: Släpp mitt folk, så att de kunna hålla guds tjänst åt mig.
Ty om du icke släpper mitt folk, de, då skall jag sända svärmar av flugor över dig och dina tjänare och ditt folk och dina hus, så att egyptiernas hus skola bliva uppfyllda av flugsvärmar, ja, själva marken på vilken de stå.
Men på den dagen skall jag göra ett undantag för landet Gosen, där mitt folk bor, så att inga flugsvärmar skola finnas där, på det att du må förnimma att jag är HERREN här i landet.
Så skall jag förlossa mitt folk och göra en åtskillnad mellan mitt folk och ditt.
I morgon skall detta tecken ske.»
Och HERREN gjorde så: stora flugsvärmar kommo in i Faraos och i hans tjänares hus; och överallt i Egypten blev landet fördärvat av flugsvärmarna.
Då kallade Farao Mose och Aron till sig och sade: »Gån åstad och offren åt eder Gud här i landet.»
Men Mose svarade: »Det går icke an att vi göra så; ty vi offra åt HERREN, vår Gud, sådant som för egyptierna är en styggelse.
Om vi nu inför egyptiernas ögon offra sådant som för dem är en styggelse, skola de säkert stena oss.
Så låt oss nu gå tre dagsresor in i öknen och offra åt HERREN, vår Gud, såsom han befaller oss.»
Då sade Farao: »Jag vill släppa eder, så att I kunnen offra åt HERREN, eder Gud, i öknen; allenast mån I icke gå alltför långt bort.
Bedjen för mig.
Mose svarade: »Ja, när jag kommer ut från dig, skall jag bedja till HERREN, så att flugsvärmarna i morgon vika bort ifrån Farao, ifrån hans tjänare och hans folk.
Allenast må Farao icke mer handla svikligt och vägra att släppa folket, så att de kunna offra åt HERREN.
Och Mose gick ut ifrån Farao och bad till HERREN.
Och HERREN gjorde såsom Mose sade begärt: han skaffade bort flugsvärmarna ifrån Farao, ifrån hans tjänare och hans folk, så att icke en enda fluga blev kvar.
Men Farao tillslöt sitt hjärta också denna gång och släppte icke folket.
Därefter sade HERREN till Mose: »Gå till Farao och tala till honom: Så säger HERREN, hebréernas Gud: Släpp mitt folk, så att de kunna hålla gudstjänst åt mig.
Ty om du icke vill släppa dem, utan kvarhåller dem längre,
se, då skall HERRENS hand med en mycket svår pest komma över din boskap på marken, över hästar, åsnor och kameler, över fäkreatur och får.
Men HERREN skall därvid göra en åtskillnad mellan israeliternas boskap och egyptiernas, så att intet av de djur som tillhöra Israels barn skall dö.»
Och HERREN bestämde en tid och sade: »I morgon skall HERREN göra så i landet.»
Och dagen därefter gjorde HERREN så, och all egyptiernas boskap dog.
Men av Israels barns boskap dog icke ett enda djur;
när Farao sände och hörde efter, se, då hade icke så mycket som ett enda djur av Israels boskap dött.
Men Faraos hjärta var tillslutet, och han släppte icke folket
Därefter sade HERREN till Mose och Aron: »Tagen edra händer fulla med sot ur smältugnen, och må sedan Mose strö ut det, upp mot himmelen, inför Faraos ögon,
så skall därav bliva ett damm över hela Egyptens land, och därav skola uppstå bulnader, som slå ut med blåsor, på människor och boskap i hela Egyptens land.»
Då togo de sot ur smältugnen och trädde inför Farao, och Mose strödde ut det, upp mot himmelen; och därav uppstodo bulnader, som slogo ut med blåsor, på människor och boskap.
Och spåmännen kunde icke hålla stånd mot Mose för bulnadernas skull, ty bulnader uppstodo på spåmännen såväl som på alla andra egyptier.
Men HERREN förstockade Faraos hjärta, så att han icke hörde på dem, såsom HERREN hade sagt till Mose.
Därefter sade HERREN till Mose: »Träd i morgon bittida fram inför Farao och säg till honom: Så säger HERREN, hebréernas Gud: Släpp mitt folk, så att de kunna hålla gudstjänst åt mig.
Annars skall jag nu sända alla mina hemsökelser över dig själv och över dina tjänare och ditt folk, på det att du må förnimma att ingen är såsom jag på hela jorden.
Ty jag hade redan räckt ut min land för att slå dig och ditt folk med pest, så att du skulle bliva utrotad från jorden;
men jag skonade dig, just därför att jag ville låta min kraft bliva uppenbarad för dig och mitt namn bliva förkunnat på hela jorden.
Om du ytterligare lägger hinder i vägen för mitt folk och icke släpper dem,
se, då skall jag i morgon vid denna tid låta ett mycket svårt hagel komma, sådant att dess like icke har varit i Egypten, allt ifrån den dag dess grund blev lagd ända till nu.
Så sänd nu bort och låt bärga din boskap och allt vad du annars har ute på marken.
Ty alla människor och all boskap som då finnas ute på marken och icke hava kommit under tak, de skola träffas av haglet och bliva dödade.»
Den som nu bland Faraos tjänare fruktade HERRENS ord, han lät sina tjänare och sin boskap söka skydd i husen;
men den som icke aktade på HERRENS ord, han lät sina tjänare och sin boskap bliva kvar ute på marken.
Och HERREN sade till Mose: »Räck din hand upp mot himmelen, så skall hagel falla över hela Egyptens land, över människor och boskap och över alla markens örter i Egyptens land.»
Då räckte Mose sin stav upp mot himmelen, och HERREN lät det dundra och hagla, och eld for ned mot jorden, så lät HERREN hagel komma över Egyptens land.
Och det haglade, och bland hagelskurarna flammade eld; och haglet var så svårt, att dess like icke hade varit i hela Egyptens land från den tid det blev befolkat.
Och i hela Egyptens land slog haglet ned allt som fanns på marken, både människor och djur; och haglet slog ned alla markens örter och slog sönder alla markens träd.
Allenast i landet Gosen, där Israels barn voro, haglade det icke.
Då sände Farao och lät kalla till sig Mose och Aron och sade till dem: »Jag har syndat denna gång.
Det är HERREN som är rättfärdig; jag och mitt folk hava gjort orätt.
Bedjen till HERREN, ty hans dunder och hagel har varat länge nog; så skall jag släppa eder, och I skolen icke behöva bliva kvar längre.»
Mose svarade honom: »När jag kommer ut ur staden, skall jag uträcka mina händer till HERREN; då skall dundret upphöra och intet hagel mer komma, på det att du må förnimma att landet är HERRENS.
Dock vet jag väl att du och dina tjänare ännu icke frukten för HERREN Gud.»
Så slogos då linet och kornet ned, ty kornet hade gått i ax och linet stod i knopp;
men vetet och spälten slogos icke ned, ty de äro sensäd.
Och Mose gick ifrån Farao ut ur staden och uträckte sina händer till HERREN; och dundret och haglet upphörde, och regnet strömmade icke mer ned på jorden.
Men när Farao såg att regnet och haglet och dundret hade upphört, framhärdade han i sin synd och tillslöt sitt hjärta, han själv såväl som hans tjänare.
Så förblev Faraos hjärta förstockat, och han släppte icke Israels barn, såsom HERREN hade sagt genom Mose.
Därefter sade HERREN till Mose: »Gå till Farao; ty jag har tillslutit hans och hans tjänares hjärtan, för att jag skulle göra dessa mina tecken mitt ibland dem,
och för att du sedan skulle kunna förtälja för din son och din sonson vilka stora gärningar jag har utfört bland egyptierna, och vilka tecken jag har gjort bland dem, så att I förnimmen att jag är HERREN.»
Då gingo Mose och Aron till Farao och sade till honom: »Så säger HERREN, hebréernas Gud: Huru länge vill du vara motsträvig och icke ödmjuka dig inför mig?
Släpp mitt folk, så att de kunna hålla gudstjänst åt mig.
Ty om du icke vill släppa mitt folk, se, då skall jag i morgon låta gräshoppor komma över ditt land.
Och de skola övertäcka marken så att man icke kan se marken; och de skola äta upp återstoden av den kvarleva som har blivit över åt eder efter haglet, och de skola aväta alla edra träd, som växa på marken.
Och dina hus skola bliva uppfyllda av dem, så ock alla dina tjänares hus och alla egyptiers hus, så att dina fäder och dina faders fäder icke hava sett något sådant, från den dag de blevo till på jorden ända till denna dag.»
Och han vände sig om och gick ut ifrån Farao.
Men Faraos tjänare sade till honom: »Huru länge skall denne vara oss till förfång?
Släpp männen, så att de kunna hålla gudstjänst åt HERREN, sin Gud.
Inser du icke ännu att Egypten bliver fördärvat?»
Då hämtade man Mose och Aron tillbaka till Farao.
Och han sade till dem: »I mån gå åstad och hålla gudstjänst åt HERREN, eder Gud.
Men vilka äro nu de som skola gå?»
Mose svarade: »Vi vilja gå både unga och gamla; vi vilja gå med söner och döttrar, med får och fäkreatur; ty en HERRENS högtid skola vi hålla.»
Då sade han till dem: »Må HERREN: vara med eder lika visst som jag släpper eder med edra kvinnor och barn!
Där ser man att I haven ont i sinnet!
Nej; I män mån gå åstad och hålla gudstjänst åt HERREN; det var ju detta som I begärden.»
Och man drev dem ut ifrån Farao.
Och HERREN sade till Mose: »Räck ut din hand över Egyptens land, så att gräshoppor komma över Egyptens land och äta upp alla örter i landet, allt vad haglet har lämnat kvar.»
Då räckte Mose ut sin stav över Egyptens land, och HERREN lät en östanvind blåsa över landet hela den dagen och hela natten; och när det blev morgon, förde östanvinden gräshopporna fram med sig.
Och gräshopporna kommo över hela Egyptens land och slogo i stor mängd ned över hela Egyptens område; en sådan myckenhet av gräshoppor hade aldrig tillförne kommit och skall icke heller hädanefter komma.
De övertäckte hela marken, så att marken blev mörk; och de åto upp alla örter i landet och all frukt på träden, allt som haglet hade lämnat kvar; intet grönt blev kvar på träden eller på markens örter i hela Egyptens land.
Då kallade Farao med hast Mose och Aron till sig och sade: »Jag har syndat mot HERREN, eder Gud, och mot eder.
Men förlåt nu min synd denna enda gång; och bedjen till HERREN, eder Gud, att han avvänder allenast denna dödsplåga ifrån mig.»
Då gick han ut ifrån Farao och bad till HERREN.
Och HERREN vände om vinden och lät en mycket stark västanvind komma; denna fattade i gräshopporna och kastade dem i Röda havet, så att icke en enda gräshoppa blev kvar inom Egyptens hela område.
Men HERREN förstockade Faraos hjärta, så att han icke släppte Israels barn.
Därefter sade HERREN till Mose: »Räck din hand upp mot himmelen, så skall över Egyptens land komma ett sådant mörker, att man kan taga på det.»
Då räckte Mose sin hand upp mot himmelen, och ett tjockt mörker kom över hela Egyptens land i tre dagar.
Ingen kunde se den andre, och ingen kunde röra sig från sin plats i tre dagar.
Men alla Israels barn hade ljust där de bodde.
Då kallade Farao Mose till sig och sade: »Gån åstad och hållen gudstjänst åt HERREN; låten allenast edra får och fäkreatur bliva kvar.
Också edra kvinnor och barn må gå med eder.»
Men Mose sade: »Du måste ock låta oss få slaktoffer och brännoffer att offra åt HERREN, vår Gud.
Också vår boskap måste gå med oss, och icke en klöv får bliva kvar; ty därav måste vi taga det varmed vi skola hålla gudstjänst åt HERREN, vår Gud.
Och förrän vi komma dit, veta vi själva icke vad vi böra offra åt HERREN.»
Men HERREN förstockade Faraos hjärta, så att han icke ville släppa dem.
Och Farao sade till honom: »Gå bort ifrån mig, och tag dig till vara för att ännu en gång komma inför mitt ansikte; ty på den dag du kommer inför mitt ansikte skall du dö.»
Mose svarade: »Du har talat rätt; jag skall icke vidare komma inför ditt ansikte.»
Därefter sade HERREN till Mose: »Ännu en plåga skall jag låta komma över Farao och över Egypten; sedan skall han släppa eder härifrån; ja, han skall till och med driva eder ut härifrån, när han släpper eder.
Så tala nu till folket, och säg att var och en av dem, man såväl som kvinna, skall av sin nästa begära klenoder av silver och guld.»
Och HERREN lät folket finna nåd för egyptiernas ögon.
Ja, mannen Mose hade stort anseende i Egyptens land, både hos Faraos tjänare och hos folket.
Och Mose sade: »Så säger HERREN: Vid midnattstid skall jag gå fram genom Egypten.
Och då skall allt förstfött i Egyptens land dö, från den förstfödde hos Farao, som sitter på tronen, ända till den förstfödde hos tjänstekvinnan, som arbetar vid handkvarnen, så ock allt förstfött ibland boskapen.
Och ett stort klagorop skall upphävas i hela Egyptens land, sådant att dess like aldrig har varit hört och aldrig mer skall höras.
Men icke en hund skall gläfsa mot någon av Israels barn, varken mot människor eller mot boskap.
Så skolen I förnimma att HERREN gör en åtskillnad mellan Egypten och Israel.
Då skola alla dina tjänare här komma ned till mig och buga sig för mig och säga: 'Drag ut, du själv med allt folket som följer dig.'
Och sedan skall jag draga ut.»
Därefter gick han bort ifrån Farao i vredesmod.
Men HERREN sade till Mose: »Farao skall neka att höra eder, på det att jag må låta många under ske i Egyptens land.»
Och Mose och Aron gjorde alla dessa under inför Farao; men HERREN förstockade Faraos hjärta, så att han icke släppte Israels barn ut ur sitt land.
Och HERREN talade till Mose och Aron i Egyptens land och sade:
Denna månad skall hos eder vara den främsta månaden, den skall hos eder vara den första av årets månader.
Talen till Israels hela menighet och sägen: På tionde dagen i denna månad skall var husfader taga sig ett lamm, så att vart hushåll får ett lamm.
Men om hushållet är för litet till ett lamm, så skola husfadern och hans närmaste granne taga ett lamm tillsammans, efter personernas antal.
För vart lamm skolen I beräkna ett visst antal, i mån av vad var och en äter.
Ett felfritt årsgammalt lamm av hankön skolen I utvälja; av fåren eller av getterna skolen I taga det.
Och I skolen förvara det intill fjortonde dagen i denna månad; då skall man -- Israels hela församlade menighet -- slakta det vid aftontiden.
Och man skall taga av blodet och stryka på båda dörrposterna och på övre dörrträet i husen där man äter det.
Och man skall äta köttet samma natt; det skall vara stekt på eld, och man skall äta det med osyrat bröd jämte bittra örter.
I skolen icke äta något därav rått eller kokt i vatten, utan det skall vara stekt på eld, med huvud, fötter och innanmäte.
Och I skolen icke lämna något därav kvar till morgonen; skulle något därav bliva kvar till morgonen, skolen I bränna upp det i eld.
Och I skolen äta det så: I skolen vara omgjordade kring edra länder, hava edra skor på fötterna och edra stavar i händerna.
Och I skolen äta det med hast.
Detta är HERRENS Påsk.
Ty jag skall på den natten gå fram genom Egyptens land och slå allt förstfött i Egyptens land, både människor och boskap; och över Egyptens alla gudar skall jag hålla dom; jag är HERREN.
Och blodet skall vara ett tecken, eder till räddning, på de hus i vilka I ären; ty när jag ser blodet, skall jag gå förbi eder.
Och ingen hemsökelse skall drabba eder med fördärv, när jag slår Egyptens land.
Och I skolen hava denna dag till en åminnelsedag och fira den såsom en HERRENS högtid.
Såsom en evärdlig stiftelse skolen I fira den, släkte efter släkte.
I sju dagar skolen I äta osyrat bröd; redan på första dagen skolen I skaffa bort all surdeg ur edra hus.
Ty var och en som äter något syrat, från den första dagen till den sjunde, han skall utrotas ur Israel.
På den första dagen skolen I hålla en helig sammankomst; I skolen ock på den sjunde dagen hålla en helig sammankomst.
På dem skall intet arbete göras; allenast det som var och en behöver till mat, det och intet annat må av eder tillredas.
Och I skolen hålla det osyrade brödets högtid, eftersom jag på denna samma dag har fört edra härskaror ut ur Egyptens land.
Därför skolen I, släkte efter släkte, hålla denna dag såsom en evärdlig stiftelse.
I första månaden, på fjortonde dagen i månaden, om aftonen, skolen I äta osyrat bröd, och I skolen fortfara därmed ända till aftonen på tjuguförsta dagen i månaden.
I sju dagar må ingen surdeg finnas i edra hus; ty var och en son äter något syrligt, han skall utrotas ur Israels menighet, evad han är främling eller inföding i landet.
Intet syrligt skolen I äta; var I än ären bosatta skolen I äta osyrat bröd.
Och Mose kallade till sig alla de äldste i Israel och sade till dem: »Begiven eder hem, och tagen eder ett lamm för vart hushåll och slakten påskalammet.
Och tagen en knippa isop och doppen den i blodet som är i skålen, och bestryken det övre dörr träet och båda dörrposterna med blodet som är i skålen; och ingen av eder må gå ut genom sin hus dörr intill morgonen.
Ty HERREN skall gå fram för att hemsöka Egypten; men när ha ser blodet på det övre dörrträet och på de två dörrposterna, skall HERREN gå förbi dörren och icke tillstädja Fördärvaren att komma i i edra hus och hemsöka eder.
Detta skolen I hålla; det skall vara en stadga för dig och dina barn till evärdlig tid.
Och när I kommen in i det land som HERREN skall giva åt eder, såsom han har lovat, skolen I hålla denna gudstjänst.
När då edra barn fråga eder: 'Vad betyder denna eder gudstjänst?',
skolen I svara: 'Det är ett påskoffer åt HERREN, därför att han gick förbi Israels barns hus i Egypten, när han hemsökte Egypten, men skonade våra hus.'»
Då böjde folket sig ned och tillbad.
Och Israels barn gingo åstad och gjorde så; de gjorde såsom HERREN hade bjudit Mose och Aron.
Och vid midnattstiden slog HERREN allt förstfött i Egyptens land, från den förstfödde hos Farao, som satt på tronen, ända till den förstfödde hos fången, som satt i fängelset, så ock allt förstfött ibland boskapen.
Då stod Farao upp om natten jämte alla sina tjänare och alla egyptier, och ett stort klagorop upphävdes i Egypten; ty intet hus fanns, där icke någon död låg.
Och han kallade Mose och Aron till sig om natten och sade: »Stån upp och dragen ut från mitt folk, I själva och Israels barn; och gån åstad och hållen gudstjänst åt HERREN, såsom I haven begärt.
Tagen ock edra får och edra fäkreatur, såsom I haven begärt, och gån åstad, och välsignen därvid mig.»
Och egyptierna trängde på folket för att med hast få dem ut ur landet, ty de tänkte: »Eljest dö vi allasammans.»
Och folket tog med sig sin deg, innan den ännu hade blivit syrad; de togo sina baktråg och lindade in dem i mantlarna och buro dem på sina axlar.
Och Israels barn hade gjort såsom Mose sade: de hade av egyptierna begärt deras klenoder av silver och guld, så ock kläder.
Och HERREN hade låtit folket finna nåd för egyptiernas ögon, så att de gåvo dem vad de begärde.
Så togo de byte från egyptierna.
Och Israels barn bröto upp och drogo från Rameses till Suckot, vid pass sex hundra tusen män till fots, förutom kvinnor och barn.
En hop folk av allahanda slag drog ock åstad med dem, därtill får och fäkreatur, boskap i stor myckenhet.
Och av degen som de hade fört med sig ur Egypten bakade de osyrade kakor, ty den hade icke blivit syrad; de hade ju drivits ut ur Egypten utan att få dröja; ej heller hade de kunnat tillreda någon reskost åt sig.
Men den tid Israels barn hade bott i Egypten var fyra hundra trettio år.
Just på den dag då de fyra hundra trettio åren voro förlidna drogo alla HERRENS härskaror ut ur Egyptens land.
En HERRENS vakenatt var detta, när han skulle föra dem ut ur Egyptens land; denna samma natt är HERRENS, en högtidsvaka för alla Israels barn, släkte efter släkte.
Och HERREN sade till Mose och Aron: »Detta är stadgan om påskalammet: Ingen utlänning skall äta därav;
men en träl som är köpt för penningar må äta därav, sedan du ha omskurit honom.
En inhysesman och en legodräng må icke äta därav.
I ett och samma hus skall det ätas; du skall icke föra något av köttet ut ur huset, och intet ben skolen I sönderslå därpå.
Israels hela menighet skall iakttaga detta.
Och om någon främling bor hos dig och vill hålla HERRENS påskhögtid, så skall allt mankön hos honom omskäras, och sedan må han komma och hålla den; han skall då vara såsom en inföding i landet.
Men ingen oomskuren må äta därav.
En och samma lag skall gälla för infödingen och för främlingen som bor ibland eder.»
Och alla Israels barn gjorde så; de gjorde såsom HERREN hade bjudit Mose och Aron.
Så förde då HERREN på denna samma dag Israels barn ut ur Egyptens land, efter deras härskaror.
Och HERREN talade till Mose och sade:
»Helga åt mig allt förstfött, allt hos Israels barn, som öppnar moderlivet, evad det är människor eller boskap; mig tillhör det.
Och Mose sade till folket: »Kommen ihåg denna dag, på vilken I haven dragit ut ur Egypten, ur träldomshuset; ty med stark hand har HERREN fört eder ut därifrån.
Fördenskull må intet syrat ätas.
På denna dag i månaden Abib dragen I nu ut.
Och när HERREN låter dig komma in i kananéernas, hetiternas, amoréernas, hivéernas och jebuséernas land, som han med ed har lovat dina fäder att giva dig, ett land som flyter av mjölk och honung, då skall du hålla denna gudstjänst i denna månad:
I sju dagar skall du äta osyrat bröd, och på sjunde dagen skall hållas en HERRENS högtid.
Under de sju dagarna skall man äta osyrat bröd; intet syrat skall man se hos dig, ej heller skall man se någon surdeg hos dig, i hela ditt land.
Och du skall på den dagen berätta för din son och säga: 'Sådant gör jag av tacksamhet för vad HERREN gjorde med mig, när jag drog ut ur Egypten.'
Och det skall vara för dig såsom ett tecken på din hand och såsom ett påminnelsemärke på din panna, för att HERRENS lag må vara i din mun; ty med stark hand har HERREN fört dig ut ur Egypten.
Och denna stadga skall du hålla på bestämd tid, år efter år.
Och när HERREN låter dig komma in i kananéernas land, såsom han med ed har lovat dig och dina fäder, och giver det åt dig,
då skall du överlämna åt HERREN allt det som öppnar moderlivet.
Allt som öppnar moderlivet av det som födes bland din boskap skall, om det är hankön, höra HERREN till.
Men allt bland åsnor som öppnar moderlivet skall du lösa med ett får, och om du icke vill lösa det, skall du krossa nacken på det.
Och allt förstfött av människa bland dina söner skall du lösa.
Och när din son i framtiden frågar dig: 'Vad betyder detta?', skall du svara honom så: 'Med stark hand har HERREN fört oss ut ur Egypten, ur träldomshuset;
ty då Farao i sin hårdnackenhet icke ville släppa oss, dräpte HERREN allt förstfött i Egyptens land, det förstfödda såväl ibland människor som ibland boskap.
Därför offrar jag åt HERREN allt som öppnar moderlivet och är hankön, och allt förstfött bland mina söner löser jag.'
Och det skall vara såsom ett tecken på din hand och såsom ett märke på din panna; ty med stark hand har HERREN fört oss ut ur Egypten.»
När Farao nu hade släppt folket, förde Gud dem icke på den väg som gick igenom filistéernas land, fastän denna var den genaste; ty Gud tänkte att folket, när det fick se krig hota, kunde ångra sig och vända tillbaka till Egypten;
därför lät Gud folket taga en omväg genom öknen åt Röda havet till.
Och Israels barn drogo väpnade upp ur Egyptens land.
Och Mose tog med sig Josefs ben; ty denne hade tagit en ed av Israels barn och sagt: »När Gud ser till eder, fören då mina ben härifrån med eder.»
Så bröto de upp från Suckot och lägrade sig i Etam, där öknen begynte.
Och HERREN gick framför dem, om dagen i en molnstod, för att leda dem på vägen, och om natten i en eldstod, för att lysa dem; så kunde de tåga både dag och natt.
Molnstoden upphörde icke om dagen att gå framför folket, ej heller eldstoden om natten.
Och HERREN talade till Mose och sade:
»Säg till Israels barn att de skola vända om och lägra sig framför Pi-Hahirot, mellan Migdol och havet; mitt framför Baal-Sefon skolen I lägra eder vid havet.
Men Farao skall tänka att Israels barn hava farit vilse i landet och blivit instängda i öknen.
Och jag skall förstocka Faraos hjärta, så att han förföljer dem; och jag skall förhärliga mig på Farao och hela hans här, på det att egyptierna må förnimma att jag är HERREN.»
Och de gjorde så.
Då man nu berättade för konungen i Egypten att folket hade flytt, förvandlades Faraos och hans tjänares hjärtan mot folket, och de sade: »Huru illa gjorde vi icke, när vi släppte Israel, så att de nu icke mer skola tjäna oss!»
Och han lät spänna för sina vagnar och tog sitt folk med sig;
han tog sex hundra utvalda vagnar, och alla vagnar som eljest funnos i Egypten, och kämpar på dem alla.
Ty HERREN förstockade Faraos, den egyptiske konungens, hjärta, så att han förföljde Israels barn, när de nu drogo ut med upplyft hand.
Och egyptierna, alla Faraos hästar, vagnar och ryttare och hela hans här, förföljde dem och hunno upp dem, där de voro lägrade vid havet, vid Pi-Hahirot, framför Baal-Sefon.
När så Farao var helt nära, lyfte Israels barn upp sina ögon och fingo se att egyptierna kommo tågande efter dem.
Då blevo Israels barn mycket förskräckta och ropade till HERREN.
Och de sade till Mose: »Funnos då inga gravar i Egypten, eftersom du har fört oss hit till att dö i öknen?
Huru illa gjorde du icke mot oss, när du förde oss ut ur Egypten!
Var det icke det vi sade till dig i Egypten?
Vi sade ju: 'Låt oss vara, så att vi få tjäna egyptierna.'
Ty det vore oss bättre att tjäna egyptierna än att dö i öknen.»
Då svarade Mose folket: »Frukten icke; stån fasta, så skolen I se vilken frälsning HERREN i dag skall bereda eder; ty aldrig någonsin skolen I mer få se egyptierna så, som I sen dem i dag.
HERREN skall strida för eder, och I skolen vara stilla därvid.»
Och HERREN sade till Mose: »Varför ropar du till mig?
Säg till Israels barn att de draga vidare.
Men lyft du upp din stav, och räck ut din hand över havet, och klyv det itu, så att Israels barn kunna gå mitt igenom havet på torr mark.
Och se, jag skall förstocka egyptiernas hjärtan, så att de följa efter dem; och jag skall förhärliga mig på Farao och hela hans här, på hans vagnar och ryttare.
Och egyptierna skola förnimma att jag är HERREN, när jag förhärligar mig på Farao, på hans vagnar och ryttare.»
Och Guds ängel, som hade gått framför Israels här, flyttade sig nu och gick bakom dem; molnstoden, som hade gått framför dem, flyttade sig och tog plats bakom dem.
Den kom så emellan egyptiernas här och Israels här; och molnet var där med mörker, men tillika upplyste det natten.
Så kunde den ena hären icke komma inpå den andra under hela natten.
Och Mose räckte ut sin hand över havet; då drev HERREN undan havet genom en stark östanvind som blåste hela natten, och han gjorde så havet till torrt land; och vattnet klövs itu.
Och Israels barn gingo mitt igenom havet på torr mark, under det att vattnet stod såsom en mur till höger och till vänster om dem.
Och egyptierna, alla Faraos hästar, vagnar och ryttare, förföljde dem och kommo efter dem ut till mitten av havet.
Men när morgonväkten var inne, blickade HERREN på egyptiernas här ur eldstoden och molnskyn och sände förvirring i egyptiernas här;
och han lät hjulen falla ifrån deras vagnar, så att det blev dem svårt att komma framåt.
Då sade egyptierna: »Låt oss fly för Israel, ty HERREN strider för dem mot egyptierna.»
Men HERREN sade till Mose: »Räck ut din hand över havet, så att vattnet vänder tillbaka och kommer över egyptierna, över deras vagnar och ryttare.»
Då räckte Mose ut sin hand över havet, och mot morgonen vände havet tillbaka till sin vanliga plats, och egyptierna som flydde möttes därav; och HERREN kringströdde egyptierna mitt i havet.
Och vattnet som vände tillbaka övertäckte vagnarna och ryttarna, hela Faraos här, som hade kommit efter dem ut i havet; icke en enda av dem kom undan.
Men Israels barn gingo på torr mark mitt igenom havet, och vattnet stod såsom en mur till höger och till vänster om dem.
Så frälste HERREN på den dagen Israel från egyptiernas hand, och Israel såg egyptierna ligga döda på havsstranden.
Och när Israel såg huru HERREN hade bevisat sin stora makt på egyptierna, fruktade folket HERREN; och de trodde på HERREN och på hans tjänare Mose.
Då sjöngo Mose och Israels barn denna lovsång till HERRENS ära; de sade: »Jag vill sjunga till HERRENS ära, ty högt är han upphöjd.
Häst och man störtade han i havet.
HERREN är min starkhet och min lovsång, Och han blev mig till frälsning.
Han är min Gud, jag vill ära honom, min faders Gud, jag vill upphöja honom.
HERREN är en stridsman, 'HERREN' är hans namn.
Faraos vagnar och härsmakt kastade han i havet, hans utvalda kämpar dränktes i Röda havet.
De övertäcktes av vattenmassor, sjönko i djupet såsom stenar.
Din högra hand, HERRE, du härlige och starke, din högra hand, HERRE, krossar fienden.
Genom din stora höghet slår du ned dina motståndare; du släpper lös din förgrymmelse, den förtär dem såsom strå.
För en fnysning av din näsa uppdämdes vattnen, böljorna reste sig och samlades hög, vattenmassorna stelnade i havets djup.
Fienden sade: 'Jag vill förfölja dem, hinna upp dem, jag vill utskifta byte, släcka min hämnd på dem; jag vill draga ut mitt svärd, min hand skall förgöra dem.'
Du andades på dem, då övertäckte dem havet; de sjönko såsom bly i de väldiga vattnen.
Vilken bland gudar liknar dig, HERRE?
Vem är dig lik, du härlige och helige, du fruktansvärde och högtlovade, du som gör under?
Du räckte ut din högra hand, då uppslukades de av jorden.
Men du ledde med din nåd det folk du hade förlossat, du förde dem med din makt till din heliga boning.
Folken hörde det och måste då darra, av ångest grepos Filisteens inbyggare.
Då förskräcktes Edoms furstar, Moabs hövdingar grepos av bävan, alla Kanaans inbyggare försmälte av ångest.
Ja, över dem faller förskräckelse och fruktan; för din arms väldighet stå de såsom förstenade, medan ditt folk tågar fram, o HERRE medan det tågar fram, det folk du har förvärvat.
Du för dem in och planterar dem på din arvedels berg, på den plats, o HERRE, som du har gjort till din boning, i den helgedom, Herre, som dina händer hava berett.
HERREN är konung alltid och evinnerligen!»
Ty när Faraos hästar med hans vagnar och ryttare hade kommit ned i havet, lät HERREN havets vatten vända tillbaka och komma över dem, sedan Israels barn på torr mark hade gått mitt igenom havet.
Och profetissan Mirjam, Arons syster, tog en puka i sin hand, och alla kvinnorna följde efter henne med pukor och dans.
Och Mirjam sjöng för dem: »Sjungen till HERRENS ära, ty högt är han upphöjd.
Häst och man störtade han i havet.»
Därefter lät Mose israeliterna bryta upp från Röda havet, och de drogo ut i öknen Sur; och tre dagar vandrade de i öknen utan att finna vatten.
Så kommo de till Mara; men de kunde icke dricka vattnet i Mara, ty det var bittert.
Därav fick stället namnet Mara.
Då knorrade folket emot Mose och sade: »Vad skola vi dricka?»
Men han ropade till HERREN; och HERREN visade honom ett visst slags trä, som han kastade i vattnet, och så blev vattnet sött.
Där förelade han folket lag och rätt, och där satte han det på prov.
Han sade: »Om du hör HERRENS, din Guds, röst och gör vad rätt är i hans ögon och lyssnar till hans bud och håller alla hans stadgar, så skall jag icke lägga på dig någon av de sjukdomar som jag lade på egyptierna, ty jag är HERREN, din läkare.»
Sedan kommo de till Elim; där funnos tolv vattenkällor och sjuttio palmträd.
Och de lägrade sig där vid vattnet.
Därefter bröt Israels barns hela menighet upp från Elim och kom till öknen Sin, mellan Elim och Sinai, på femtonde dagen i andra månaden efter sitt uttåg ur Egyptens land.
Och Israels barns hela menighet knorrade emot Mose och Aron i öknen;
Israels barn sade till dem: »Ack att vi hade fått dö för HERRENS hand i Egyptens land, där vi sutto vid köttgrytorna och hade mat nog att äta!
Men I haven fört oss hitut i öknen för att låta hela denna hop dö av hunger.»
Då sade HERREN till Mose: »Se, jag vill låta bröd från himmelen regna åt eder.
Och folket skall gå ut och samla för var dag så mycket som behöves.
Så skall jag sätta dem på prov, för att se om de vilja vandra efter min lag eller icke.
Och när de på den sjätte dagen tillreda vad de hava fört hem, skall det vara dubbelt mot vad de eljest för var dag samla in.»
Och Mose och Aron sade till alla Israels barn: »I afton skolen I förnimma att det är HERREN som har fört eder ut ur Egyptens land,
och i morgon skolen I se HERRENS härlighet, HERREN har nämligen hört huru I knorren mot honom.
Ty vad äro vi, att I knorren mot oss?»
Och Mose sade ytterligare: »Detta skall ske därigenom att HERREN i afton giver eder kött att äta, och i morgon bröd att mätta eder med då nu HERREN har hört huru I knorren mot honom.
Ty vad äro vi?
Det är icke mot oss I knorren, utan mot HERREN.»
Och Mose sade till Aron: »Säg till Israels barns hela menighet Träden fram inför HERREN, ty han har hört huru I knorren.»
När sedan Aron talade till Israels barns hela menighet, vände de sig mot öknen, och se, då visade sig HERRENS härlighet i molnskyn.
Och HERREN talade till Mose och sade:
»Jag har hört huru Israels barn knorra.
Tala till dem och säg: Vid aftontiden skolen I få kött att äta och i morgon skolen I få bröd att mätta eder med; så skolen I förnimma att jag är HERREN, eder Gud.»
Och om aftonen kommo vaktlar och övertäckte lägret, och följande morgon låg dagg fallen runt omkring lägret.
Och när daggen som hade fallit gick bort, se, då låg över öknen på jorden något fint, såsom fjäll, något fint, likt rimfrost.
När Israels barn sågo detta, frågade de varandra: »Vad är det?»
Ty de visste icke vad det var.
Men Mose sade till dem: »Detta är brödet som HERREN har givit eder till föda.
Och så har HERREN bjudit: Samlen därav, var och en så mycket han behöver till mat; en gomer på var person skolen I taga, efter antalet av edert husfolk, var och en åt så många som han har i sitt tält.»
Och Israels barn gjorde så, och den ene samlade mer, den andre mindre.
Men när de mätte upp det med gomer-mått, hade den som hade samlat mycket intet till överlopps, och de som hade samlat litet, honom fattades intet; var och en hade så mycket samlat, som han behövde till mat.
Och Mose sade till dem: »Ingen må behålla något kvar härav till i morgon.
Men de lydde icke Mose, utan somliga behöllo något därav kvar till följande morgon.
Då växte maskar däri, och det blev illaluktande.
Och Mose blev förtörnad på dem.
Så samlade de därav var morgon, var och en så mycket han behövde till mat.
Men när solhettan kom smälte det bort.
På den sjätte dagen hade de samlat dubbelt så mycket av brödet, två gomer för var och en.
Och menighetens hövdingar kommo alla och omtalade detta för Mose.
Då sade han till dem: »Detta är efter HERRENS ord; i morgon är sabbatsvila, en HERRENS heliga sabbat.
Baken nu vad I viljen baka, och koken vad I viljen koka, men allt som är till överlopps skolen I ställa i förvar hos eder till i morgon.»
Och de ställde det i förvar till följande morgon, såsom Mose hade bjudit; och nu blev det icke illaluktande, ej heller kom mask däri.
Och Mose sade: »Äten det i dag, ty i dag är HERRENS sabbat; i dag skolen I intet finna på marken.
I sex dagar skolen I samla därav, men på sjunde dagen är sabbat; då skall intet vara att finna.»
Likväl gingo några av folket på den sjunde dagen ut för att samla, men de funno intet.
Då sade HERREN till Mose: »Huru länge viljen I vara motsträviga och icke hålla mina bud och lagar?
Se, HERREN har givit eder sabbaten; därför giver han eder på den sjätte dagen bröd för två dagar.
Så stannen då hemma, var och en hos sig; ingen må gå hemifrån på den sjunde dagen.»
Alltså höll folket sabbat på den sjunde dagen.
Och Israels barn kallade det manna .
Och det liknade korianderfrö, det var vitt, och det smakade såsom semla med honung.
Och Mose sade: »Så har HERREN bjudit: En gomer härav skall förvaras åt edra efterkommande, för att de må se det bröd som jag gav eder att äta i öknen, när jag förde eder ut ur Egyptens land.
Och Mose sade till Aron: »Tag ett kärl och lägg däri en gomer manna, och ställ det inför HERREN till att förvaras åt edra efterkommande.»
Då gjorde man såsom HERREN hade bjudit Mose, och Aron ställde det framför vittnesbördet till att förvaras.
Och Israels barn åto manna i fyrtio år, till dess de kommo till bebott land; de åto manna, till dess de kommo till gränsen av Kanaans land. --
En gomer är tiondedelen av en efa.
Därefter bröt Israels barns hela menighet upp från öknen Sin och tågade från lägerplats till lägerplats, efter HERRENS befallning.
Och de lägrade sig i Refidim; där hade folket intet vatten att dricka.
Då begynte folket tvista med Mose och sade: »Given oss vatten att dricka.»
Mose svarade dem: »Varför tvisten I med mig?
Varför fresten I HERREN?»
Men eftersom folket där törstade efter vatten, knorrade de ytterligare emot Mose och sade: »Varför har du fört oss upp ur Egypten, så att vi, våra barn och vår boskap nu måste dö av törst?»
Då ropade Mose till HERREN och sade: »Vad skall jag göra med detta folk?
Det fattas icke mycket i att de stena mig.»
HERREN svarade Mose: »Gå framför folket, och tag med dig några av de äldste i Israel.
Och tag i din hand staven med vilken du slog Nilfloden, och begiv dig åstad.
Se, jag vill stå där framför dig på Horebs klippa, och du skall slå på klippan, och vatten skall då komma ut ur den, så att folket får dricka.»
Och Mose gjorde så inför de äldste i Israel.
Och han gav stället namnet Massa och Meriba , därför att Israels barn hade tvistat och frestat HERREN och sagt: »Är HERREN ibland oss eller icke?»
Därefter kom Amalek och gav sig i strid med Israel i Refidim.
Då sade Mose till Josua: »Välj ut manskap åt oss, och drag så åstad till strid mot Amalek.
I morgon skall jag ställa mig överst på höjden, med Guds stav i min hand.»
Och Josua gjorde såsom Mose hade tillsagt honom, och gav sig i strid med Amalek.
Men Mose, Aron och Hur stego upp överst på höjden.
Och så länge Mose höll upp sin hand, rådde Israel, men när han lät sin hand sjunka, rådde Amalek.
Och när Moses händer blevo tunga, togo de en sten och lade under honom, och på den satte han sig; sedan stödde Aron och Hur hans händer, en på vardera sidan.
Så höllos hans händer stadiga, till dess solen gick ned.
Och Josua slog Amalek och dess folk med svärdsegg.
Och HERREN sade till Mose: »Teckna upp detta till en åminnelse i en bok, och inprägla det hos Josua, ty jag skall så i grund utplåna minnet av Amalek, att det icke mer skall finnas under himmelen.»
Och Mose byggde ett altare och gav det namnet HERREN mitt baner.
Och han sade: »Ja, jag lyfter min hand upp mot HERRENS tron och betygar att HERREN skall strida mot Amalek från släkte till släkte.»
Och Jetro, prästen i Midjan, Moses svärfader, fick höra allt vad Gud hade gjort med Mose och med sitt folk Israel, huru HERREN hade fört Israel ut ur Egypten.
Då tog Jetro, Moses svärfader, med sig Sippora, Moses hustru, som denne förut hade sänt hem,
så ock hennes två söner -- av dessa hade den ene fått namnet Gersom, »ty», sade Mose, »jag är en främling i ett land som icke är mitt»,
och den andre namnet Elieser, »ty», sade han, »min faders Gud blev mig till hjälp och räddade mig ifrån Faraos svärd». --
Då så Jetro, Moses svärfader, kom med Moses söner och hans hustru till honom i öknen, där han hade slagit upp sitt läger vid Guds berg,
lät han säga till Mose: »Jag, din svärfader Jetro, kommer till dig med din hustru och hennes båda söner.»
Då gick Mose sin svärfader till mötes och bugade sig för honom och kysste honom.
Och när de hade hälsat varandra, gingo de in i tältet.
Och Mose förtäljde för sin svärfader allt vad HERREN hade gjort med Farao och egyptierna, för Israels skull, och alla de vedermödor som de hade haft att utstå på vägen, och huru HERREN hade räddat dem.
Och Jetro fröjdade sig över allt det goda som HERREN hade gjort mot Israel, i det han hade räddat dem ur egyptiernas hand.
Och Jetro sade: »Lovad vare HERREN, som har räddat eder ur egyptiernas hand och ur Faraos hand, HERREN, som har räddat folket undan egyptiernas hand!
Nu vet jag att HERREN är större än alla andra gudar, ty så bevisade han sig, när man handlade övermodigt mot detta folk.»
Och Jetro, Moses svärfader, frambar ett brännoffer och några slaktoffer åt Gud; och Aron och alla de äldste i Israel kommo och höllo måltid med Moses svärfader inför Gud.
Dagen därefter satte Mose sig för att döma folket, och folket stod omkring Mose från morgonen ända till aftonen.
Då nu Moses svärfader såg allt vad han hade att beställa med folket, sade han: »Vad är det allt du har att bestyra med folket?
Varför sitter du här till doms ensam under det att allt folket måste stå omkring dig från morgonen ända till aftonen?»
Mose svarade sin svärfader: »Folket kommer till mig för att fråga Gud.
De komma till mig, när de hava någon rättssak, och jag dömer då mellan dem; och jag kungör då för dem Guds stadgar och lagar.»
Då sade Moses svärfader till honom: »Du går icke till väga på det rätta sättet.
Både du själv och folket omkring dig måsten ju bliva uttröttade; ett sådant förfaringssätt är dig för svårt, du kan icke ensam bestyra detta.
Så lyssna nu till mina ord; jag vill giva dig ett råd, och Gud skall vara med dig.
Du må vara folkets målsman inför Gud och framlägga deras ärenden inför Gud.
Och du må upplysa dem om stadgar och lagar och kungöra dem den väg de skola vandra och vad de skola göra.
Men sök ut åt dig bland allt folket dugande män som frukta Gud, pålitliga män som hata orätt vinning, och sätt dessa till föreståndare för dem, somliga över tusen, andra över hundra, andra över femtio och andra över tio.
Dessa må alltid döma folket.
Kommer något viktigare ärende före, må de hänskjuta det till dig, men alla ringare ärenden må de själva avdöma.
Så skall du göra din börda lättare, därigenom att de bära den med dig.
Om du vill så göra och Gud så bjuder dig, skall du kunna hålla ut; och allt folket här skall då kunna gå hem i frid.»
Och Mose lyssnade till sin svärfaders ord och gjorde allt vad denne hade sagt.
Mose utvalde dugande män ur hela Israel och gjorde dem till huvudmän för folket, till föreståndare somliga över tusen, andra över hundra, andra över femtio och andra över tio.
Dessa skulle alltid döma folket.
Alla svårare ärenden skulle de hänskjuta till Mose, men alla ringare ärenden skulle de själva avdöma.
Därefter lät Mose sin svärfader fara hem, och denne begav sig till sitt land igen.
På den dag då den tredje månaden ingick efter Israels barns uttåg ur Egyptens land kommo de in i Sinais öken.
Ty de bröto upp från Refidim och kommo så till Sinais öken och lägrade sig i öknen; Israel lägrade sig där mitt emot berget.
Och Mose steg upp till Gud; då ropade HERREN till honom uppifrån berget och sade: »Så skall du säga till Jakobs hus, så skall du förkunna för Israels barn:
'I haven själva sett vad jag har gjort med egyptierna, och huru jag har burit eder på örnvingar och fört eder till mig.
Om I nu hören min röst och hållen mitt förbund, så skolen I vara min egendom framför alla andra folk, ty hela jorden är min;
Och I skolen vara mig ett rike av präster och ett heligt folk.'
Detta är vad du skall tala till Israels barn.
När Mose kom tillbaka, sammankallade han de äldste i folket och förelade dem allt detta som HERREN hade bjudit honom.
Då svarade allt folket med en mun och sade: »Allt vad HERREN har talat vilja vi göra.»
Och Mose gick tillbaka till HERREN med folkets svar.
Och HERREN sade till Mose: »Se, jag skall komma till dig i en tjock molnsky, för att folket skall höra, när jag talar med dig, och så tro på dig evärdligen.»
Och Mose framförde folkets svar till HERREN.
Då sade HERREN till Mose: »Gå till folket, och helga dem i dag och i morgon, och I åt dem två sina kläder.
Och må de hålla sig redo till i övermorgon; ty i övermorgon skall HERREN stiga ned på Sinai berg inför allt folkets ögon.
Och du skall märka ut en gräns för folket runt omkring och säga: 'Tagen eder till vara för att stiga upp på berget eller komma vid dess fot.
Var och en som kommer vid berget skall straffas med döden;
men ingen hand må komma vid honom, utan han skall stenas eller skjutas ihjäl.
Evad det är djur eller människa, skall en sådan mista livet.'
När jubelhornet ljuder med utdragen ton, då må de stiga upp på berget.»
Och Mose steg ned från berget till folket och helgade folket, och de tvådde sina kläder.
Och han sade till folket: »Hållen eder redo till i övermorgon; ingen komme vid en kvinna.»
På tredje dagen, när det hade blivit morgon, begynte det dundra och blixtra, och en tung molnsky kom över berget, och ett mycket starkt basunljud hördes; och allt folket i lägret bävade.
Men Mose förde folket ut ur lägret, Gud till mötes; och de ställde sig nedanför berget.
Och hela Sinai berg höljdes i rök, vid det att HERREN kom ned därpå i eld; och en rök steg upp därifrån, lik röken från en smältugn, och hela berget bävade storligen.
Och basunljudet blev allt starkare och starkare.
Mose talade, och Gud svarade honom med hög röst.
Och HERREN steg ned på Sinai berg, på toppen av berget, och HERREN kallade Mose upp till bergets topp; då steg Mose ditupp.
Och HERREN sade till Mose: »Stig ned och varna folket, så att de icke tränga sig fram för att se HERREN, ty då skola många av dem falla.
Jämväl prästerna, som få nalkas HERREN, skola helga sig, för att HERREN icke må låta dem drabbas av fördärv.»
Men Mose svarade HERREN: »Folket kan icke stiga upp på Sinai berg, ty du har själv varnat oss och sagt att jag skulle märka ut en gräns omkring berget och helga det.»
Då sade HERREN till honom: »Gå ditned, och kom sedan åter upp och hav Aron med dig.
Men prästerna och folket må icke tränga sig fram för att stiga upp till HERREN på det att han icke må låta dem drabbas av fördärv.»
Och Mose steg ned till folket och sade dem detta.
Och Gud talade alla dessa ord och sade:
Jag är HERREN, din Gud, som har fört dig ut ur Egyptens land, ur träldomshuset.
Du skall inga andra gudar hava jämte mig.
Du skall icke göra dig något beläte eller någon bild, vare sig av det som är uppe i himmelen, eller av det som är nere på jorden, eller av det som är i vattnet under jorden.
Du skall icke tillbedja sådana, ej heller tjäna dem; ty jag, HERREN, din Gud, är en nitälskande Gud, som hemsöker fädernas missgärning på barn och efterkommande i tredje och fjärde led, när man hatar mig,
men som gör nåd med tusenden, när man älskar mig och håller mina bud.
Du skall icke missbruka HERRENS, din Guds, namn, ty HERREN skall icke låta den bliva ostraffad, som missbrukar hans namn.
Tänk på sabbatsdagen, så att du helgar den.
Sex dagar skall du arbeta och förrätta alla dina sysslor;
men den sjunde dagen är HERRENS, din Guds, sabbat; då skall du ingen syssla förrätta, ej heller din son eller din dotter, ej heller din tjänare eller din tjänarinna eller din dragare, ej heller främlingen som är hos dig inom dina portar.
Ty på sex dagar gjorde HERREN himmelen och jorden och havet och allt vad i dem är, men han vilade på sjunde dagen; därför har HERREN välsignat sabbatsdagen och helgat den.
Hedra din fader och din moder, för att du må länge leva i det land som HERREN, din Gud, vill giva dig.
Du skall icke dräpa.
Du skall icke begå äktenskapsbrott.
Du skall icke stjäla.
Du skall icke bära falskt vittnesbörd mot din nästa.
Du skall icke hava begärelse till din nästas hus.
Du skall icke hava begärelse till din nästas hustru, ej heller till hans tjänare eller hans tjänarinna, ej heller till hans oxe eller hans åsna, ej heller till något annat som tillhör din nästa.
Och allt folket förnam dundret och eldslågorna och basunljudet och röken från berget; och när folket förnam detta, bävade de och höllo sig på avstånd.
Och de sade till Mose: »Tala du till oss, så vilja vi höra, men låt icke Gud tala till oss, på det att vi icke må dö.»
Men Mose sade till folket: »Frukten icke, ty Gud har kommit för att sätta eder på prov, och för att I skolen hava hans fruktan för ögonen, så att I icke synden.»
Alltså höll folket sig på avstånd, under det att Mose gick närmare till töcknet i vilket Gud var.
Och HERREN sade till Mose: Så skall du säga till Israels barn: I haven själva förnummit att jag har talat till eder från himmelen.
I skolen icke göra eder gudar jämte mig; gudar av silver eller guld skolen I icke göra åt eder.
Ett altare av jord skall du göra åt mig och offra därpå dina brännoffer och tackoffer, din småboskap och dina fäkreatur.
Överallt på den plats där jag stiftar en åminnelse åt mitt namn skall jag komma till dig och välsigna dig.
Men om du vill göra åt mig ett altare av stenar, så må du icke bygga det av huggen sten; ty om du kommer vid stenen med din mejsel, så oskärar du den.
Icke heller må du stiga upp till mitt altare på trappor, på det att icke din blygd må blottas därinvid.
Dessa äro de rätter som du skall förelägga dem:
Om du köper en hebreisk träl, skall han tjäna i sex år, men på det sjunde skall han givas fri, utan lösen.
Har han kommit allena, så skall han givas fri allena; var han gift, så skall hans hustru givas fri med honom.
Har hans herre givit honom en hustru, och har denna fött honom söner eller döttrar, så skola hustrun och hennes barn tillhöra hennes herre, och allenast mannen skall givas fri.
Men om trälen säger: »Jag har min herre, min hustru och mina barn så kära, att jag icke vill givas fri»,
då skall hans herre föra honom fram för Gud och ställa honom vid dörren eller dörrposten, och hans herre skall genomborra hans öra med en syl; därefter vare han hans träl evärdligen.
Om någon säljer sin dotter till trälinna, så skall hon icke givas fri såsom trälarna givas fria.
Misshagar hon sin herre, sedan denne förut har ingått förbindelse med henne, så låte han henne köpas fri.
Till främmande folk have han icke makt att sälja henne, när han så har handlat trolöst mot henne.
Men om han låter sin son ingå förbindelse med henne, så förunne han henne döttrars rätt.
Tager han sig ännu en hustru, så göre han icke någon minskning i den förras kost, beklädnad eller äktenskapsrätt.
Om han icke låter henne njuta sin rätt i dessa tre stycken, så skall hon givas fri, utan lösen och betalning.
Den som slår någon, så att han dör, han skall straffas med döden.
Men om han icke traktade efter den andres liv, utan Gud lät denne oförvarandes träffas av hans hand, så skall jag anvisa dig en ort dit han kan fly.
Men om någon begår det dådet att han dräper sin nästa med list, så skall du gripa honom, vore han ock invid mitt altare, och han måste dö.
Den som slår sin fader eller sin moder, han skall straffas med döden.
Den som stjäl en människa, vare sig han sedan säljer den stulne, eller denne finnes kvar hos honom, han skall straffas med döden.
Den som uttalar förbannelser över sin fader eller sin moder, han skall straffas med döden.
Om män tvista med varandra, och den ene slår den andre med en sten eller med knuten hand, så att denne väl icke dör, men bliver sängliggande,
dock att han sedan kommer sig och kan gå ute, stödd vid sin stav, så skall den som slog honom vara fri ifrån straff; allenast ersätte han honom för den tid han har förlorat och besörje sjukvård åt honom.
Om någon slår sin träl eller sin trälinna med en käpp, så att den slagne dör under hans hand, så skall han straffas därför.
Men om den slagne lever en eller två dagar, skall han icke straffas, ty det var hans egna penningar.
Om män träta med varandra, och någon av dem stöter till en havande kvinna, så att hon föder fram sitt foster, men eljest ingen olycka sker, så böte han vad kvinnans man ålägger honom och betale efter skiljedomares prövning.
Men om olycka sker, skall liv givas för liv,
öga för öga, tand för tand, hand för hand, fot för fot,
brännskada för brännskada, sår för sår, blånad för blånad.
Om någon slår sin träl eller sin trälinna i ögat och fördärvar det, så släppe han den skadade fri, till ersättning för ögat.
Sammalunda, om någon slår ut en tand på sin träl eller sin trälinna, så släppe han den skadade fri, till ersättning för tanden.
Om en oxe stångar någon till döds, man eller kvinna, så skall oxen stenas, och köttet må icke ätas; men oxens ägare vara fri ifrån straff.
Men om oxen förut har haft vanan att stångas, och hans ägare har blivit varnad, men denne ändå icke tager vara på honom, och oxen så dödar någon, man eller kvinna, då skall oxen stenas, och hans ägare skall ock dödas.
Men skulle lösepenning bliva denne ålagd, så give han till lösen för sitt liv så mycket som ålägges honom.
Är det en gosse eller en flicka som har blivit stångad av oxen, så skall med denne förfaras efter samma lag.
Men om oxen stångar en träl eller en trälinna, så skall ägaren giva åt den stångades herre trettio siklar silver, och oxen skall stenas.
Om någon öppnar en brunn, eller om någon gräver en ny brunn och icke täcker över den, och sedan en oxe eller en åsna faller däri,
så skall brunnens ägare giva ersättning i penningar åt djurets ägare, men den döda kroppen skall vara hans.
Om någons oxe stångar en annans oxe, så att denne dör, så skola de sälja den levande oxen och dela betalningen för honom och därjämte dela den döda kroppen.
Var det däremot känt att oxen förut hade vanan att stångas, men tog hans ägare ändå icke vara på honom, så skall han ersätta oxe med oxe, men den döda kroppen skall vara hans.
Om någon stjäl en oxe eller ett får och slaktar eller säljer djuret, så skall han giva fem oxar i ersättning för oxen, och fyra får för fåret.
Ertappas tjuven vid inbrottet och bliver slagen till döds, så vilar ingen blodskuld på dråparen.
Men hade solen gått upp, när de skedde, då är det blodskuld.
Tjuven skall giva full ersättning; äger han intet, så skall han säljas, till gäldande av vad han har stulit.
Om det stulna djuret, det må vara oxe eller åsna eller får, påträffas levande i hans våld, skall han giva dubbel ersättning.
Om någon låter avbeta en åker eller vingård, eller släpper sin boskap lös, så att denna betar på en annans åker, då skall han ersätta skadan med det bästa från sin åker och med det bästa från sin vingård.
Om eld kommer lös och fattar i törnhäckar, och därvid sädesskylar bliva uppbrända eller oskuren säd eller annat på åkern, så skall den som har vållat branden giva full ersättning.
Om någon giver åt en annan penningar eller gods att förvara, och detta bliver stulet ur hans hus, så skall tjuven, om han ertappas, giva dubbel ersättning.
Ertappas icke tjuven, då skall man föra husets ägare fram för Gud, på det att det må utrönas om han icke har förgripit sig på sin nästas tillhörighet.
Om fråga uppstår angående orättrådigt tillgrepp -- det må gälla oxe eller åsna eller får eller kläder eller något annat som har förlorats -- och någon påstår att en orättrådighet verkligen har ägt rum, så skall båda parternas sak komma inför Gud.
Den som Gud dömer skyldig, han skall ersätta den andre dubbelt.
Om någon giver åt en annan i förvar en åsna eller en oxe eller ett får, eller vilket annat husdjur det vara må, och detta dör eller bliver skadat eller bortrövat, utan att någon ser det,
Så skall det dem emellan komma till en ed vid HERREN, för att det må utrönas om den ene icke har förgripit sig på den andres tillhörighet; denna ed skall ägaren antaga och den andre behöver icke giva någon ersättning.
Men om det har blivit bortstulet från honom, då skall han ersätta ägaren därför.
Har det blivit ihjälrivet, skall han föra fram det ihjälrivna djuret såsom bevis; han behöver då icke giva ersättning därför.
Om någon lånar ett djur av en annan, och detta bliver skadat eller dör, och dess ägare därvid icke är tillstädes, så skall han giva full ersättning.
Är dess ägare tillstädes, då behöver han icke giva ersättning.
Var djuret lejt, då är legan ersättning.
Om någon förför en jungfru som icke är trolovad och lägrar henne, så skall han giva brudgåva för henne och taga henne till hustru.
Vägrar hennes fader att giva henne åt honom, då skall han gälda en så stor penningsumma som man plägar giva i brudgåva för en jungfru.
En trollkvinna skall du icke låta leva.
Var och en som beblandar sig med något djur skall straffas med döden.
Den som offrar åt andra gudar än åt HERREN allena, han skall givas till spillo.
En främling skall du icke förorätta eller förtrycka; I haven ju själva varit främlingar i Egyptens land.
Änkor och faderlösa skolen I icke behandla illa.
Behandlar du dem illa, så skall jag förvisso höra deras rop, när de ropa till mig;
och min vrede skall upptändas, och jag skall dräpa eder med svärd; så att edra egna hustrur bliva änkor och edra barn faderlösa.
Lånar du penningar åt någon fattig hos dig bland mitt folk, så skall du icke handla mot honom såsom en ockrare; I skolen icke pålägga honom någon ränta.
Har du av din nästa tagit hans mantel i pant, så skall du giva den tillbaka åt honom, innan solen går ned;
den är ju det enda täcke han har, och med den skyler han sin kropp.
Vad skall han eljest hava på sig, när han ligger och sover?
Om han måste ropa till mig, så skall jag höra, ty jag är barmhärtig.
Gud skall du icke häda, och över en hövding i ditt folk skall du icke uttala förbannelser.
Av det som fyller din lada och av det som flyter ifrån din press skall du utan dröjsmål frambära din gåva.
Den förstfödde bland dina söner skall du giva åt mig.
På samma sätt skall du göra med dina fäkreatur och din småboskap.
I sju dagar skola de stanna hos sina mödrar; på åttonde dagen skall du giva dem åt mig.
Och I skolen vara mig ett heligt: folk; kött av ett djur som har blivit ihjälrivet på marken skolen I icke äta, åt hundarna skolen I kasta det.
Du skall icke utsprida falskt rykte; åt den som har en orätt sak skall du icke giva ditt bistånd genom att bliva ett orättfärdigt vittne.
Du skall icke följa med hopen i vad ont är, eller vittna så i någon sak, att du böjer dig efter hopen och vränger rätten.
Du skall icke vara partisk för den ringe i någon hans sak.
Om du träffar på din fiendes oxe eller åsna som har kommit vilse, så skall du föra djuret tillbaka till honom.
Om du ser din oväns åsna ligga dignad under sin börda, så skall du ingalunda lämna mannen ohulpen, utan hjälpa honom att lösa av bördan.
Du skall icke i någon sak vränga rätten för den fattige som du har hos dig.
Du skall hålla dig fjärran ifrån orätt sak; du skall icke dräpa den som är oskyldig och har rätt, ty jag skall icke giva rätt åt någon som är skyldig.
Du skall icke taga mutor, ty mutor förblinda de seende och förvrida de rättfärdigas sak.
En främling skall du icke förtrycka; I veten ju huru främlingen känner det, eftersom I själva haven varit främlingar i Egyptens land.
I sex år skall du beså din jord och inbärga dess gröda;
men under det sjunde året skall du låta den vila och ligga orörd, för att de fattiga bland ditt folk må äta därav; vad de lämna kvar, det må ätas av markens djur.
Så skall du ock göra med din vingård och med din olivplantering.
Sex dagar skall du göra ditt arbete, men på sjunde dagen skall du hålla vilodag, för att din oxe och din åsna må hava ro, och din tjänstekvinnas son och främlingen må njuta vila.
I alla de stycken om vilka jag har talat till eder skolen I taga eder till vara.
Och andra gudars namn skolen I icke nämna; de skola icke höras i din mun.
Tre gånger om året skall du hålla högtid åt mig.
Det osyrade brödets högtid skall du hålla: i sju dagar skall du äta osyrat bröd, såsom jag har bjudit dig, på den bestämda tiden i månaden Abib, eftersom du då drog ut ur Egypten; men med tomma händer skall ingen träda fram inför mitt ansikte.
Du skall ock hålla skördehögtiden, när du skördar förstlingen av ditt arbete, av det du har sått på marken.
Bärgningshögtiden skall du ock hålla, vid årets utgång, när du inbärgar frukten av ditt arbete från marken.
Tre gånger om året skall allt ditt mankön träda fram inför HERRENS, din Herres, ansikte.
Du skall icke offra blodet av mitt slaktoffer jämte något som är syrat.
Och det feta av mitt högtidsoffer skall icke lämnas kvar över natten till morgonen.
Det första av din marks förstlingsfrukter skall du föra till HERRENS, din Guds, hus.
Du skall icke koka en killing i dess moders mjölk.
Se, jag skall sända en ängel framför dig, som skall bevara dig på vägen och föra dig till den plats som jag har utsett.
Tag dig till vara inför honom och hör hans röst, var icke gensträvig mot honom, han skall icke hava fördrag med edra överträdelser, ty mitt namn är i honom.
Men om du hör hans röst och gör allt vad jag säger, så skall jag bliva en fiende till dina fiender och en ovän till dina ovänner.
Ty min ängel skall gå framför dig och skall föra dig till amoréernas, hetiternas, perisséernas, kananéernas, hivéernas och jebuséernas land, och jag skall utrota dem.
Du må icke tillbedja deras gudar eller tjäna dem eller göra såsom man där gör, utan du skall slå dem ned i grund och bryta sönder deras stoder.
Men HERREN, eder Gud, skolen I tjäna, så skall han för dig välsigna både mat och dryck; sjukdom skall jag då ock avvända från dig.
I ditt land skall då icke finnas någon kvinna som föder i otid eller är ofruktsam.
Dina dagars mått skall jag göra fullt.
Förskräckelse för mig skall jag sända framför dig och vålla förvirring bland alla de folk som du kommer till, och jag skall driva alla dina fiender på flykten för dig.
Jag skall sända getingar framför dig, och de skola förjaga hivéerna, kananéerna och hetiterna undan för dig.
Dock skall jag icke på ett och samma år förjaga dem för dig, på det att icke landet så må bliva en ödemark och vilddjuren föröka sig till din skada;
utan småningom skall jag förjaga dem för dig, till dess du har förökat dig, så att du kan taga landet till din arvedel.
Och jag skall låta ditt lands gränser gå från Röda havet till filistéernas hav, och från öknen till floden; ty jag skall giva landets inbyggare i eder hand, och du skall förjaga dem, så att de fly för dig.
Du må icke sluta förbund med dem eller deras gudar.
De skola icke få bo kvar i ditt land, på det att de icke må förleda dig till synd mot mig; ty du kunde ju komma att tjäna deras gudar, och detta skulle bliva dig till en snara.
Och han sade till Mose: »Stig upp till HERREN, du själv jämte Aron, Nadab och Abihu och sjuttio av de äldste i Israel; och I skolen tillbedja på avstånd.
Mose allena må träda fram till HERREN, de andra må icke träda fram; ej heller må folket stiga ditupp med honom.»
Och Mose kom till folket och förkunnade för det alla HERRENS ord och alla hans rätter.
Då svarade allt folket med en mun och sade: »Efter alla de ord HERREN har talat vilja vi göra.»
Därefter upptecknade Mose alla HERRENS ord.
Och följande morgon stod han bittida upp och byggde ett altare nedanför berget.
Och han reste där tolv stoder, efter Israels tolv stammar.
Och han sände israeliternas unga män åstad till att offra brännoffer, så ock slaktoffer av tjurar till tackoffer åt HERREN.
Och Mose tog hälften av blodet och slog det i skålarna, och den andra hälften av blodet stänkte han på altaret.
Och han tog förbundsboken och, föreläste den för folket.
Och de sade: »Allt vad HERREN har sagt vilja vi göra och lyda.
Då tog Mose blodet och stänkte därav på folket och sade: »Se, detta är förbundets blod, det förbunds som HERREN har slutit med eder, i enlighet med alla dessa ord.»
Och Mose och Aron, Nadab och Abihu och sjuttio av de äldste i Israel stego ditupp.
Och de fingo se Israels Gud; och under hans fötter var likasom ett inlagt golv av safirer, likt själva himmelen i klarhet.
Men han lät icke sin hand drabba Israels barns ypperste, utan sedan de hade skådat Gud, åto de och drucko.
Och HERREN sade till Mose: »Stig upp till mig på berget och bliv kvar där, så skall jag giva dig stentavlorna och lagen och budorden som jag har skrivit, till undervisning för dessa.»
Då begav sig Mose åstad med sin tjänare Josua; och Mose steg upp på Guds berg.
Men till de äldste sade han: »Vänten här på oss, till dess att vi komma tillbaka till eder.
Se, Aron och Hur äro hos eder; den som har något att andraga, han må vända sig till dem.»
Så steg Mose upp på berget, och molnskyn övertäckte berget.
Och HERRENS härlighet vilade på Sinai berg, och molnskyn övertäckte det i sex dagar; men den sjunde dagen kallade han på Mose ur skyn.
Och HERRENS härlighet tedde sig inför Israels barns ögon såsom en förtärande eld, på toppen av berget.
Och Mose gick mitt in i skyn och steg upp på berget.
Sedan blev Mose kvar på berget i fyrtio dagar och fyrtio nätter.
Och HERREN talade till Mose och sade:
Säg till Israels barn att de upptaga en gärd åt mig; av var och en som har ett därtill villigt hjärta skolen I upptaga denna gärd åt mig.
Och detta är vad I skolen upptaga av dem såsom gärd: guld, silver och koppar
mörkblått, purpurrött, rosenrött och vitt garn och gethår,
rödfärgade vädurskinn, tahasskinn, akacieträ,
olja till ljusstaken, kryddor till smörjelseoljan och till den välluktande rökelsen,
äntligen onyxstenar och infattningsstenar, till att användas för efoden och för bröstskölden.
Och de skola göra åt mig en helgedom, för att jag må bo mitt ibland dem.
Tabernaklet och alla dess tillbehör skolen I göra alldeles efter de mönsterbilder som jag visar dig.
De skola göra en ark av akacieträ, två och en halv aln lång, en och en halv aln bred och en och en halv aln hög.
Och du skall överdraga den med rent guld, innan och utan skall du överdraga den; och du skall på den göra en rand av guld runt omkring.
Och du skall till den gjuta fyra ringar av guld och sätta dem över de fyra fötterna, två ringar på ena sidan och två ringar på andra sidan.
Och du skall göra stänger av akacieträ och överdraga dem med guld.
Och stängerna skall du skjuta in i ringarna, på sidorna av arken, så att man med dem kan bära arken.
Stängerna skola sitta kvar i ringarna på arken; de få icke dragas ut ur dem.
Och i arken skall du lägga vittnesbördet, som jag skall giva dig.
Och du skall göra en nådastol av rent guld, två och en halv aln lång och en och en halv aln bred.
Och du skall göra två keruber av guld; i drivet arbete skall du göra dem och sätta dem vid de båda ändarna av nådastolen.
Du skall göra en kerub till att sätta vid ena ändan, och en kerub till att sätta vid andra ändan.
I ett stycke med nådastolen skolen I göra keruberna vid dess båda ändar.
Och keruberna skola breda ut sina vingar och hålla dem uppåt, så att de övertäcka nådastolen med sina vingar, under det att de hava sina ansikten vända mot varandra; ned mot nådastolen skola keruberna vända sina ansikten.
Och du skall sätta nådastolen ovanpå arken, och i arken skall du lägga vittnesbördet, som jag skall giva dig.
Och där skall jag uppenbara mig för dig; från nådastolen, från platsen mellan de två keruberna, som stå på vittnesbördets ark, skall jag tala med dig om alla bud som jag genom dig vill giva Israels barn.
Du skall ock göra ett bord av akacieträ, två alnar långt, en aln brett och en och en halv aln högt.
Och du skall överdraga det med rent guld; och du skall göra en rand av guld därpå runt omkring
Och runt omkring det skall du göra en list av en hands bredd, och runt omkring listen skall du göra en rand av guld.
Och du skall till bordet göra fyra ringar av guld och sätta ringarna i de fyra hörnen vid de fyra fötterna.
Invid listen skola ringarna sitta, för att stänger må skjutas in i dem, så att man kan bära bordet.
Och du skall göra stängerna av akacieträ och överdraga dem med guld, och med dem skall bordet bäras.
Du skall ock göra därtill fat och skålar, kannor och bägare, med vilka man skall utgjuta drickoffer; av rent guld skall du göra dem.
Och du skall beständigt hava skådebröd liggande på bordet inför mitt ansikte.
Du skall ock göra en ljusstake av rent guld.
I drivet arbete skall ljusstaken göras, med sin fotställning och sitt mittelrör; kalkarna därpå, kulor och blommor skola vara i ett stycke med den.
Och sex armar skola utgå från ljusstakens sidor, tre armar från ena sidan och tre armar från andra sidan.
På den ena armen skola vara tre kalkar, liknande mandelblommor, vardera bestående av en kula och en blomma, och på den andra armen sammalunda tre kalkar, liknande mandelblommor, vardera bestående av en kula och en blomma så skall det vara på de sex arma som utgå från ljusstaken.
Men på själva ljusstaken skola vara fyra kalkar, liknande mandelblommor, med sina kulor och blommor.
En kula skall sättas under del första armparet som utgår från ljusstaken, i ett stycke med den, och en kula under det andra armparet som utgår från ljusstaken, i ett stycke med den, och en kula under det tredje armparet som utgår från ljusstaken, i ett stycke med den: alltså under de sex armar som utgå från ljusstaken.
Deras kulor och armar skola vara: i ett stycke med den, alltsammans ett enda stycke i drivet arbete av rent guld.
Och du skall till den göra sju lampor, och lamporna skall man sätta upp så, att den kastar sitt sken över platsen därframför.
Och lamptänger och brickor till den skall du göra av rent guld.
Av en talent rent guld skall man göra den med alla dessa tillbehör.
Och se till, att du gör detta efter de mönsterbilder som hava blivit dig visade på berget.
Tabernaklet skall du göra av tio tygvåder; av tvinnat vitt garn och av mörkblått, purpurrött och rosenrött garn skall du göra dem, med keruber på, i konstvävnad.
Var våd skall vara tjuguåtta alnar lång och fyra alnar bred; alla våderna skola hava samma mått.
Fem av våderna skola fogas tillhopa med varandra; likaså skola de fem övriga våderna fogas tillhopa med varandra.
Och du skall sätta öglor av mörkblått garn i kanten på den ena våden, ytterst på det hopfogade stycket; så skall du ock göra i kanten på den våd som sitter ytterst i det andra hopfogade stycket.
Femtio öglor skall du sätta på den ena våden, och femtio öglor skall du sätta ytterst på motsvarande våd i det andra hopfogade stycket, så att öglorna svara emot varandra.
Och du skall göra femtio häktor av guld och foga tillhopa våderna med varandra medelst häktorna, så att tabernaklet utgör ett helt.
Du skall ock göra tygvåder av gethår till ett täckelse över tabernaklet; elva sådana våder skall du göra.
Var vad skall vara trettio alnar lång och fyra alnar bred; de elva våderna skola hava samma mått.
Fem av våderna skall du foga tillhopa till ett särskilt stycke, och likaledes de sex övriga våderna till ett särskilt stycke, och den sjätte våden skall du lägga dubbel på framsidan av tältet.
Och du skall satta femtio öglor i kanten på den ena våden, den som sitter ytterst i det ena hopfogade stycket, och femtio öglor i kanten på motsvarande våd i det andra hopfogade stycket.
Och du skall göra femtio häktor av koppar och haka in häktorna i öglorna och foga täckelset tillhopa, så att det utgör ett helt.
Men vad överskottet av täckelsets våder angår, det som räcker över, så skall den halva våd som räcker över hänga ned på baksidan av tabernaklet.
Och den aln på vardera sidan, som på längden av täckelsets våder räcker över, skall hänga ned på båda sidorna av tabernaklet för att övertäcka det.
Vidare skall du göra ett överdrag av rödfärgade vädurskinn till täckelset, och ytterligare ett överdrag av tahasskinn att lägga ovanpå detta.
Bräderna till tabernaklet skall du göra av akacieträ, och de skola ställas upprätt.
Tio alnar långt och en och en halv aln brett skall vart bräde vara.
Vart bräde skall hava två tappar, förbundna sinsemellan med en list; så skall du göra på alla bräderna till tabernaklet.
Och av tabernaklets bräder skall du sätta tjugu på södra sidan, söderut.
Och du skall göra fyrtio fotstycken av silver att sätta under de tjugu bräderna, två fotstycken under vart bräde för dess två tappar.
Likaledes skall du på tabernaklets andra sida, den norra sidan, sätta tjugu bräder,
med deras fyrtio fotstycken av silver, två fotstycken under vart bräde.
Men på baksidan av tabernaklet, västerut, skall du sätta sex bräder.
Och två bräder skall du sätta på tabernaklets hörn, på baksidan;
och vartdera av dessa skall vara sammanfogat av två nedtill, och likaledes sammanhängande upptill, till den första ringen.
Så skall det vara med dem båda.
Dessa skola sättas i de båda hörnen.
Således bliver det åtta bräder med tillhörande fotstycken av silver, sexton fotstycken, nämligen två fotstycken under vart bräde.
Och du skall göra tvärstänger av akacieträ, fem till de bräder som äro på tabernaklets ena sida
och fem tvärstänger till de bräder som äro på tabernaklets andra sida, och fem tvärstänger till de bräder som äro på tabernaklets baksida, västerut.
Och den mellersta tvärstången, den som sitter mitt på bräderna, skall gå tvärs över, från den ena ändan till den andra.
Och bräderna skall du överdraga med guld, och ringarna på dem, i vilka tvärstängerna skola skjutas in, skall du göra av guld, och tvärstängerna skall du överdraga med guld.
Och du skall sätta upp tabernaklet, sådant det skall vara, såsom det har blivit dig visat på berget.
Du skall ock göra en förlåt av mörkblått, purpurrött, rosenrött och tvinnat vitt garn; den skall göras i konstvävnad, med keruber på.
Och du skall hänga upp den på fyra stolpar av akacieträ, som skola vara överdragna med guld och hava bakar av guld och stå på fyra fotstycken av silver.
Och du skall hänga upp förlåten under häktorna, och föra dit vittnesbördets ark och ställa den innanför förlåten; och så skall förlåten för eder vara en skiljevägg mellan det heliga och det allraheligaste.
Och du skall sätta nådastolen på vittnesbördets ark inne i det allraheligaste.
Men bordet skall du ställa utanför förlåten, och ljusstaken mitt emot bordet, på tabernaklets södra sida; bordet skall du alltså ställa på norra sidan.
Och du skall göra ett förhänge för ingången till tältet, i brokig vävnad av mörkblått, purpurrött, rosenrött och tvinnat vitt garn.
Och du skall till förhänget göra fem stolpar av akacieträ och överdraga dem med guld, och hakarna på dem skola vara av guld, och du skall till dem gjuta fem fotstycken av koppar.
Du skall ock göra ett altare av akacieträ, fem alnar långt och fem alnar brett -- så att altaret bildar en liksidig fyrkant -- och tre alnar högt.
Och du skall göra hörn därtill, Som skola sitta i dess fyra hörn; i ett stycke därmed skola hörnen vara.
Och du skall överdraga det med koppar.
Och kärl till att föra bort askan skall du göra därtill, så ock skovlar, skålar, gafflar och fyrfat.
Alla dess tillbehör skall du göra av koppar.
Och du skall göra ett galler därtill, ett nätverk av koppar, och på nätet skall du sätta fyra ringar av koppar i dess fyra hörn.
Och du skall sätta det under avsatsen på altaret, nedtill, så att nätet räcker upp till mitten av altaret.
Och du skall göra stänger till altaret, stänger av akacieträ, och överdraga dem med koppar.
Och stängerna skola skjutas in i ringarna, så att stängerna sitta på altarets båda sidor, när man bär det.
Ihåligt skall du göra det, av plankor.
Såsom det har blivit dig visat på berget, så skall det göras.
Du skall ock göra en förgård till tabernaklet.
För den södra sidan, söderut, skola omhängen till förgården göras av tvinnat vitt garn, hundra alnar långa -- detta för den ena sidan;
Och stolparna till dem skola vara tjugu och dessas fotstycken tjugu, av koppar, men stolparnas hakar och kransar skola vara av silver.
Likaledes skola för norra långsidan omhängen göras, hundra alnar långa; och stolparna till dem skola vara tjugu och dessas fotstycken tjugu, av koppar, men stolparnas hakar och kransar skola vara av silver.
Och förgårdens västra kortsida skall hava omhängen som äro femtio alnar långa; stolparna till dem skola vara tio och dessas fotstycken tio.
Och förgårdens bredd på fram sidan, österut, skall vara femtio alnar
Och omhängena skola vara femton alnar långa på ena sidan därav, med tre stolpar på tre fotstycken;
likaledes skola omhängena på andra sidan vara femton alnar långa med tre stolpar på tre fotstycken.
Och till förgårdens port skall göras ett förhänge, tjugu alnar långt i brokig vävnad av mörkblått, purpurrött, rosenrött och tvinnat vitt garn, med fyra stolpar på fyra fotstycken.
Alla stolparna runt omkring för gården skola vara försedda med kransar av silver och hava hakar av silver; men deras fotstycken skola vara av koppar.
Förgården skall vara hundra alnar lång och femtio alnar bred utefter hela längden; omhägnaden skall vara fem alnar hög, av tvinnat vitt garn; och fotstyckena skola vara av koppar.
Alla tabernaklets tillbehör för allt arbete därvid, så ock alla dess pluggar och alla förgårdens pluggar skola vara av koppar.
Och du skall bjuda Israels barn att bära till dig ren olja, av stötta oliver, till ljusstaken, så att lamporna dagligen kunna sättas upp.
I uppenbarelsetältet, utanför den förlåt som hänger framför vittnesbördet, skola Aron och hans söner sköta den, från aftonen till morgonen, inför HERRENS ansikte.
Detta skall vara en evärdlig stadga från släkte till släkte, en gärd av Israels barn.
Och du skall låta din broder Aron och hans söner med honom, träd fram till dig ur Israels barns krets för att de må bliva plåster åt mig Aron själv och hans söner: Nadab och Abihu, Eleasar och Itamar.
Och du skall göra åt din broder Aron heliga kläder, till ära och prydnad.
Och du skall tillsäga alla edra konstförfarna män, som jag har uppfyllt med vishetens ande, att de skola göra kläder åt Aron, för att har må helgas till att bliva präst åt mig.
Och dessa äro de kläder som de skola göra: bröstsköld, efod, kåpa, rutig livklädnad, huvudbindel och bälte.
De skola göra heliga kläder åt din broder Aron och hans söner, för att han må bliva präst åt mig.
Och härtill skola de taga av guldet och av det mörkblåa, det purpurröda, det rosenröda och det vita garnet.
Efoden skola de göra av guld och av mörkblått purpurrött, rosenrött och tvinnat vitt garn, i konstvävnad.
Den skall vid sina båda ändar hava två axelstycken, som skola fästas ihop, så att den hållen hopfäst.
Och skärpet, som skall sitta på efoden och sammanhålla den, skall vara av samma slags vävnad och i ett stycke med den: av guld och av mörkblått, purpurrött, rosenrött och tvinnat vitt garn.
Och du skall taga två onyxstenar och på dem inrista Israels söners namn,
sex av namnen på den ena stenen och de sex övrigas namn på den andra stenen, efter ättföljd.
Med stensnidarkonst, såsom man graverar signetringar, skall du inrista Israels söners namn på de två stenarna.
Med nätverk av guld skall du omgiva dessa.
Och du skall satta de båda stenarna på efodens axelstycken, för att stenarna må bringa Israels barn i åminnelse; Aron skall bära deras namn inför HERRENS ansikte på sina båda axlar, för att bringa dem i åminnelse.
Och du skall göra flätverk av guld,
så ock två kedjor av rent guld; i virat arbete skall du göra dessa, såsom man gör snodder.
Och du skall fästa de snodda kedjorna vid flätverken.
En domssköld skall du göra i konstvävnad; du skall göra den i samma slags vävnad som efoden: av guld och av mörkblått, purpurrött, rosenrött och tvinnat vitt garn skall du göra den.
Den skall vara liksidigt fyrkantig och hava form av en väska, ett kvarter lång och ett kvarter bred.
Och du skall besätta den med infattade stenar, ordnade på fyra rader: i första raden en karneol, en topas och en smaragd;
i andra raden en karbunkel, en safir och en kalcedon;
i tredje raden en hyacint, en agat och en ametist;
i fjärde raden en krysolit, en onyx och en jaspis.
Omgivna med flätverk av guld skola de sitta i sin infattning.
Stenarna skola vara tolv, efter Israels söners namn, en för vart namn; var sten skall bära namnet på en av de tolv stammarna, inristat på samma sätt som man graverar signetringar.
Och du skall till bröstskölden göra kedjor i virat arbete, såsom man gör snodder, av rent guld.
Vidare skall du till bröstskölden göra två ringar av guld och sätta dessa båda ringar i två av bröstsköldens hörn.
Och du skall fästa de båda guldsnodderna vid de båda ringarna, i bröstsköldens hörn.
Och de två snoddernas båda andra ändar skall du fästa vid de två flätverken och så fästa dem vid efodens axelstycken på dess framsida.
Och du skall göra två andra ringar av guld och sätta dem i bröstsköldens båda andra hörn, vid den kant därpå, som är vänd inåt mot efoden.
Och ytterligare skall du göra två ringar av guld och fästa dem vid efodens båda axelstycken, nedtill på dess framsida, där den fästes ihop, ovanför efodens skärp.
Och man skall knyta fast bröstskölden med ett mörkblått snöre, Som går från dess ringar in i efodens ringar, så att den sitter ovanför efodens skärp, på det att bröstskölden icke må lossna från efoden.
Aron skall så bära Israels söners namn i domsskölden på sitt hjärta, när han går in helgedomen, för att bringa dem i åminnelse inför HERRENS ansikte beständigt.
Och du skall lägga urim och tummim in i domsskölden, så att de ligga på Arons hjärta, när han ingår inför HERRENS ansikte; och Aron skall så bära Israels barns dom på sitt hjärta inför HERRENS ansikte beständigt.
Efodkåpan skall du göra helt och hållet av mörkblått tyg;
och mitt på den skall vara en öppning för huvudet, och denna öppning skall omgivas med en vävd kant, likasom öppningen på en pansarskjorta, för att den icke slitas sönder.
Och på dess nedre fåll skall du sätta granatäpplen, gjorda av mörkblått, purpurrött och rosenrött garn, runt omkring fållen, och bjällror av guld mellan dessa runt omkring:
en bjällra av guld och så ett granatäpple, sedan en bjällra av guld och så åter ett granatäpple, runt omkring fållen på kåpan.
Och denna skall Aron hava på sig, när han gör tjänst, så att det höres, när han går in i helgedomen inför HERRENS ansikte, och när han går ut -- detta på det att han icke må dö.
Du skall ock göra en plåt av rent guld, och på den skall du rista, såsom man graverar signetringar: »Helgad åt HERREN.»
Och du skall fästa den vid ett mörkblått snöre, och den skall sitta på huvudbindeln; på framsidan av huvudbindeln skall den sitta.
Den skall sitta på Arons panna, och Aron skall bära den missgärning som vidlåder de heliga gåvor Israels barn bära fram, när de giva några heliga gåvor; den skall sitta på hans panna beständigt, för att de må bliva välbehagliga inför HERRENS ansikte.
Du skall ock väva en rutig livklädnad av vitt garn, och du skall göra en huvudbindel av vitt garn; och ett bälte skall du göra i brokig vävnad.
Också åt Arons söner skall du göra livklädnader, och du skall göra bälten åt dem; och huvor skall du göra åt dem, till ära och prydnad.
Och detta skall du kläda på din broder Aron och hans söner jämte honom;
och du skall smörja dem och företaga handfyllning med dem och helga dem till att bliva präster åt mig.
Och du skall göra åt dem benkläder av linne, som skyla deras blygd; dessa skola räcka från länderna ned på låren.
Och Aron och hans söner skola hava dem på sig, när de gå in i uppenbarelsetältet eller träda fram till altaret för att göra tjänst i helgedomen -- detta på det att de icke må komma att bära på missgärning och så träffas av döden.
Detta skall vara en evärdlig stadga för honom och hans avkomlingar efter honom.
Och detta är vad du skall göra med dem för att helga dem till att bliva präster åt mig: Tag en ungtjur och två vädurar, felfria djur,
och osyrat bröd och osyrade kakor, begjutna med olja, och osyrade tunnkakor, smorda med olja; av fint vetemjöl skall du baka dem.
Och du skall lägga dem i en och samma korg och bära fram dem i korgen såsom offergåva, när du för fram tjuren och de två vädurarna.
Därefter skall du föra Aron och hans söner fram till uppenbarelsetältets ingång och två dem med vatten.
Och du skall taga kläderna och sätta på Aron livklädnaden och efodkåpan och själva efoden och bröstskölden; och du skall fästa ihop alltsammans på honom med efodens skärp.
Och du skall sätta huvudbindeln på hans huvud och fästa det heliga diademet på huvudbindeln.
Och du skall taga smörjelseoljan och gjuta på hans huvud och smörja honom.
Och du skall föra fram hans söner och sätta livklädnader på dem.
Och du skall omgjorda dem, Aron och hans söner, med bälten och binda huvor på dem.
Och de skola hava prästadömet såsom en evärdlig rätt.
Så skall du företaga handfyllning med Aron och hans söner.
Och du skall föra tjuren fram inför uppenbarelsetältet, och Aron och hans söner skola lägga sina händer på tjurens huvud.
Sedan skall du slakta tjuren inför HERRENS ansikte, vid ingången till uppenbarelsetältet.
Och du skall taga av tjurens blod och stryka med ditt finger på altarets hörn; men allt det övriga skall du gjuta ut vid foten av altaret.
Och du skall taga allt det fett som omsluter inälvorna, så ock leverfettet och båda njurarna med det fett som sitter på dem, och förbränna det på altaret.
Men köttet av tjuren och hans hud och hans orenlighet skall du bränna upp i eld utanför lägret.
Det är ett syndoffer.
Och du skall taga den ena väduren, och Aron och hans söner skola lägga sina händer på vädurens huvud.
Sedan skall du slakta väduren och taga hans blod och stänka på altaret runt omkring;
men själva väduren skall du dela i dess stycken, och du skall två inälvorna och fötterna och lägga dem på styckena och huvudet.
Och du skall förbränna hela väduren på altaret; det är ett brännoffer åt HERREN.
En välbehaglig lukt, ett eldsoffer åt HERREN är det.
Därefter skall du taga den andra väduren, och Aron och hans söner skola lägga sina händer på vädurens huvud.
Sedan skall du slakta väduren och taga av hans blod och bestryka Arons högra örsnibb och hans söners högra örsnibb och tummen på deras högra hand och stortån på deras högra fot; men det övriga blodet skall det stänka på altaret runt omkring.
Och du skall taga av blodet på altaret och av smörjelseoljan och stänka på Aron och hans kläder, och likaledes på hans söner och hans söners kläder; så bliver han helig, han själv såväl som hans kläder, och likaledes hans söner såväl som hans söners kläder.
Och du skall taga fettet av väduren, svansen och det fett som omsluter inälvorna, så ock leverfettet och båda njurarna med fettet på dem, därtill det högra lårstycket ty detta är handfyllningsväduren.
Och du skall taga en rundkaka, en oljebrödskaka och en tunnkaka ur korgen med de osyrade bröden, som står inför HERRENS ansikte.
Och du skall lägga alltsammans på Arons och hans söners händer och vifta det såsom ett viftoffer inför HERRENS ansikte.
Sedan skall du taga det ur deras: händer och förbränna det på altaret ovanpå brännoffret, till en välbehaglig lukt inför HERREN; det är ett eldsoffer åt HERREN.
Och du skall taga bringan av Arons handfyllningsvädur och vifta den såsom ett viftoffer inför HERRENS ansikte, och detta skall vara din del.
Så skall du helga viftoffersbringan och offergärdslåret, det som viftas och det som gives såsom offergärd, de delar av handfyllningsväduren, som skola tillhöra Aron och hans söner.
Och detta skall tillhöra Aron och; hans söner såsom en evärdlig rätt av Israels barn, ty det är en offergärd.
Det skall vara en gärd av Israels barn, av deras tackoffer, en gärd av dem åt HERREN.
Och Arons heliga kläder skola hans söner hava efter honom, för att de i dem må bliva smorda och mottaga handfyllning.
I sju dagar skall den av hans söner, som bliver präst i hans ställe, ikläda sig dem, den som skall gå in i uppenbarelsetältet för att göra tjänst i helgedomen.
Och du skall taga handfyllningsväduren och koka hans kött på en helig plats.
Och vädurens kött jämte brödet: som är i korgen skola Aron och hans söner äta vid ingången till uppenbarelsetältet; de skola äta detta,
det som har använts till att bringa försoning vid deras handfyllning och helgande, men ingen främmande får ta därav, ty det är heligt.
Och om något av handfyllningsköttet eller av brödet bliver över till följande morgon, så skall du i eld bränna upp detta som har blivit över; det får icke ätas, ty det är heligt.
Så skall du göra med Aron och hans söner, i alla stycken såsom jag har bjudit dig.
Sju dagar skall deras handfyllning vara.
Och var dag skall du offra en tjur såsom syndoffer till försoning och rena altaret, i det du bringar försoning för det; och du skall smörja det för att helga det.
I sju dagar skall du bringa försoning för altaret och helga det.
Så bliver altaret högheligt; var och en som kommer vid altaret bliver helig.
Och detta är vad du skall offra på altaret: två årsgamla lamm för var dag beständigt.
Det ena lammet skall du offra om morgonen, och det andra lammet skall du offra vid aftontiden,
och till det första lammet en tiondedels efa fint mjöl, begjutet med en fjärdedels hin olja av stötta oliver, och såsom drickoffer en fjärdedels hin vin.
Det andra lammet skall du offra vid aftontiden; med likadant spisoffer och drickoffer som om morgonen skall du offra det, till en välbehaglig lukt, ett eldsoffer åt HERREN.
Detta skall vara edert dagliga brännoffer från släkte till släkte, vid ingången till uppenbarelsetältet, inför HERRENS ansikte, där jag skall uppenbara mig för eder, för att där tala med dig.
Där skall jag uppenbara mig för Israels barn, och det rummet skall bliva helgat av min härlighet.
Och jag skall helga uppenbarelsetältet och altaret, och Aron och hans söner skall jag helga till att bliva präster åt mig.
Och jag skall bo mitt ibland Israels barn och vara deras Gud.
Och de skola förnimma att jag är HERREN, deras Gud, som förde dem ut ur Egyptens land, för att jag skulle bo mitt ibland dem.
Jag är HERREN, deras Gud.
Och du skall göra ett altare för att antända rökelse därpå, av akacieträ skall du göra det.
Det skall vara en aln långt och en aln brett -- en liksidig fyrkant -- och två alnar högt; dess horn skola vara i ett stycke därmed.
Och du skall överdraga det med rent guld, dess skiva, dess väggar runt omkring och dess hörn; och du skall göra en rand av guld därpå runt omkring.
Och du skall till det göra två ringar av guld och sätta dem nedanför randen, på dess båda sidor; på de båda sidostyckena skall du sätta dem.
De skola vara där, för att stänger må skjutas in i dem, så att man med dem kan bära altaret.
Och du skall göra stängerna av akacieträ och överdraga dem med guld.
Och du skall ställa det framför den förlåt som hänger framför vittnesbördets ark, så att det står framför nådastolen, som är ovanpå vittnesbördet, där jag skall uppenbara mig för dig.
Och Aron skall antända välluktande rökelse därpå; var morgon, när han tillreder lamporna, skall han antända rökelse;
och likaledes skall Aron antända rökelse, när han vid aftontiden sätter upp lamporna.
Detta skall vara det dagliga rökoffret inför HERRENS ansikte, från släkte till släkte.
I skolen icke låta någon främmande rökelse komma därpå, ej heller brännoffer eller spisoffer; och intet drickoffer skolen utgjuta därpå.
Och Aron skall en gång om året bringa försoning för dess horn; med blod av försoningssyndoffret skall han en gång om året bringa försoning för det, släkte efter släkte.
Det är högheligt för HERREN.
Och HERREN talade till Mose och sade:
När du räknar antalet av Israels barn, nämligen av dem som inmönstras, skall vid mönstringen var och en giva åt HERREN en försoningsgåva för sig, på det att ingen hemsökelse må drabba dem vid mönstringen.
Detta är vad var och en som upptages bland de inmönstrade skall giva: en halv sikel, efter helgedomssikelns vikt -- sikeln räknad till tjugu gera -- en halv sikel såsom offergärd åt HERREN,
Var och en som upptages bland de inmönstrade, var och en som är tjugu år gammal eller därutöver, skall giva detta såsom offergärd åt HERREN.
Den rike skall icke giva mer och den fattige icke mindre än en halv sikel, när I given offergärden åt HERREN, till att bringa försoning för eder.
Och du skall taga försoningspenningarna av Israels barn och använda dem till arbetet vid uppenbarelsetältet.
Så skall ske, för att Israels barn må vara i åminnelse inför HERRENS ansikte, och för att försoning må bringas för eder.
Och HERREN talade till Mose och sade:
Du skall ock göra ett bäcken av koppar med en fotställning av koppar, till tvagning, och ställa det mellan uppenbarelsetältet och altaret och gjuta vatten däri.
Och Aron och hans söner skola två sina händer och fötter med vatten därur.
När de gå in i uppenbarelsetältet, skola de två sig med vatten, på del att de icke må dö; så ock när de träda fram till altaret för att göra tjänst genom att antända eldsoffer åt HERREN.
De skola två sina händer och fötter, på det att de icke må dö.
Och detta skall vara en evärdlig stadga för dem: för honom själv och hans avkomlingar från släkte till släkte.
Och HERREN talade till Mose och sade:
Tag dig ock kryddor av yppersta slag: fem hundra siklar myrradropp, hälften så mycket kanel av finaste slag, alltså två hundra femtio siklar, likaledes två hundra femtio siklar kalmus av finaste slag,
därtill fem hundra siklar kassia, efter helgedomssikelns vikt, och en hin olivolja.
Och du skall av detta göra en helig smörjelseolja, en konstmässigt beredd salva; det skall vara en helig smörjelseolja.
Och du skall därmed smörja uppenbarelsetältet, vittnesbördets ark,
bordet med alla dess tillbehör, ljusstaken med dess tillbehör, rökelsealtaret,
brännoffersaltaret med alla dess tillbehör, äntligen bäckenet med dess fotställning.
Och du skall helga dem, så att de bliva högheliga; var och en som sedan kommer vid dem bliver helig.
Och Aron och hans söner skall du smörja, och du skall helga dem till att bliva präster åt mig.
Och till Israels barn skall du tala och säga: Detta skall vara min heliga smörjelseolja hos eder, från släkte till släkte.
På ingen annan människas kropp må den komma, ej heller mån I göra någon annan så sammansatt som denna.
Helig är den, helig skall den vara för eder.
Den som bereder en sådan salva, och den som använder något därav på någon främmande, han skall utrotas ur sin släkt.
Ytterligare sade HERREN till Mose: Tag dig välluktande kryddor, stakte och sjönagel och galban, och jämte dessa vällukter rent rökelseharts, lika mycket av vart slag,
och gör därav rökelse, en konstmässigt beredd blandning, saltad, ren, helig.
Och en del av den skall du stöta till pulver och lägga framför vittnesbördet i uppenbarelsetältet, där jag vill uppenbara mig för dig.
Höghelig skall den vara för eder.
Och ingen annan rökelse mån I göra åt eder så sammansatt som denna skall vara.
Helig skall den vara dig för HERREN.
Den som gör sådan för att njuta av dess lukt, han skall utrotas ur sin släkt.
Och HERREN talade till Mose och sade:
Se, jag har kallat och nämnt Besalel, son till Uri, son till Hur, av Juda stam;
och jag har uppfyllt honom med Guds Ande, med vishet och förstånd och kunskap och med allt slags slöjdskicklighet,
till att tänka ut konstarbeten, till att arbeta i guld, silver och koppar,
till att snida stenar för infattning och till att snida i trä, korteligen, till att utföra alla slags arbeten.
Och se, jag har givit honom till medhjälpare Oholiab, Ahisamaks son, av Dans stam, och åt alla edra konstförfarna män har jag givit vishet i hjärtat.
Dessa skola kunna göra allt vad jag har bjudit dig:
uppenbarelsetältet, vittnesbördets ark, nådastolen därpå, alla uppenbarelsetältets tillbehör,
bordet med dess tillbehör, den gyllene ljusstaken med alla dess tillbehör, rökelsealtaret,
brännoffersaltaret med alla dess tillbehör, bäckenet med dess fotställning,
de stickade kläderna och prästen Arons andra heliga kläder, så och hans söners prästkläder,
äntligen smörjelseoljan och den välluktande rökelsen till helgedomen.
De skola utföra sitt arbete i alla stycken såsom jag har bjudit dig.
Och HERREN talade till Mose och sade:
Tala du till Israels barn och säg: Mina sabbater skolen I hålla, ty de äro ett tecken mellan mig och eder, från släkte till släkte, för att I skolen veta att jag är HERREN, som helgar eder.
Så hållen nu sabbaten, ty den skall vara eder helig.
Den som ohelgar den skall straffas med döden; ty var och en som på den dagen gör något arbete, han skall utrotas ur sin släkt.
Sex dagar skall arbete göras, men på sjunde dagen är vilosabbat, en HERRENS helgdag.
Var och en som gör något arbete på sabbatsdagen skall straffas med döden.
Och Israels barn skola hålla sabbaten, så att de fira den släkte efter släkte, såsom ett evigt förbund.
Den skall vara ett evärdligt tecken mellan mig och Israels barn; ty på sex dagar gjorde HERREN himmel och jord, men på sjunde dagen vilade han och tog sig ro.
När han nu hade talat ut med; Mose på Sinai berg, gav han honom vittnesbördets två tavlor, tavlor av sten, på vilka Gud hade skrivit med sitt finger.
Men när folket såg att Mose dröjde att komma ned från berget, församlade de sig omkring Aron och sade till honom: »Upp, gör oss en gud som kan gå framför oss; ty vi veta icke vad som har vederfarits denne Mose, honom som förde oss upp ur Egyptens land.»
Då sade Aron till dem: »Tagen guldringarna ut ur öronen på edra hustrur, edra söner och edra döttrar, och bären dem till mig.
Då tog allt folket av sig guldringarna som de hade i öronen, och de buro dem till Aron;
och han tog emot guldet av dem och formade det med en mejsel och gjorde därav en gjuten kalv.
Och de sade: »Detta är din Gud, Israel, han som har fört dig upp ur Egyptens land.»
När Aron såg detta, byggde han ett altare åt honom.
Och Aron lät utropa och säga: »I morgon bliver en HERRENS högtid.»
Dagen därefter stodo de bittida upp och offrade brännoffer och buro fram tackoffer, och folket satte sig ned till att äta och dricka, och därpå stodo de upp till att leka.
Då sade HERREN till Mose: »Gå ditned, ty ditt folk, som du har fört upp ur Egyptens land, har tagit sig till, vad fördärvligt är.
De hava redan vikit av ifrån den väg som jag bjöd dem gå; de hava gjort sig en gjuten kalv.
Den hava de tillbett, åt den hava de offrat, och sagt: 'Detta är din Gud, Israel, han som har fört dig upp ur Egyptens land.»
Och HERREN sade ytterligare till Mose: »Jag ser att detta folk är ett hårdnackat folk.
Så låt mig nu vara, på det att min vrede må brinna mot dem, och på det att jag må förgöra dem; dig vill jag sedan göra till ett stort folk.»
Men Mose bönföll inför HERREN, sin Gud, och sade: »HERRE, varför skulle din vrede brinna mot ditt folk, som du med stor kraft och stark hand har fört ut ur Egyptens land?
Varför skulle egyptierna få säga: 'Till deras olycka har han fört dem ut, till att dräpa dem bland bergen och förgöra dem från jorden'?
Vänd dig ifrån din vredes glöd, och ångra det onda du nu har i sinnet mot ditt folk.
Tänk på Abraham, Isak och Israel, dina tjänare, åt vilka du med ed vid dig själv har givit det löftet: 'Jag skall göra eder säd talrik såsom stjärnorna på himmelen, och hela det land som jag har talat om skall jag giva åt eder säd, och de skola få det till evärdlig arvedel.'»
Då ångrade HERREN det onda som han hade hotat att göra mot sitt folk.
Och Mose vände sig om och steg ned från berget, och han hade med sig vittnesbördets två tavlor.
Och på tavlornas båda sidor var skrivet både på den ena sidan och på den andra var skrivet.
Och tavlorna voro gjorda av Gud, och skriften var Guds skrift, inristad på tavlorna.
När Josua nu hörde huru folket skriade, sade han till Mose: »Krigsrop höres i lägret.»
Men han svarade: »Det är varken segerrop som höres, ej heller är det ett ropande såsom efter nederlag; det är sång jag hör.»
När sedan Mose kom närmare lägret och fick se kalven och dansen, upptändes hans vrede, och han kastade tavlorna ifrån sig och slog sönder dem nedanför berget.
Sedan tog han kalven som de hade gjort, och brände den i eld och krossade den till stoft; detta strödde han i vattnet och gav det åt Israels barn att dricka.
Och Mose sade till Aron: »Vad har folket gjort dig, eftersom du har kommit dem att begå en så stor synd?»
Aron svarade: »Min herres vrede må icke upptändas; du vet själv att detta folk är ont.
De sade till mig: 'Gör oss en gud som kan gå framför oss; ty vi veta icke vad som har vederfarits denne Mose, honom som förde oss upp ur Egyptens land.'
Då sade jag till dem: 'Den som har guld tage det av sig'; och de gåvo det åt mig.
Och jag kastade det i elden, och så kom kalven till.»
Då nu Mose såg att folket var lössläppt, eftersom Aron, till skadeglädje för deras fiender, hade släppt dem lösa,
ställde han sig i porten till lägret och ropade: »Var och en som hör HERREN till komme hit till mig.»
Då församlade sig till honom alla Levi barn.
Och han sade till dem: »Så säger HERREN, Israels Gud: Var och en binde sitt svärd vid sin länd.
Gån så igenom lägret, fram och tillbaka, från den ena porten till den andra, Och dräpen vem I finnen, vore det också broder eller vän eller frände.
Och Levi barn gjorde såsom Mose hade sagt; och på den dagen föllo av folket vid pass tre tusen män.
Och Mose sade: »Eftersom I nu haven stått emot edra egna söner och bröder, mån I i dag taga handfyllning till HERRENS tjänst, för att välsignelse i dag må komma över eder.»
Dagen därefter sade Mose till folket: »I haven begått en stor synd.
Jag vill nu stiga upp till HERREN och se till, om jag kan bringa försoning för eder synd.»
Och Mose gick tillbaka till HERREN och sade: »Ack, detta folk har begått en stor synd; de hava gjort sig en gud av guld.
Men förlåt dem nu deras synd; varom icke, så utplåna mig ur boken som du skriver i.»
Men HERREN svarade Mose: »Den som har syndat mot mig, honom skall jag utplåna ur min bok.
Gå nu och för folket dit jag har sagt dig; se, min ängel skall gå framför dig.
Men när min hemsökelses dag kommer, skall jag på dem hemsöka deras synd.»
Så straffade HERREN folket, därför att de hade gjort kalven, den som Aron gjorde.
Och HERREN sade till Mose: »Upp, drag åstad härifrån med folket som du har fört upp ur Egyptens land, och begiv dig till det land som jag med ed har lovat åt Abraham, Isak och Jakob, i det jag sade: 'Åt din säd skall jag giva det.'
Jag skall sända en ängel framför dig och förjaga kananéerna, amoréerna, hetiterna, perisséerna, hivéerna och jebuséerna,
för att du må komma till ett land som flyter av mjölk och honung.
Ty eftersom du är ett hårdnackat folk, vill jag icke själv draga upp med dig; jag kunde då förgöra dig under vägen.»
När folket hörde detta stränga tal, blevo de sorgsna, och ingen tog sina smycken på sig.
Och HERREN sade till Mose: »Säg till Israels barn: I ären ett hårdnackat folk.
Om jag allenast ett ögonblick droge med dig, skulle jag förgöra dig.
Men lägg nu av dig dina smycken, så vill jag se till, vad jag skall göra med dig.»
Så togo då Israels barn av sig sina smycken och voro utan dem allt ifrån vistelsen vid Horebs berg.
Men Mose hade för sed att taga tältet och slå upp det ett stycke utanför lägret; och han kallade det »uppenbarelsetältet».
Och var och en som ville rådfråga HERREN måste gå ut till uppenbarelsetältet utanför lägret.
Och så ofta Mose gick ut till tältet, stod allt folket upp, och var och en ställde sig vid ingången till sitt tält och skådade efter Mose, till dess han hade kommit in i tältet.
Och så ofta Mose kom in i tältet, steg molnstoden ned och blev stående vid ingången till tältet; och han talade med Mose.
Och allt folket såg molnstoden stå vid ingången till tältet; då föll allt folket ned och tillbad, var och en vid ingången till sitt tält.
Och HERREN talade med Mose ansikte mot ansikte, såsom när den ena människan talar med den andra.
Sedan vände Mose tillbaka till lägret; men hans tjänare Josua, Nuns son, en ung man, lämnade icke tältet.
Och Mose sade till HERREN: »Väl säger du till mig: 'För detta folk ditupp'; men du har icke låtit mig veta vem du vill sända med mig Du har dock sagt: 'Jag känner dig vid namn, och du har funnit nåd för mina ögon.'
Om jag alltså har funnit nåd för dina ögon, så låt mig se dina vägar och lära känna dig; jag vill ju finna nåd för dina ögon.
Och se därtill, att detta folk är ditt folk.»
Han sade: »Skall jag då själv gå med och föra dig till ro?»
Han svarade honom: »Om du icke själv vill gå med, så låt oss alls icke draga upp härifrån.
Ty varigenom skall man kunna veta att jag och ditt folk hava funnit nåd för dina ögon, om icke därigenom att du går med oss, så att vi, jag och ditt folk, utmärkas framför alla andra folk på jorden?»
HERREN svarade Mose: »Vad du nu har begärt skall jag ock göra; ty du har funnit nåd för mina ögon, och jag känner dig vid namn.»
Då sade han: »Låt mig alltså se din härlighet.»
Han svarade: »Jag skall låta all min skönhet gå förbi dig där du står, och jag skall utropa namnet 'HERREN' inför dig; jag skall vara nådig mot den jag vill vara nådig emot, och skall förbarma mig över den jag vill förbarma mig över.
Ytterligare sade han: »Mitt ansikte kan du dock icke få se, ty ingen människa kan se mig och leva.»
Därefter sade HERREN: »Se, här är en plats nära intill mig; ställ dig där på klippan.
När nu min härlighet går förbi, skall jag låta dig stå där i en klyfta på berget, och jag skall övertäcka dig med min hand, till dess jag har gått förbi.
Sedan skall jag taga bort min hand, och då skall du få se mig på ryggen; men mitt ansikte kan ingen se.»
Och HERREN sade till Mose: »Hugg ut åt dig två stentavlor, likadana som de förra voro, så vill jag skriva på tavlorna samma ord som stodo på de förra tavlorna, vilka du slog sönder.
Och var redo till i morgon, du skall då på morgonen stiga upp på Sinai berg och ställa dig på toppen av berget, mig till mötes,
men ingen må stiga upp med dig, och på hela berget för ingen annan visa sig; ej heller må får och fäkreatur gå i bet framemot detta berg.»
Och han högg ut två stentavlor likadana som de förra voro.
Och bittida följande morgon begav sig Mose upp på Sinai berg, såsom HERREN hade bjudit honom, och tog de två stentavlorna med sig.
Då steg HERREN ned i molnskyn.
Och han ställde sig där nära intill honom och åkallade HERRENS namn.
Och HERREN gick förbi honom, där han stod, och utropade: »HERREN!
HERREN! -- en Gud, barmhärtig och nådig, långmodig och stor i mildhet och trofasthet,
som bevarar nåd mot tusenden, som förlåter missgärning och överträdelse och synd, men som ingalunda låter någon bliva ostraffad, utan hemsöker fädernas missgärning på barn och barnbarn och efterkommande i tredje och fjärde led.»
Då böjde Mose sig med hast ned mot jorden och tillbad
och sade: »Om jag har funnit nåd för dina ögon, Herre, så må Herren gå med oss.
Ty väl är det ett hårdnackat folk, men du vill ju förlåta oss vår missgärning och synd och taga oss till din arvedel.»
Han svarade: »Välan, jag vill sluta ett förbund.
Inför hela ditt folk skall jag göra under, sådana som icke hava blivit gjorda i något land eller bland något folk.
Och hela det folk som du tillhör skall se att HERRENS gärningar äro underbara, de som jag skall göra med dig.
Håll de bud som jag i dag giver dig.
Se, jag skall förjaga för dig amoréerna, kananéerna, hetiterna, perisséerna, hivéerna och jebuséerna.
Tag dig till vara för att sluta förbund med inbyggarna i det land dit du kommer, och låt dem icke bliva till en snara bland eder.
Fastmer skolen I bryta ned deras altaren och slå sönder deras stoder och hugga ned deras Aseror.
Ja, du skall icke tillbedja någon annan gud, ty HERREN heter Nitälskare; en nitälskande Gud är han.
Du må icke sluta något förbund med landets inbyggare.
Ty i trolös avfällighet löpa de efter sina gudar och offra åt sina gudar; och när de då inbjuda dig, kommer du att äta av deras offer;
du tager ock deras döttrar till hustrur åt dina söner, och när då deras döttrar i avfällighet löpa efter sina gudar, skola de förleda dina söner till att likaledes löpa efter deras gudar.
Gjutna gudar skall du icke göra åt dig.
Det osyrade brödets högtid skall, du hålla: i sju dagar skall du äta osyrat bröd, såsom jag har bjudit dig, på den bestämda tiden i månaden Abib; ty i månaden Abib drog du ut ur Egypten.
Allt det som öppnar moderlivet skall höra mig till, också allt hankön bland din boskap, som öppnar moderlivet, såväl av fäkreaturen som av småboskapen.
Men vad som bland åsnor öppnar moderlivet skall du lösa med ett får, och om du icke vill lösa det, skall du krossa nacken på det.
Var förstfödd bland dina söner skall du läsa.
Och ingen skall med tomma händer träda fram inför mitt ansikte.
Sex dagar skall du arbeta, men på sjunde dagen skall du hålla vilodag; både under plöjningstiden och under skördetiden skall du hålla vilodag.
Och veckohögtiden skall du hålla, för förstlingen av veteskörden, så ock bärgningshögtiden, när året har gått till ända.
Tre gånger om året skall allt ditt mankön träda fram inför HERRENS, din herres, Israels Guds, ansikte.
Ty jag skall fördriva folk för dig och utvidga ditt område; och ingen skall stå efter ditt land, när du drager upp, tre gånger om året, för att träda fram inför HERRENS, din Guds, ansikte.
Du skall icke offra blodet av mitt slaktoffer jämte något som är syrat.
Och påskhögtidens slaktoffer skall icke lämnas kvar över natten till morgonen.
Det första av din marks förstlingsfrukter skall du föra till HERRENS, din Guds, hus.
Du skall icke koka en killing i dess moders mjölk.»
Och HERREN sade till Mose: »Teckna upp åt dig dessa ord; ty i enlighet med dessa ord har jag slutit ett förbund med dig och med Israel.»
Och han blev kvar där hos HERREN i fyrtio dagar och fyrtio nätter, utan att äta och utan att dricka.
Och han skrev på tavlorna förbundets ord, de tio orden.
När sedan Mose steg ned från Sinai berg, och på vägen ned från berget hade vittnesbördets två tavlor med sig, visste han icke att hans ansiktes hy hade blivit strålande därav att han hade talat med honom.
Och när Aron och alla Israels barn sågo huru Moses ansiktes hy strålade, fruktade de för att komma honom nära.
Men Mose ropade till dem; då vände Aron och menighetens alla hövdingar tillbaka till honom, och Mose talade till dem.
Därefter kommo alla Israels barn fram till honom, och han gav dem alla de bud som HERREN hade förkunnat för honom på Sinai berg.
Och när Mose hade slutat sitt tal till dem, hängde han ett täckelse för sitt ansikte.
Men så ofta Mose skulle träda inför HERRENS ansikte för att tala med honom, lade han av täckelset, till dess han åter gick ut.
Och sedan han hade kommit ut, förkunnade han för Israels barn det som hade blivit honom bjudet.
Då sågo Israels barn var gång huru Moses ansiktes by strålade, och Mose hängde då åter täckelset över sitt ansikte, till dess han ånyo skulle gå in för att tala med honom.
Och Mose församlade Israels barns hela menighet och sade till dem: »Detta är vad HERREN har bjudit eder att göra:
Sex dagar skall arbete göras, men på sjunde dagen skolen I hava helgdag, en HERRENS vilosabbat.
Var och en som på den dagen gör något arbete skall dödas.
I skolen icke tända upp eld på: sabbatsdagen, var I än ären bosatta.
Och Mose sade till Israels barns hela menighet: »Detta är vad HERREN har bjudit och sagt:
Låten bland eder upptaga en gärd åt HERREN, så att var och en som har ett därtill villigt hjärta bär fram denna gård åt HERREN: guld, silver och koppar,
mörkblått, purpurrött, rosenrött och vitt garn och gethår,
rödfärgade vädurskinn, tahasskinn, akacieträ,
olja till ljusstaken, kryddor till smörjelseoljan och till den välluktande rökelsen,
äntligen onyxstenar och infattningsstenar, till att användas för efoden och för bröstskölden.
Och alla konstförfarna män bland eder må komma och förfärdiga allt vad HERREN har bjudit:
tabernaklet, dess täckelse och överdraget till detta, dess häktor, bräder, tvärstänger, stolpar och fotstycken,
arken med dess stänger, nådastolen och den förlåt som skall hänga framför den,
bordet med dess stänger och alla dess tillbehör och skådebröden,
ljusstaken med dess tillbehör och dess lampor, oljan till ljusstaken,
rökelsealtaret med dess stänger, smörjelseoljan och den välluktande rökelsen, förhänget för ingången till tabernaklet,
brännoffersaltaret med tillhörande koppargaller, dess stänger och alla dess tillbehör, bäckenet med dess fotställning,
omhängena till förgården, dess stolpar och fotstycken, förhänget för porten till förgården,
tabernaklets pluggar och förgårdens pluggar med deras streck,
äntligen de stickade kläderna till tjänsten i helgedomen och prästen Arons andra heliga kläder, så ock hans söners prästkläder.»
Och Israels barns hela menighet gick sin väg bort ifrån Mose.
Sedan kommo de tillbaka, var och en som av sitt hjärta manades därtill; och var och en som hade en därtill villig ande bar fram en gärd åt HERREN till förfärdigande av uppenbarelsetältet och till allt arbete därvid och till de heliga kläderna.
De kommo, både män och kvinnor, och framburo, var och en efter sitt hjärtas villighet, spännen, örringar, fingerringar och halssmycken, alla slags klenoder av guld, var och en som kunde offra åt HERREN någon gåva av guld.
Och var och en som hade i sin ägo mörkblått, purpurrött, rosenrött eller vitt garn eller gethår eller rödfärgade vädurskinn eller tahasskinn bar fram det.
Och var och en som kunde giva såsom gärd något av silver eller koppar bar fram sin gärd åt HERREN.
Och var och en som hade i sin ägo akacieträ till förfärdigande av något slags arbete bar fram det.
Och alla konstförfarna kvinnor spunno med sina händer mörkblått, purpurrött, rosenrött och vitt garn och buro fram sin spånad;
och alla kvinnor som av sitt hjärta manades därtill och hade lärt konsten spunno gethår.
Och hövdingarna buro fram onyxstenar och infattningsstenar, till att användas för efoden och för bröstskölden,
vidare kryddor och olja, till att användas för ljusstaken och smörjelseoljan och den välluktande rökelsen.
Var och en av Israels barn, man eller kvinna, vilkens hjärta var villigt att bära fram något till förfärdigande av allt det som HERREN genom Mose hade bjudit att man skulle göra, bar fram sin frivilliga gåva åt HERREN.
och Mose sade till Israels barn: »Sen, HERREN har kallat och nämnt Besalel, son till Uri, son till Hur, av Juda stam;
och han har uppfyllt honom med Guds Ande, med vishet, med förstånd och kunskap och med allt slags slöjdskicklighet,
både till att tänka ut konstarbeten och till att arbeta i guld, silver och koppar,
till att smida stenar för infattning: och till att snida i trä, korteligen, till att utföra alla slags konstarbeten.
Åt honom och åt Oholiab, Ahisamaks son, av Dans stam, har han ock givit förmåga att undervisa andra.
Han har uppfyllt deras hjärtan med vishet till att utföra alla slags snideriarbeten och konstvävnader och brokiga vävnader av mörkblått, purpurrött, rosenrött och vitt garn, så ock andra vävnader, korteligen, alla slags arbeten och särskilt konstvävnadsarbeten.
Och Besalel och Oholiab och alla andra konstförfarna män, åt vilka HERREN har givit vishet och förstånd till att veta huru de skola utföra allt arbete vid helgedomens förfärdigande, skola utföra det, i alla stycken såsom HERREN har bjudit.»
Därefter kallade Mose till sig Besalel och Oholiab och alla de andra konstförfarna männen, åt vilka HERREN hade givit vishet i hjärtat, alla som av sitt hjärta manades att träda fram för att utföra arbetet.
Och de mottogo från Mose hela den gärd som Israels barn hade burit fram till utförande av arbetet vid helgedomens förfärdigande.
Men man fortfor att bära fram till honom frivilliga gåvor, morgon efter morgon.
Då kommo alla de konstförfarna män som utförde allt arbetet till helgedomen, var och en från det arbete som han utförde,
och sade till Mose: »Folket bär fram mer än som behöves för att verkställa det arbete som HERREN har bjudit oss att utföra.»
Då bjöd Mose att man skulle låta utropa i lägret: »Ingen, vare sig man eller kvinna, må vidare arbeta för att göra något till helgedomen.»
Så avhölls folket ifrån att bära fram flera gåvor.
Ty vad man hade skaffat samman var tillräckligt för allt det arbete som skulle göras, och man hade till och med över.
Så gjorde nu alla de konstförfarna arbetarna tabernaklet av tio tygvåder; av tvinnat vitt garn och av mörkblått, purpurrött och rosenrött garn gjorde man dem, med keruber på, i konstvävnad.
Var våd gjordes tjuguåtta alnar lång och fyra alnar bred; alla våderna fingo samma mått.
Och man fogade tillhopa fem av våderna med varandra; likaså fogade man tillhopa de fem övriga våderna med varandra.
Och man satte öglor av mörkblått garn i kanten på den ena våden, ytterst på det hopfogade stycket; så gjorde man ock i kanten på den våd som satt ytterst i det andra hopfogade stycket.
Femtio öglor satte man på den ena våden, och femtio öglor satte man ytterst på motsvarande våd i det andra hopfogade stycket, så att öglorna svarade emot varandra.
Och man gjorde femtio häktor av guld och fogade våderna tillhopa med varandra medelst häktorna, så att tabernaklet utgjorde ett helt.
Man gjorde och tygvåder av gethår till ett täckelse över tabernaklet; elva sådana våder gjorde man.
Var våd gjordes trettio alnar lång och fyra alnar bred, de elva våderna fingo samma mått.
Fem av våderna fogade man tillhopa till ett särskilt stycke,
och likaledes de sex övriga våderna till ett särskilt stycke.
Och man satte femtio öglor i kanten på den våd som satt ytterst i det ena hopfogade stycket, och femtio öglor satte man i kanten på motsvarande våd i det andra hopfogade stycket.
Och man gjorde femtio häktor av koppar för att foga tillhopa täckelset, så att det kom att utgöra ett helt.
Vidare gjorde man ett överdrag av rödfärgade vädurskinn till täckelset, och ytterligare ett överdrag av tahasskinn att lägga ovanpå detta.
Bräderna till tabernaklet gjorde man av akacieträ och ställde dem upprätt.
Tio alnar långt och en och en halv aln brett gjordes vart bräde.
På vart bräde sattes två tappar, förbundna sinsemellan med en list; så gjorde man på alla bräderna till tabernaklet.
Och av tabernaklets bräder satte man tjugu på södra sidan, söderut.
Och man gjorde fyrtio fotstycken av silver att sätta under de tjugu bräderna, två fotstycken under vart bräde för dess två tappar.
Likaledes satte man på tabernaklets andra sida, den norra sidan, tjugu bräder,
med deras fyrtio fotstycken av silver, två fotstycken under vart bräde.
Men på baksidan av tabernaklet, västerut, satte man sex bräder.
Och två bräder satte man på tabernaklets hörn, på baksidan;
och vartdera av dessa var sammanfogat av två nedtill, och likaledes sammanhängande upptill, till den första ringen.
Så gjorde man med dem båda, i de båda hörnen.
Således blev det åtta bräder med tillhörande fotstycken av silver, sexton fotstycken, nämligen två fotstycken under vart bräde.
Och man gjorde tvärstänger av akacieträ, fem till de bräder som voro på tabernaklets ena sida,
och fem tvärstänger till de bräder som voro på tabernaklets andra sida, och fem tvärstänger till de bräder som voro på tabernaklets baksida, västerut.
Och man satte den mellersta tvärstången så, att den gick tvärs över, mitt på bräderna, från den ena ändan till den andra.
Och bräderna överdrog man med guld, och ringarna på dem, i vilka tvärstängerna skulle skjutas in, gjorde man av guld, och tvärstängerna överdrog man med guld.
Man gjorde ock förlåten av mörkblått, purpurrött, rosenrött och tvinnat vitt garn; man gjorde den i konstvävnad, med keruber på.
Och man gjorde till den fyra stolpar av akacieträ och överdrog dem med guld, och hakarna till dem gjordes av guld, och man göt till dem fyra fotstycken av silver.
Och man gjorde ett förhänge för ingången till tältet, i brokig vävnad av mörkblått, purpurrött, rosenrött och tvinnat vitt garn,
och till detta fem stolpar med deras hakar; och deras knoppar och deras kransar överdrog man med guld, och deras fem fotstycken gjordes av koppar.
Och Besalel gjorde arken av akacieträ, två och en halv aln lång, en och en halv aln bred och en och en halv aln hög.
Och han överdrog den med rent guld innan och utan; och han gjorde på den en rand av guld runt omkring.
Och han göt till den fyra ringar: av guld och satte dem över de fyra fötterna, två ringar på ena sidan och två ringar på andra sidan.
Och han gjorde stänger av akacieträ och överdrog dem med guld.
Och stängerna sköt han in i ringarna, på sidorna av arken, så att man kunde bära arken.
Och han gjorde en nådastol av rent guld, två och en halv aln lång och en och en halv aln bred.
Och han gjorde två keruber av guld; i drivet arbete gjorde han dem och satte dem vid de båda ändarna av nådastolen,
en kerub vid ena ändan och en kerub vid andra ändan.
I ett stycke med nådastolen gjorde han keruberna vid dess båda ändar.
Och keruberna bredde ut sina vingar och höllo dem uppåt, så att de övertäckte nådastolen med sina vingar, under det att de hade sina ansikten vända mot varandra; ned mot nådastolen vände keruberna sina ansikten.
Han gjorde ock bordet av akacieträ, två alnar långt, en aln brett och en och en halv aln högt.
Och han överdrog det med rent guld; och han gjorde en rand av guld därpå runt omkring.
Och runt omkring det gjorde han en list av en hands bredd, och runt omkring listen gjorde han en rand av guld.
Och han göt till bordet fyra ringar av guld och satte ringarna i de fyra hörnen vid de fyra fötterna.
Invid listen sattes ringarna, för att stängerna skulle skjutas in i dem, så att man kunde bära bordet.
Och han gjorde stängerna av akacieträ och överdrog dem med guld; så kunde man bära bordet.
Och han gjorde kärlen till bordet av rent guld, faten och skålarna, bägarna och kannorna med vilka man skulle utgjuta drickoffer.
Han gjorde ock ljusstaken av rent guld.
I drivet arbete gjorde han ljusstaken med dess fotställning och dess mittelrör; kalkarna därpå, kulor och blommor, gjordes i ett stycke med den.
Och sex armar utgingo från ljusstakens sidor, tre armar från ena sidan och tre armar från andra sidan.
På den ena armen sattes tre kalkar, liknande mandelblommor, vardera bestående av en kula och en blomma, och på den andra armen sammalunda tre kalkar, liknande mandelblommor, vardera bestående av en kula och en blomma; så gjordes på de sex armar som utgingo från ljusstaken
Men på själva ljusstaken sattes fyra kalkar, liknande mandelblommor, med sina kulor och blommor.
En kula sattes under det första armparet som utgick från ljusstaken, i ett stycke med den, och en kula under det andra armparet som utgick från ljusstaken, i ett stycke med den, och en kula under det tredje armparet som utgick från ljusstaken, i ett stycke med den: alltså under de sex armar som utgingo från den.
Deras kulor och armar gjordes i ett stycke med den, alltsammans ett enda stycke i drivet arbete av rent guld.
Och han gjorde till den sju lampor, så ock lamptänger och brickor till den av rent guld.
Av en talent rent guld gjorde han den med alla dess tillbehör.
Och han gjorde rökelsealtaret av akacieträ, en aln långt och en aln brett -- en liksidig fyrkant -- och två alnar högt; dess horn gjordes i ett stycke därmed.
Och han överdrog det med rent guld, dess skiva, dess väggar runt omkring och dess hörn; och han gjorde en rand av guld därpå runt omkring.
Och han gjorde till det två ringar av guld och satte dem nedanför randen, på dess båda sidor, på de båda sidostyckena, för att stänger skulle skjutas in i dem, så att män med dem kunde bära altaret.
Och han gjorde stängerna av akacieträ och överdrog dem med guld.
Han gjorde ock den heliga smörjelseoljan och den rena, välluktande rökelsen, konstmässigt beredda.
Han gjorde ock brännoffersaltaret av akacieträ, fem alnar långt och fem alnar brett -- en liksidig fyrkant -- och tre alnar högt.
Och han gjorde hörn därtill och satte dem i dess fyra hörn; i ett stycke därmed gjordes hörnen.
Och han överdrog det med koppar.
Och han gjorde altarets alla tillbehör, askkärlen, skovlarna, skålarna, gafflarna och fyrfaten.
Alla dess tillbehör gjorde han av koppar.
Och han gjorde till altaret ett galler, ett nätverk av koppar, och satte det under dess avsats, nedtill, så att det räckte upp till mitten.
Och han göt fyra ringar och satte dem i de fyra hörnen på koppargallret, för att stängerna skulle skjutas in i dem.
Och han gjorde stängerna av akacieträ och överdrog dem med koppar.
Och han sköt stängerna in i ringarna på altarets sidor, så att man kunde bära det med dem.
Ihåligt gjorde han det, av plankor.
Han gjorde ock bäckenet av koppar med dess fotställning av koppar och använde därtill speglar, som hade tillhört de kvinnor vilka hade tjänstgöring vid ingången till uppenbarelsetältet.
Han gjorde ock förgården.
För den södra sidan, söderut, gjordes omhängena till förgården av tvinnat sitt garn, hundra alnar långa;
till dem gjordes tjugu stolpar, och till dessa tjugu fotstycken, av koppar, men stolparnas hakar och kransar gjordes av silver.
Likaledes gjordes de för norra sidan hundra alnar långa; till dem gjordes tjugu stolpar, och till dessa tjugu fotstycken, av koppar, men stolparnas hakar och kransar gjordes av silver.
Och för västra sidan gjordes omhängen som voro femtio alnar långa; till dem gjordes tio stolpar, och till dessa tio fotstycken, men stolparnas hakar och kransar gjordes av silver.
Och för framsidan, österut, gjordes de femtio alnar långa.
Omhängena gjordes femton alnar långa på ena sidan därav, med tre stolpar på tre fotstycken; likaledes gjordes omhängena på andra sidan femton alnar långa -- alltså lika på båda sidor om porten till förgården -- med tre stolpar på tre fotstycken.
Alla omhängena runt omkring förgården gjordes av tvinnat vitt garn;
och fotstyckena till stolparna gjordes av koppar, men stolparnas hakar och kransar gjordes av silver, och deras knoppar överdrogos med silver;
alla förgårdens stolpar försågos med kransar av silver.
Och förhänget för porten till förgården gjordes i brokig vävnad av mörkblått, purpurrött, rosenrött och tvinnat vitt garn, tjugu alnar långt och fem alnar högt, efter tygets bredd, i likhet med förgårdens omhängen;
och till det gjordes fyra stolpar på fyra fotstycken, av koppar; men deras hakar gjordes av silver, och deras knoppar överdrogos med silver, och deras kransar gjordes av silver.
Alla pluggarna till tabernaklet och till förgården runt omkring gjordes av koppar.
Följande är vad som beräknas hava åtgått till tabernaklet, vittnesbördets tabernakel, vilken beräkning gjordes efter Moses befallning genom leviternas försorg, under ledning av Itamar, prästen Arons son;
och Besalel, son till Uri, son till Hur, av Juda stam, förfärdigade allt vad HERREN hade bjudit Mose,
och till medhjälpare hade han Oholiab, Ahisamaks son, av Dans stam, en man kunnig i snideri och konstvävnad och i konsten att väva brokigt med mörkblått, purpurrött, rosenrött och vitt garn.
Det guld som användes till arbetet, vid förfärdigandet av hela helgedomen, det guld som hade blivit givet såsom offer, utgjorde sammanlagt tjugunio talenter och sju hundra trettio siklar, efter helgedomssikelns vikt.
Och det silver som gavs av dem i menigheten, vilka inmönstrades, utgjorde ett hundra talenter och ett tusen sju hundra sjuttiofem siklar, efter helgedomssikelns vikt.
En beka, det är en halv sikel, efter helgedomssikelns vikt, kom på var person, på var och en som upptogs bland de inmönstrade, var och en som var tjugu år gammal eller därutöver: sex hundra tre tusen fem hundra femtio personer.
Och de hundra talenterna silver användes till gjutningen av fotstyckena för helgedomen och av fotstyckena för förlåten, ett hundra talenter till ett hundra fotstycken, en talent till vart fotstycke.
Och de ett tusen sju hundra sjuttiofem siklarna användes till att göra hakar till stolparna och till att överdraga deras knoppar och göra kransar till dem.
Och den koppar som hade blivit given såsom offer utgjorde sjuttio talenter och två tusen fyra hundra siklar.
Därav gjorde man fotstyckena till uppenbarelsetältets ingång, så ock kopparaltaret med tillhörande koppargaller och altarets alla tillbehör,
vidare fotstyckena till förgården, runt omkring, och fotstyckena till förgårdens port, äntligen alla tabernaklets pluggar och alla förgårdens pluggar, runt omkring.
Och av det mörkblåa, det purpurröda och det rosenröda garnet gjorde man stickade kläder till tjänsten i helgedomen; och man gjorde de andra heliga kläderna som Aron skulle hava, såsom HERREN hade bjudit Mose.
Efoden gjorde man av guld och av mörkblått, purpurrött, rosenrött och tvinnat vitt garn.
Man hamrade ut guldet till tunna plåtar och skar dessa i trådar, så att man kunde väva in det i det mörkblåa, det purpurröda, det rosenröda och det vita garnet, med konstvävnad.
Till den gjorde man axelstycken, som skulle fästas ihop; vid sina båda ändar fästes den ihop.
Och skärpet, som skulle sitta på efoden och sammanhålla den, gjordes i ett stycke med den och av samma slags vävnad: av guld och av mörkblått, purpurrött, rosenrött och tvinnat vitt garn, allt såsom HERREN hade bjudit Mose.
Och onyxstenarna omgav man med flätverk av guld; på dem voro Israels söners namn inristade, på samma sätt som man graverar signetringar.
Och man satte dem på efodens axelstycken, för att stenarna skulle bringa Israels barn i åminnelse, allt såsom HERREN hade bjudit Mose.
Bröstskölden gjorde man i konstvävnad, i samma slags vävnad som efoden: av guld och av mörkblått, purpurrött, rosenrött och tvinnat vitt garn.
Bröstskölden gjordes liksidigt fyrkantig, i form av en väska gjorde man den: ett kvarter lång och ett kvarter bred, i form av en väska.
Och man besatte den med fyra rader stenar: i första raden en karneol, en topas och en smaragd;
i andra raden en karbunkel, en safir och en kalcedon;
i tredje raden en hyacint, en agat och en ametist;
i fjärde raden en krysolit, en onyx och en jaspis.
Med flätverk av guld blevo de omgivna i sina infattningar.
Stenarna voro tolv, efter Israels söners namn, en för vart namn; var sten bar namnet på en av de tolv stammarna, inristat på samma sätt som man graverar signetringar.
Och man gjorde till bröstskölden kedjor i virat arbete, såsom man gör snodder, av rent guld.
Man gjorde vidare två flätverk av guld och två ringar av guld och satte dessa båda ringar i två av bröstsköldens hörn.
Och man fäste de båda guldsnodderna vid de båda ringarna, i bröstsköldens hörn.
Och de två snoddernas båda andra ändar fäste man vid de två flätverken och fäste dem så vid efodens axelstycken på dess framsida.
Och man gjorde två andra ringar av guld och satte dem i bröstsköldens båda andra hörn, vid den kant därpå, som var vänd inåt mot efoden.
Och ytterligare gjorde man två ringar av guld och fäste dem vid efodens båda axelstycken, nedtill på dess framsida, där den fästes ihop, ovanför efodens skärp.
Och man knöt fast bröstskölden med ett mörkblått snöre, som gick från dess ringar in i efodens ringar, så att den satt ovanför efodens skärp, på det att bröstskölden icke skulle lossna från efoden, allt såsom HERREN hade bjudit Mose.
Efodkåpan gjorde man av vävt tyg, helt och hållet mörkblått.
Och mitt på kåpan gjordes en öppning, lik öppningen på en pansarskjorta; öppningen omgavs nämligen med en kant, för att den icke skulle slitas sönder.
Och på kåpans nedre fåll satte man granatäpplen, gjorda av mörkblått, purpurrött och rosenrött tvinnat garn.
Och man gjorde bjällror av rent guld och satte dessa bjällror mellan granatäpplena runt omkring fållen på kåpan, mellan granatäpplena:
en bjällra och så ett granatäpple, sedan en bjällra och så åter ett granatäpple, runt omkring fållen på kåpan, att bäras vid tjänstgöringen, såsom HERREN hade bjudit Mose.
Och man gjorde åt Aron och hans söner livklädnaderna av vitt garn, i vävt arbete,
huvudbindeln av vitt garn, högtidshuvorna av vitt garn och linnebenkläderna av tvinnat vitt garn,
äntligen bältet av tvinnat vitt garn och av mörkblått, purpurrött och rosenrött garn, i brokig vävnad, allt såsom HERREN hade bjudit Mose.
Och man gjorde plåten till det heliga diademet av rent guld, och på den skrev man, såsom man graverar signetringar: »Helgad åt HERREN.»
Och man fäste vid den ett mörkblått snöre och satte den ovanpå huvudbindeln, allt såsom HERREN hade bjudit Mose.
Så blev då allt arbetet på uppenbarelsetältets tabernakel fullbordat.
Israels barn utförde det; de gjorde i alla stycken såsom HERREN hade bjudit Mose.
Och de förde fram till Mose tabernaklet, dess täckelse och alla dess tillbehör, dess häktor, bräder, tvärstänger, stol par och fotstycken,
överdraget av rödfärgade vädurskinn och överdraget av tahasskinn och den förlåt som skulle hänga framför arken,
vidare vittnesbördets ark med dess stänger, så ock nådastolen,
bordet med alla dess tillbehör och skådebröden,
den gyllene ljusstaken, lamporna som skulle sättas på den och alla dess andra tillbehör, oljan till ljusstaken,
det gyllene altaret, smörjelseoljan och den välluktande rökelsen, förhänget för ingången till tältet,
kopparaltaret med tillhörande koppargaller, dess stänger och alla dess tillbehör, bäckenet med dess fotställning.
omhängena till förgården, dess stolpar och fotstycken, förhänget för porten till förgården, dess streck och pluggar, alla redskap till arbetet vid uppenbarelsetältets tabernakel
äntligen de stickade kläderna till tjänsten i helgedomen och prästen Arons andra heliga kläder, så ock hans söners prästkläder.
Såsom HERREN hade bjudit Mose så hade Israels barn i alla stycken gjort allt arbete.
Och Mose besåg allt arbetet och fann att de hade utfört det, att de hade gjort såsom HERREN hade bjudit.
Och Mose välsignade dem
Och HERREN talade till Mose och sade:
»När den första månaden ingår, skall du på första dagen i månaden uppsätta uppenbarelsetältets tabernakel.
Och du skall däri sätta vittnesbördets ark och hänga förlåten framför arken.
Och du skall föra bordet ditin och lägga upp på detta vad där skall vara upplagt; och du skall föra ditin ljusstaken och sätta upp lamporna på den.
Och du skall ställa det gyllene rökelsealtaret framför vittnesbördets ark; och du skall sätta upp förhänget för ingången till tabernaklet.
Och brännoffersaltaret skall du ställa framför ingången till uppenbarelsetältets tabernakel.
Och du skall ställa bäckenet mellan uppenbarelsetältet och altaret och gjuta vatten däri.
Och du skall sätta upp förgårdshägnaden runt omkring och hänga upp förhänget för porten till förgården.
Och du skall taga smörjelseoljan och smörja tabernaklet och allt vad däri är och helga det jämte alla dess tillbehör, så att det bliver heligt.
Du skall ock smörja brännoffersaltaret jämte alla dess tillbehör och helga altaret; så bliver altaret högheligt.
Du skall ock smörja bäckenet jämte dess fotställning och helga det.
Därefter skall du föra Aron och hans söner fram till uppenbarelsetältets ingång och två dem med vatten.
Och du skall sätta på Aron del heliga kläderna, och smörja honom och helga honom till att bliva präst åt mig
Och du skall föra fram hans söner och sätta livklädnader på dem.
Och du skall smörja dem, såsom du smorde deras fader, till att bliva präster åt mig.
Så skall denna deras smörjelse bliva för dem en invigning till ett evärdligt prästadöme, släkte efter släkte.
Och Mose gjorde detta; han gjorde i alla stycken såsom HERREN hade bjudit honom.
Så blev då tabernaklet uppsatt i första månaden av andra året, på första dagen i månaden.
Då satte Mose upp tabernaklet.
Han lade ut dess fotstycken, ställde fast dess bräder, sköt in dess tvärstänger och satte upp dess stolpar.
Och han bredde täckelset över tabernaklet och lade ovanpå täckelset dess överdrag allt såsom HERREN hade bjudit Mose.
Och han tog vittnesbördet och lade det in i arken och satte stängerna på arken; och han satte nådastolen ovanpå arken.
Sedan förde han arken in i tabernaklet och satte upp förlåten som skulle hänga framför arken, och hängde så för vittnesbördets ark, allt såsom HERREN hade bjudit Mose.
Och han satte bordet i uppenbarelsetältet, vid tabernaklets norra sida, utanför förlåten,
och lade upp på detta de bröd som skulle vara upplagda inför HERRENS ansikte, allt såsom HERREN hade bjudit Mose.
Och han ställde ljusstaken in i uppenbarelsetältet, mitt emot bordet, på tabernaklets södra sida,
och satte upp lamporna inför HERRENS ansikte, såsom HERREN hade bjudit Mose.
Och han ställde det gyllene altaret in i uppenbarelsetältet, framför förlåten,
och antände välluktande rökelse därpå, såsom HERREN hade bjudit Mose.
Och han satte upp förhänget för ingången till tabernaklet.
Och brännoffersaltaret ställde han vid ingången till uppenbarelsetältets tabernakel och offrade brännoffer och spisoffer därpå, såsom HERREN hade bjudit Mose.
Och han ställde bäckenet mellan uppenbarelsetältet och altaret och göt vatten till tvagning däri.
Och Mose och Aron och hans söner tvådde sedermera sina händer och fötter med vatten därur;
så ofta de skulle gå in i uppenbarelsetältet eller träda fram till altaret, tvådde de sig, såsom HERREN hade bjudit Mose.
Och han satte upp förgårdshägnaden runt omkring tabernaklet och altaret, och hängde upp förhänget för porten till förgården.
Så fullbordade Mose allt arbetet.
Då övertäckte molnskyn uppenbarelsetältet, och HERRENS härlighet uppfyllde tabernaklet;
och Mose kunde icke gå in i uppenbarelsetältet, eftersom molnskyn vilade däröver och HERRENS härlighet uppfyllde tabernaklet.
Och så ofta molnskyn höjde sig från tabernaklet, bröto Israels barn upp; så gjorde de under hela sin vandring.
Men så länge molnskyn icke höjde sig, bröto de icke upp, utan stannade ända till den dag då den åter höjde sig.
Ty HERRENS molnsky vilade om dagen över tabernaklet, och om natten var eld i den; så var det inför alla Israels barns ögon under hela deras vandring.
Och HERREN kallade på Mose och talade till honom ur uppenbarelsetältet och sade:
Tala till Israels barn och säg till dem: När någon bland eder vill bära fram ett offer åt HERREN, skolen I taga edert offer av boskapen, antingen av fäkreaturen eller av småboskapen.
Om han vill bära fram ett brännoffer av fäkreaturen, så skall han därtill taga ett felfritt djur av hankön och föra det fram till uppenbarelsetältets ingång, för att han må bliva välbehaglig inför HERRENS ansikte.
Och han skall lägga sin hand på brännoffersdjurets huvud; så bliver det välbehagligt, och försoning bringas för honom.
Och han skall slakta ungtjuren inför HERRENS ansikte; och Arons söner, prästerna, skola bära fram blodet, och de skola stänka blodet runt omkring på det altare som står vid ingången till uppenbarelsetältet.
Och han skall draga av huden på brännoffersdjuret och dela det i dess stycken.
Och prästen Arons söner skola göra upp eld på altaret och lägga ved på elden.
Och Arons söner, prästerna, skola lägga styckena, huvudet och istret ovanpå veden som ligger på altarets eld.
Men inälvorna och fötterna skola tvås i vatten.
Och prästen skall förbränna alltsammans på altaret: ett brännoffer, ett eldsoffer till en välbehaglig lukt för HERREN.
Men om han vill bära fram ett brännoffer av småboskapen, vare sig av fåren eller av getterna, så skall han därtill taga ett felfritt djur av hankön.
Och han skall slakta det vid sidan av altaret, norrut, inför HERRENS ansikte, och Arons söner, prästerna, skola stänka dess blod på altaret runt omkring.
Och han skall dela det i dess stycken och frånskilja dess huvud och ister; och prästen skall lägga detta ovanpå veden som ligger på altarets eld.
Men inälvorna och fötterna skola tvås i vatten.
Och prästen skall offra alltsammans och förbränna det på altaret; det är ett brännoffer, ett eldsoffer till en välbehaglig lukt för HERREN.
Men om han vill bära fram åt HERREN ett brännoffer av fåglar, så skall han taga sitt offer av turturduvor eller av unga duvor.
Och prästen skall bära fram djuret till altaret och vrida huvudet av det och förbränna det på altaret.
Och dess blod skall utkramas på altarets vägg.
Men dess kräva med orenligheten däri skall han taga ut, och han skall kasta den vid sidan av altaret, österut, på askhögen.
Och han skall fläka upp det invid vingarna, dock utan att frånskilja dessa; och prästen skall förbränna det på altaret, ovanpå veden som ligger på elden.
Det är ett brännoffer, ett eldsoffer till en välbehaglig lukt för HERREN.
Och när någon vill bära fram ett spisoffer åt HERREN skall hans offer vara av fint mjöl, och han skall gjuta olja därpå och lägga rökelse därpå.
Och han skall bära det fram till Arons söner, prästerna; och prästen skall taga en handfull därav, nämligen av mjölet och oljan, därtill all rökelsen, och skall på altaret förbränna detta, som utgör själva altaroffret: ett eldsoffer till en välbehaglig lukt för HERREN.
Och det som är över av spisoffret skall tillhöra Aron och hans söner.
Bland HERRENS eldsoffer är det högheligt.
Men när du vill bära fram ett spisoffer av det som bakas i ugn, skall det vara av fint mjöl, osyrade kakor, begjutna med olja, och osyrade tunnkakor, smorda med olja.
Och om ditt offer är ett spisoffer som tillredes på plåt, så skall det vara av fint mjöl, begjutet med olja, osyrat.
Du skall bryta sönder det i stycken och gjuta olja därpå.
Det är ett spisoffer.
Och om ditt offer är ett spisoffer som tillredes i panna, så skall det tillredas av fint mjöl med olja.
Det spisoffer som är tillrett på något av dessa sätt skall du föra fram till HERREN; det skall bäras fram till prästen, och han skall hava det fram till altaret.
Och prästen skall av spisoffret taga den del som utgör själva altaroffret och förbränna den på altaret: ett eldsoffer till en välbehaglig lukt för HERREN.
Och det som är över av spisoffret skall tillhöra Aron och hans söner.
Bland HERRENS eldsoffer är det högheligt.
Intet spisoffer som I viljen bära fram åt HERREN skall vara syrat, ty varken av surdeg eller av honung skolen I förbränna något såsom eldsoffer åt HERREN.
Såsom förstlingsoffer mån I bära fram sådant åt HERREN, men på altaret må det icke komma för att vara en välbehaglig lukt.
Och alla dina spisoffer skall du beströ med salt; du må icke låta din Guds förbunds salt fattas på ditt spisoffer.
Till alla dina offer skall du offra salt.
Men om du vill bära fram åt HERREN ett spisoffer av förstlingsfrukter, skall du såsom ett sådant spisoffer av dina förstlingsfrukter böra fram ax, rostade vid eld, sönderstötta, av grönskuren säd.
Och du skall gjuta olja därpå och lägga rökelse därpå.
Det är ett spisoffer.
Och prästen skall förbränna den del av de sönderstötta axen och av oljan, som utgör själva altaroffret, jämte all rökelsen därpå: ett eldsoffer åt Herren.
Och om någon vill bära fram ett tackoffer, och han vill taga sitt offer av fäkreaturen, så skall han ställa fram inför HERRENS ansikte ett felfritt djur, antingen av hankön eller av honkön.
Och han skall lägga sin hand på sitt offerdjurs huvud och sedan slakta det vid ingången till uppenbarelsetältet; och Arons söner, prästerna, skola stänka blodet på altaret runt omkring.
Och av tackoffret skall han såsom eldsoffer åt Herren bära fram det fett som omsluter inälvorna, och allt det fett som sitter på inälvorna,
och båda njurarna med det fett som sitter på dem invid länderna, så ock leverfettet, vilket han skall frånskilja invid njurarna.
Och Arons söner skola förbränna det på altaret, ovanpå brännoffret, på veden som ligger på elden: ett eldsoffer till en välbehaglig lukt för Herren.
Men om någon vill bära fram åt HERREN ett tackoffer av småboskapen, så skall han därtill taga ett felfritt djur, av hankön eller av honkön.
Om det är ett får som han vill offra, så skall han ställa fram det inför HERRENS ansikte.
Och han skall lägga sin hand på sitt offerdjurs huvud och sedan slakta det framför uppenbarelsetältet; och Arons söner skola stänka dess blod på altaret runt omkring.
Och av tackoffersdjuret skall han såsom eldsoffer åt HERREN offra dess fett, hela svansen, frånskild invid ryggraden, och det fett som omsluter inälvorna, och allt det fett som sitter på inälvorna,
och båda njurarna med det fett som sitter på dem invid länderna, så ock leverfettet, vilket han skall frånskilja invid njurarna.
Och prästen skall förbränna det på altaret: en eldsoffersspis åt HERREN.
Likaledes, om någon vill offra en get, så skall han ställa fram denna inför HERRENS ansikte.
Och han skall lägga sin hand på dess huvud och sedan slakta den framför uppenbarelsetältet; och Arons söner skola stänka dess blod på altaret runt omkring.
Och han skall därav såsom eldsoffer åt HERREN offra det fett som omsluter inälvorna, och allt det fett som sitter på inälvorna,
och båda njurarna med det fett som sitter på dem invid länderna, så ock leverfettet, vilket han skall frånskilja invid njurarna.
Och prästen skall förbränna detta på altaret: en eldsoffersspis, till en välbehaglig lukt.
Allt fettet skall tillhöra HERREN.
Detta skall vara en evärdlig stadga för eder från släkte till släkte, var I än ären bosatta: intet fett och intet blod skolen I förtära.
Och HERREN talade till Mose och sade:
Tala till Israels barn och säg: Om någon ouppsåtligen syndar mot något HERRENS bud genom vilket något förbjudes, och han alltså gör något som är förbjudet, så gäller följande:
Om det är den smorde prästen som har syndat och därvid dragit skuld över folket, så skall han för den synd han har begått offra en felfri ungtjur åt HERREN till syndoffer.
Och han skall föra tjuren fram inför HERRENS ansikte, till uppenbarelsetältets ingång.
Och han skall lägga sin hand på tjurens huvud och sedan slakta tjuren inför HERRENS ansikte.
Och den smorde prästen skall taga något av tjurens blod och bära det in i uppenbarelsetältet,
och prästen skall doppa sitt finger i blodet och stänka blodet sju gånger inför HERRENS ansikte, vid förlåten till helgedomen.
Därefter skall prästen med blodet bestryka hornen på den välluktande rökelsens altare, som står inför HERRENS ansikte i uppenbarelsetältet; men allt det övriga blodet av tjuren skall han gjuta ut vid foten av brännoffersaltaret, som står vid ingången till uppenbarelsetältet.
Och allt syndofferstjurens fett skall han taga ut ur honom -- det fett som omsluter inälvorna, och allt det fett som sitter på inälvorna,
och båda njurarna med det fett som sitter på dem invid länderna, så ock leverfettet, vilket han skall frånskilja invid njurarna --
på samma sätt som detta tages ut ur tackofferstjuren; och prästen skall förbränna det på brännoffersaltaret.
Men tjurens hud och allt hans kött jämte hans huvud och hans fötter hans inälvor och hans orenlighet,
korteligen, allt det övriga av tjuren, skall han föra bort utanför lägret till en ren plats, där man slår ut askan, och bränna upp det på ved i eld; på den plats där man slår ut askan skall det brännas upp.
Och om Israels hela menighet begår synd ouppsåtligen, och utan att församlingen märker det, i det att de bryta mot något Herrens bud genom vilket något förbjudes och så ådraga sig skuld,
och den synd de hava begått sedan bliver känd, så skall församlingen offra en ungtjur till syndoffer.
De skola föra honom fram inför uppenbarelsetältet;
och de äldste i menigheten skola lägga sina händer på tjurens huvud inför Herrens ansikte, och sedan skall man slakta tjuren inför HERRENS ansikte.
Och den smorde prästen skall bära något av tjurens blod in i uppenbarelsetältet,
och prästen skall doppa sitt finger i blodet och stänka sju gånger inför HERRENS ansikte, vid förlåten.
Därefter skall han med blodet bestryka hornen på det altare som står inför HERRENS ansikte i uppenbarelsetältet; men allt det övriga blodet skall han gjuta ut vid foten av brännoffersaltaret, som står vid ingången till uppenbarelsetältet.
Och allt tjurens fett skall han taga ut ur honom och förbränna det på altaret.
Så skall han göra med tjuren; såsom han skulle göra med den förra syndofferstjuren, så skall han göra med denna.
När så prästen bringar försoning för dem, då bliver dem förlåtet.
Och han skall föra ut tjuren utanför lägret och bränna upp honom, såsom han skulle göra med den förra tjuren.
Detta är syndoffret för församlingen.
Om en hövding syndar, i det att han ouppsåtligen bryter mot något HERRENS, sin Guds, bud genom vilket något förbjudes, och han själv märker att han har ådragit sig skuld,
eller av någon får veta vilken synd han har begått, så skall han såsom sitt offer föra fram en bock, ett felfritt djur av hankön.
Och han skall lägga sin hand på bockens huvud och sedan slakta honom på samma plats där man slaktar brännoffret, inför HERRENS ansikte.
Det är ett syndoffer.
Och prästen skall taga något av syndoffrets blod på sitt finger och stryka på brännoffersaltarets horn; men det övriga blodet skall han gjuta ut vid foten av brännoffersaltaret.
Och allt fettet skall han förbränna på altaret, såsom det sker med tackoffersdjurets fett.
När så prästen bringar försoning för honom, till rening från hans synd, då bliver honom förlåtet.
Och om någon av det meniga folket syndar ouppsåtligen, därigenom att han bryter mot något HERRENS bud genom vilket något förbjudes, och han själv märker att han har ådragit sig skuld,
eller av någon får veta vilken synd han har begått, så skall han, såsom sitt offer för den synd han har begått, föra fram en felfri get, ett djur av honkön.
Och han skall lägga sin hand på syndoffersdjurets huvud och sedan slakta syndoffersdjuret på den plats där brännoffersdjuren slaktas.
Och prästen skall taga något av blodet på sitt finger och stryka det på brännoffersaltarets horn; men allt det övriga blodet skall han gjuta ut vid foten av altaret.
Och allt fettet skall han taga ut, på samma sätt som fettet tages ut ur tackoffersdjuret, och prästen skall förbränna det på altaret, till en välbehaglig lukt för HERREN.
När så prästen bringar försoning för honom, då bliver honom förlåtet.
Men om någon vill offra ett lamm till syndoffer, så skall han föra fram ett felfritt djur av honkön.
Och han skall lägga sin hand på syndoffersdjurets huvud och sedan slakta det till syndoffer på samma plats där man slaktar brännoffersdjuren.
Och prästen skall taga något av syndoffrets blod på sitt finger och stryka på brännoffersaltarets horn; men allt det övriga blodet skall han gjuta ut vid foten av altaret.
Och allt fettet skall han taga ut, på samma sätt som fettet tages ut ur tackoffersfåret, och prästen skall förbränna det på altaret, ovanpå Herrens eldsoffer.
När så prästen för honom bringar försoning för den synd han har begått, då bliver honom förlåtet.
Och om någon syndar, i det att han, när han hör edsförpliktelsen och kan vittna om något, vare sig han har sett det eller eljest förnummit det, likväl icke yppar detta och han sålunda bär på missgärning;
eller om någon, utan att märka det, kommer vid något orent -- vare sig den döda kroppen av ett orent vilddjur, eller den döda kroppen av ett orent boskapsdjur, eller den döda kroppen av något slags orent smådjur -- och han så bliver oren och ådrager sig skuld;
eller om han, utan att märka det, kommer vid en människas orenhet, det må nu vara vad som helst varigenom hon kan vara oren, och han sedan får veta det och han så ådrager sig skuld;
eller om någon, utan att märka det, svär i obetänksamhet med sina läppar något, vare sig ont eller gott -- det må nu vara vad som helst som man kan svärja i obetänksamhet -- och sedan kommer till insikt därom och han så ådrager sig skuld i något av dessa stycken:
så skall han, när han har ådragit sig skuld i något av dessa stycken, bekänna det vari han har syndat
och såsom bot för den synd han har begått föra fram åt HERREN ett hondjur av småboskapen, antingen en tacka eller en get, till syndoffer.
Och prästen skall bringa försoning för honom, till rening från hans synd.
Men om han icke förmår bekosta ett sådant djur, så skall han såsom bot för vad han har syndat bära fram åt Herren två turturduvor eller två unga duvor, en till syndoffer och en till brännoffer.
Dem skall han bära fram till prästen, och denne skall först offra den som är avsedd till syndoffer.
Han skall vrida huvudet av den invid halsen, dock utan att frånskilja det.
Och han skall stänka något av syndoffrets blod på altarets vägg; men det övriga blodet skall utkramas vid foten av altaret.
Det är ett syndoffer.
Och den andra skall han offra till ett brännoffer, på föreskrivet sätt.
När så prästen bringar försoning för honom, till rening från den synd han har begått, då bliver honom förlåtet.
Men om han icke kan anskaffa två turturduvor eller två unga duvor, så skall han såsom offer för vad han har syndat bära fram en tiondedels efa fint mjöl till syndoffer, men ingen olja skall han gjuta därpå och ingen rökelse lägga därpå, ty det är ett syndoffer.
Och han skall bära det fram till prästen, och prästen skall taga en handfull därav, det som utgör själva altaroffret, och förbränna det på altaret, ovanpå HERRENS eldsoffer.
Det är ett syndoffer.
När så prästen för honom bringar försoning för den synd han har begått i något av dessa stycken, då bliver honom förlåtet.
Och det övriga skall tillhöra prästen, likasom vid spisoffret.
Och HERREN talade till Mose och sade:
Om någon begår en orättrådighet, i det att han ouppsåtligen försyndar sig genom att undanhålla något som är helgat åt Herren, så skall han såsom bot föra fram åt HERREN till skuldoffer av småboskapen en felfri vädur, efter det värde du bestämmer i silver, till ett visst belopp siklar efter helgedomssikelns vikt.
Och han skall giva ersättning för det som han har undanhållit av det helgade och skall lägga femtedelen av värdet därtill; och detta skall han giva åt prästen.
När så prästen bringar försoning för honom genom skuldoffersväduren, då bliver honom förlåtet.
Och om någon, utan att veta det, syndar, i det att han bryter mot något HERRENS bud genom vilket något förbjudes, och han så ådrager sig skuld och bär på missgärning,
så skall han såsom skuldoffer föra fram till prästen av småboskapen en felfri vädur, efter det värde du bestämmer.
När så prästen för honom bringar försoning för den synd han har begått ouppsåtligen och utan att veta det, då bliver honom förlåtet.
Det är ett skuldoffer, ty han har ådragit sig skuld inför HERREN.
Och HERREN talade till Mose och sade:
Om någon syndar och begår en orättrådighet mot HERREN, i det att han inför sin nästa nekar angående något som denne har ombetrott honom eller överlämnat i hans hand, eller angående något som han med våld har tagit; eller i det att han med orätt avhänder sin nästa något;
eller i det att han, när han har hittat något borttappat, nekar därtill och svär falskt i någon sak, vad det nu må vara, vari en människa kan försynda sig:
så skall den som så har syndat Och därmed ådragit sig skuld återställa vad han med våld har tagit eller med orätt tillägnat sig, eller det som har varit honom ombetrott, eller det borttappade som han har hittat,
eller vad det må vara, varom han har svurit falskt; han skall ersätta det till dess fulla belopp och lägga femtedelen av värdet därtill.
Han skall giva det åt ägaren samma dag han bär fram sitt skuldoffer.
Ty sitt skuldoffer skall han föra fram inför HERREN; en felfri vädur av småboskapen, efter det värde du bestämmer, skall han såsom sitt skuldoffer föra fram till prästen.
När så prästen bringar försoning för honom inför HERRENS ansikte, då bliver honom förlåtet, vad han än må hava gjort, som har dragit skuld över honom.
Och Herren talade till Mose och sade:
Bjud Aron och hans söner och säg: Detta är lagen om brännoffret: Brännoffret skall ligga på altarets härd hela natten intill morgonen, och elden på altaret skall därigenom hållas brinnande.
Och prästen skall ikläda sig sin livrock av linne och ikläda sig benkläder av linne, för att de må skyla hans kött; därefter skall han taga bort askan vartill elden har förbränt brännoffret på altaret, och lägga den vid sidan av altaret.
Sedan skall han taga av sig sina kläder och ikläda sig andra kläder och föra askan bort utanför lägret till en ren plats.
Men elden på altaret skall hållas brinnande och får icke slockna; prästen skall var morgon antända ny ved därpå.
Och han skall lägga brännoffret därpå och förbränna fettstyckena av tackoffret därpå.
Elden skall beständigt hållas brinnande på altaret; den får icke slockna.
Och detta är lagen om spisoffret: Arons söner skola bära fram det inför HERRENS ansikte, till altaret.
Och prästen skall taga en handfull därav, nämligen av det fina mjölet som hör till spisoffret, och av oljan, därtill all rökelsen som ligger på spisoffret, och detta, som utgör själva altaroffret, skall han förbränna på altaret, till en välbehaglig lukt för HERREN.
Och det som är över därav skola Aron och hans söner äta.
Osyrat skall det ätas på en helig plats; i förgården till uppenbarelsetältet skola de äta det.
Det skall icke bakas med surdeg.
Detta är deras del, det som jag har givit dem av mina eldsoffer.
Det är högheligt likasom syndoffret och skuldoffret.
Allt mankön bland Arons barn må äta det.
Det skall vara deras evärdliga rätt av HERRENS eldsoffer, från släkte till släkte.
Var och en som kommer därvid bliver helig.
Och HERREN talade till Mose och sade:
Detta är det offer som Aron och hans söner skola offra åt HERREN på den dag då någon av dem undfår smörjelsen: en tiondedels efa fint mjöl såsom det dagliga spisoffret, hälften om morgonen och hälften om aftonen.
På plåt skall det tillredas med olja, och du skall bära fram det hopknådat; och du skall offra det sönderdelat, såsom när man offrar ett spisoffer i stycken, till en välbehaglig lukt för HERREN.
Och den präst bland hans söner, som bliver smord i hans ställe, skall göra så.
Detta skall vara en evärdlig stadga.
Såsom ett heloffer skall det förbrännas åt HERREN.
En prästs spisoffer skall alltid vara ett heloffer; det får icke ätas.
Och HERREN talade till Mose och sade:
Tala till Aron och hans söner och säg: Detta är lagen om syndoffret: På samma plats där brännoffersdjuret slaktas skall ock syndoffersdjuret slaktas, inför HERRENS ansikte.
Det är högheligt.
Den präst som offrar syndoffret skall äta det; på en helig plats skall det ätas, i förgården till uppenbarelsetältet.
Var och en som kommer vid köttet bliver helig.
Och om något av blodet stänkes på någons kläder, så skall man avtvå det bestänkta stället på en helig plats.
Ett lerkärl vari kokningen har skett skall sönderslås; men har kokningen skett i ett kopparkärl, så skall detta skuras och sköljas med vatten.
Allt mankön bland prästerna må äta det.
Det är högheligt.
Men intet syndoffer av vars blod något bäres in i uppenbarelsetältet till att bringa försoning i helgedomen får ätas; det skall brännas upp i eld.
Och detta är lagen om skuldoffret: Det är högheligt.
På samma plats där man slaktar brännoffersdjuret skall man slakta skuldoffersdjuret.
Och man skall stänka dess blod på altaret runt omkring.
Och allt dess fett skall man offra, svansen och det fett som omsluter inälvorna,
och båda njurarna med det fett som sitter på dem invid länderna, så ock leverfettet, vilket man skall frånskilja invid njurarna.
Och prästen skall förbränna det på altaret till ett eldsoffer åt HERREN.
Det är ett skuldoffer.
Allt mankön bland prästerna må äta det; på en helig plats skall det ätas; det är högheligt.
Vad som gäller om syndoffret skall ock gälla om skuldoffret; samma lag skall gälla för dem båda.
Den präst som bringar försoning därmed, honom skall det tillhöra.
Och när en präst bär fram brännoffer for någon, skall huden av det framburna brännoffersdjuret tillhöra den prästen.
Och ett spisoffer som är bakat i ugn, eller som är tillrett i panna eller på plåt, skall alltid tillfalla den präst som bär fram det.
Men ett spisoffer som är begjutet med olja, eller som frambäres torrt, skall alltid tillfalla Arons söner gemensamt, den ene likaväl som den andre.
Och detta är lagen om tackoffret, när ett sådant bäres fram åt HERREN:
Om någon vill bära fram ett sådant till lovoffer, så skall han, förutom det till lovoffret hörande slaktdjuret, bära fram osyrade kakor, begjutna med olja, och osyrade tunnkakor, smorda med olja, och fint mjöl, hopknådat, i form av kakor, begjutna med olja.
Jämte kakor av syrat bröd skall han bära fram detta sitt offer, förutom det slaktdjur som hör till det tackoffer han bär fram såsom lov offer.
Av detta offer skall han bära fram en kaka av vart slag, såsom en gärd åt HERREN; den präst som stänker tackoffrets blod på altaret, honom skall den tillhöra.
Och köttet av det slaktdjur, som hör till det tackoffer som bäres fram såsom lovoffer, skall ätas samma dag det har offrats; intet därav må lämnas kvar till följande morgon.
Om däremot det slaktoffer som någon vill bära fram år ett löftesoffer eller ett frivilligt offer, så skall offerdjuret likaledes ätas samma dag det har offrats; dock må det som har blivit över därav ätas den följande dagen.
Bliver ändå något över av offerköttet, skall detta på tredje dagen brännas upp i eld.
Om någon på tredje dagen äter av tackoffersköttet, så bliver offret icke välbehagligt; honom som har burit fram det skall det då icke räknas till godo, det skall anses såsom en vederstygglighet.
Den som äter därav kommer att bära på missgärning.
Ej heller må det kött ätas, som har kommit vid något orent, utan det skall brännas upp i eld.
För övrigt må köttet ätas av var och en som är ren.
Men den som äter kött av HERRENS tackoffer, medan orenhet låder vid honom, han skall utrotas ur sin släkt.
Och om någon har kommit vid något orent -- vare sig en människas orenhet, eller ett orent djur, eller vilken oren styggelse det vara må -- och han likväl äter kött av HERRENS tackoffer, så skall han utrotas ur sin släkt.
Och HERREN talade till Mose och sade:
Tala till Israels barn och säg: Intet fett av fäkreatur, får eller getter skolen I äta.
Fettet av ett självdött eller ihjälrivet djur må eljest användas till alla slags behov, men äta det skolen I icke.
Ty var och en som äter fettet av något djur varav man bär fram eldsoffer åt HERREN, vem det vara må som äter därav, han skall utrotas ur sin släkt.
Och intet blod skolen I förtära varken av fåglar eller av boskap, var I än ären bosatta.
Var och en som förtär något blod, han skall utrotas ur sin släkt.
Och HERREN talade till Mose och sade:
Tala till Israels barn och säg: Den som vill offra ett tackoffer åt HERREN, han skall av detta sitt tackoffer bära fram åt HERREN den vederbörliga offergåvan.
Med egna händer skall han bära fram HERRENS eldsoffer; fettet jämte bringan skall han bära fram, bringan till att viftas såsom ett viftoffer inför HERRENS ansikte.
Och prästen skall förbränna fettet på altaret, men bringan skall tillhöra Aron och hans söner.
Också det högra lårstycket skolen I giva åt prästen, såsom en gärd av edra tackoffer.
Den bland Arons söner, som offrar tackoffrets blod och fettet, han skall hava det högra lårstycket till sin del.
Ty av Israels barns tackoffer tager jag viftoffersbringan och offergärdslåret och giver dem åt prästen Aron och åt hans söner till en evärdlig rätt av Israels barn.
Detta är Arons och hans söners ämbetslott av HERRENS eldsoffer, den lott som gavs dem den dag de fördes fram till att bliva HERRENS präster
vilken lott, efter HERRENS befallning på den dag då han smorde dem, skulle givas dem av Israels barn, till en evärdlig rätt, släkte efter släkte.
Detta är lagen om brännoffret, spisoffret, syndoffret, skuldoffret, handfyllningsoffret och tackoffret,
vilken HERREN på Sinai berg gav Mose, på den dag då han bjöd Israels barn att de skulle offra sina offer åt HERREN, i Sinais öken.
Och HERREN talade till Mose och sade:
»Tag Aron och hans söner jämte honom samt deras kläder och smörjelseoljan, så ock syndofferstjuren och de två vädurarna och korgen med de osyrade bröden.
Församla sedan hela menigheten vid ingången till uppenbarelsetältet.»
Och Mose gjorde såsom HERREN hade bjudit honom, och menigheten församlade sig vid ingången till uppenbarelsetältet.
Och Mose sade till menigheten: »Detta är vad HERREN har bjudit mig att göra.»
Och Mose förde fram Aron och hans söner och tvådde dem med vatten.
Och han satte livklädnaden på honom och omgjordade honom med bältet och klädde på honom kåpan och satte på honom efoden och omgjordade honom med efodens skärp och fäste därmed ihop alltsammans på honom.
Och han satte på honom bröstskölden och lade urim och tummim in i skölden.
Och han satte huvudbindeln på hans huvud och satte på huvudbindeln framtill den gyllene plåten, det heliga diademet, såsom HERREN hade bjudit Mose.
Och Mose tog smörjelseoljan och smorde tabernaklet och allt vad däri var och helgade allt;
och han stänkte därmed sju gånger på altaret och smorde altaret och alla dess tillbehör och bäckenet jämte dess fotställning, för att helga dem.
Och han göt smörjelseolja på Arons huvud och smorde honom för att helga honom.
Och Mose förde fram Arons söner och satte livklädnader på dem och omgjordade dem med bälten och band huvor på dem, såsom HERREN hade bjudit Mose.
Och han förde fram syndofferstjuren, och Aron och hans söner lade sina händer på syndofferstjurens huvud.
Sedan slaktades den, och Mose tog blodet och strök med sitt finger på altarets horn runt omkring och renade altaret; men det övriga blodet göt han ut vid foten av altaret och helgade detta och bragte försoning för det.
Och han tog allt det fett som satt på inälvorna, så ock leverfettet och båda njurarna med fettet på dem; och Mose förbrände det på altaret.
Men det övriga av tjuren, hans hud och kött och orenlighet, brände han upp i eld utanför lägret såsom HERREN hade bjudit Mose.
Och han förde fram brännoffersväduren, och Aron och hans söner lade sina händer på vädurens huvud.
Sedan slaktades den, och Mose stänkte blodet på altaret runt omkring;
men själva väduren delade han i dess stycken.
Och Mose förbrände huvudet och styckena och istret;
inälvorna och fötterna tvådde han i vatten.
Sedan förbrände Mose hela väduren på altaret.
Det var ett brännoffer till en välbehaglig lukt, det var ett eldsoffer åt HERREN, Såsom HERREN hade bjudit Mose.
Därefter förde han fram den andra väduren, handfyllningsväduren, och Aron och hans söner lade sina händer på vädurens huvud.
Sedan slaktades den, och Mose tog av dess blod och beströk Arons högra örsnibb och tummen på hans högra hand och stortån på hans högra fot.
Därefter förde han fram Arons söner.
Och Mose beströk med blodet deras högra örsnibb och tummen på deras högra hand och stortån på deras högra fot; men det övriga blodet stänkte Mose på altaret runt omkring.
Och han tog fettet, svansen och allt det fett som satt på inälvorna, så ock leverfettet och båda njurarna med fettet på dem, därtill det högra lårstycket.
Och ur korgen med de osyrade bröden, som stod inför HERRENS ansikte, tog han en osyrad kaka, en oljebrödskaka och en tunnkaka och lade detta på fettstyckena och det högra lårstycket.
Och alltsammans lade han på Arons och hans söners händer och viftade det såsom ett viftoffer inför HERRENS ansikte.
Sedan tog Mose det ur deras händer och förbrände det på altaret, ovanpå brännoffret.
Det var ett handfyllningsoffer till en välbehaglig lukt, det var ett eldsoffer åt HERREN.
Och Mose tog bringan och viftade den såsom ett viftoffer inför HERRENS ansikte; av handfyllningsoffrets vädur fick Mose detta till sin del, såsom HERREN hade bjudit Mose.
Och Mose tog av smörjelseoljan och av blodet på altaret och stänkte på Aron -- på hans kläder -- och likaledes på hans söner och hans söners kläder; han helgade så Aron -- hans kläder -- och likaledes hans söner och hans söners kläder.
Och Mose sade till Aron och till hans söner: »Koken köttet vid ingången till uppenbarelsetältet, och äten det där jämte brödet som är i handfyllningskorgen, såsom jag har bjudit och sagt: Aron och hans söner skola äta det.
Men vad som bliver över av köttet; eller av brödet, det skolen I bränna upp i eld.
Och under sju dagar skolen I icke gå bort ifrån uppenbarelsetältets ingång, icke förrän edra handfyllningsdagar äro ute, ty sju dagar skall eder handfyllning vara.
Och HERREN har bjudit, att såsom det i dag har tillgått, så skall det ock sedan tillgå, på det att försoning må bringas för eder.
Vid ingången till uppenbarelsetältet skolen I stanna kvar i sju dygn, dag och natt, och I skolen iakttaga vad HERREN har bjudit eder iakttaga, på det att I icke mån dö; ty så är mig bjudet.»
Och Aron och hans söner gjorde allt vad HERREN hade bjudit genom Mose.
Och på åttonde dagen kallade Mose till sig Aron och hans söner och de äldste i Israel.
Och han sade till Aron: »Tag dig en tjurkalv till syndoffer och en vädur till brännoffer, båda felfria, och för dem fram inför HERRENS ansikte.
Och tala till Israels barn och säg: Tagen en bock till syndoffer och en kalv och ett lamm, båda årsgamla och felfria, till brännoffer,
så ock en tjur och en vädur till tackoffer, att offra inför HERRENS ansikte, därtill ett spisoffer, begjutet med olja; ty i dag uppenbarar sig HERREN för eder.»
Och de togo det som Mose hade givit dem befallning om och förde det fram inför uppenbarelsetältet; och hela menigheten trädde fram och ställde sig inför HERRENS ansikte.
Då sade Mose: »Detta är vad HERREN har bjudit eder göra; så skall HERRENS härlighet visa sig för eder.»
Och Mose sade till Aron: »Träd fram till altaret och offra ditt syndoffer och ditt brännoffer, och bringa försoning för dig själv och folket; offra sedan folkets offer och bringa försoning för dem, såsom HERREN har bjudit.»
Då trädde Aron fram till altaret och slaktade sin syndofferskalv.
Och Arons söner buro fram blodet till honom, och han doppade sitt finger i blodet och strök på altarets horn, men det övriga blodet göt han ut vid foten av altaret.
Och syndoffersdjurets fett, njurar och leverfett förbrände han på altaret, såsom HERREN hade bjudit Mose.
Men köttet och huden brände han upp i eld utanför lägret.
Sedan slaktade han brännoffersdjuret.
Och Arons söner räckte honom blodet, och han stänkte det på altaret runt omkring.
Och de räckte honom brännoffersdjuret, delat i sina stycken, och dess huvud, och han förbrände det på altaret.
Och han tvådde inälvorna och fötterna och förbrände dem ovanpå brännoffret, på altaret.
Därefter förde han fram folkets offer.
Han tog folkets syndoffersbock och slaktade honom och offrade honom till syndoffer, på samma sätt som det förra syndoffersdjuret.
Och han förde fram brännoffersdjuren och offrade dem på föreskrivet sätt.
Och han bar fram spisoffret och tog en handfull därav och förbrände detta på altaret, förutom morgonens brännoffer.
Sedan slaktade han tjuren och väduren, som voro folkets tackoffer.
Och Arons söner räckte honom blodet, och han stänkte det på altaret runt omkring.
Och fettstyckena av tjuren, samt av väduren svansen och vad som omsluter inälvorna, så ock njurarna och leverfettet,
dessa fettstycken lade de på bringorna; och han förbrände fettstyckena på altaret.
Men bringorna och det högra lårstycket viftade Aron till ett viftoffer inför HERRENS ansikte, såsom Mose hade bjudit.
Och Aron lyfte upp sina händer över folket och välsignade det.
Därefter steg han ned, sedan han hade offrat syndoffret, brännoffret och tackoffret.
Och Mose och Aron gingo in i uppenbarelsetältet; sedan gingo de åter ut och välsignade folket.
Då visade sig HERRENS härlighet för allt folket.
Och eld gick ut från HERREN och förtärde brännoffret och fettstyckena på altaret.
Och allt folket såg detta; då jublade de och föllo ned på sina ansikten.
Men Arons söner Nadab och Abihu togo var sitt fyrfat och lade eld i dem och strödde rökelse därpå och buro fram inför HERRENS ansikte främmande eld, annan eld än den han hade givit dem befallning om.
Då gick eld ut från HERREN och förtärde dem, så att de föllo döda ned inför HERRENS ansikte.
Och Mose sade till Aron: »Detta är vad HERREN har talat och sagt: På dem som stå mig nära vill jag bevisa mig helig, och inför allt folket bevisa mig härlig.»
Och Aron teg stilla.
Och Mose kallade till sig Misael och Elsafan, Arons farbroder Ussiels söner, och sade till dem: »Träden fram och bären edra fränder bort ifrån helgedomen och fören den utanför lägret.»
Då trädde de fram och buro bort dem i deras livklädnader, utanför lägret, såsom Mose hade sagt.
Och Mose sade till Aron och till hans söner Eleasar och Itamar: »I skolen icke hava edert hår oordnat, ej heller riva sönder edra kläder, på det att I icke mån dö och draga förtörnelse över hela menigheten.
Men edra bröder, hela Israels hus, må gråta över denna brand som HERREN har upptänt.
Och I skolen icke gå bort ifrån uppenbarelsetältets ingång, på det att I icke mån dö; ty HERRENS smörjelseolja är på eder.»
Och de gjorde såsom Mose hade sagt.
Och HERREN talade till Aron och sade:
»Varken du själv eller dina söner må dricka vin eller starka drycker, när I skolen gå in i uppenbarelsetältet, på det att I icke mån dö.
Det skall vara en evärdlig stadga för eder från släkte till släkte.
I skolen skilja mellan heligt och oheligt, mellan orent och rent;
och I skolen lära Israels barn alla de stadgar som HERREN har kungjort för dem genom Mose.»
Och Mose sade till Aron och till Eleasar och Itamar, hans kvarlevande söner: »Tagen det spisoffer som har blivit över av HERRENS eldsoffer, och äten det osyrat vid sidan av altaret, ty det är högheligt.
I skolen äta det på en helig plats; ty det är din och dina söners stadgade rätt av HERRENS eldsoffer; så är mig bjudet.
Och viftoffersbringan och offergärdslåret skola ätas av dig, och av dina söner och dina döttrar jämte dig, på en ren plats, ty de äro dig givna såsom din och dina söners stadgade rätt av Israels barns tackoffer.
Jämte eldsoffren -- fettstyckena -- skola offergärdslåret och viftoffersbringan bäras fram för att viftas såsom ett viftoffer inför HERRENS ansikte; och de skola såsom en evärdlig rätt tillhöra dig och dina söner jämte dig, såsom HERREN har bjudit.»
Och Mose frågade efter syndoffersbocken, men den befanns vara uppbränd.
Då förtörnades han på Eleasar och Itamar, Arons kvarlevande söner, och sade:
»Varför haven I icke ätit syndoffret på den heliga platsen?
Det är ju högheligt.
Och han har givit eder det, för att I skolen borttaga menighetens missgärning och bringa försoning för dem inför HERRENS ansikte.
Se, dess blod har icke blivit inburet i helgedomens inre; därför skullen I på heligt område hava ätit upp köttet, såsom jag hade bjudit.»
Men Aron sade till Mose: »Se, de hava i dag offrat sitt syndoffer och sitt brännoffer inför HERRENS ansikte, och mig har vederfarits vad du vet.
Om jag nu i dag åte syndofferskött, skulle detta vara HERREN välbehagligt?»
När Mose hörde detta, var han till freds.
Och HERREN talade till Mose och Aron och sade till dem:
Talen till Israels barn och sägen: Dessa äro de djur som I fån äta bland alla fyrfotadjur på jorden:
alla de fyrfotadjur som hava klövar och hava dem helkluvna, och som idissla, dem fån I äta.
Men dessa skolen I icke äta av de idisslande djuren och av dem som hava klövar: kamelen, ty han idisslar väl, men har icke klövar, han skall gälla för eder såsom oren; klippdassen, ty han idisslar väl
men har icke klövar, han skall gälla for eder såsom oren; haren, ty han idisslar väl,
men har icke klövar, han skall gälla för eder såsom oren; svinet,
ty det har väl klövar och har dem helkluvna, men det idisslar icke, det skall gälla för eder såsom orent.
Av dessa djurs kött skolen I icke äta, ej heller skolen I komma vid deras döda kroppar; de skola gälla för eder såsom orena.
Detta är vad I fån äta av allt det som lever i vattnet: allt det i vattnet, vare sig i sjöar eller i strömmar, som har fenor och fjäll, det fån I äta.
Men allt det i sjöar och strömmar, som icke har fenor och fjäll, bland allt det som rör sig i vattnet, bland alla levande varelser i vattnet, det skall vara en styggelse för eder.
Ja, de skola vara en styggelse för eder; av deras kött skolen I icke äta, och deras döda kroppar skolen I räkna såsom en styggelse.
Allt det i vattnet, som icke har fenor och fjäll, skall vara en styggelse för eder.
Och bland fåglarna skolen I räkna dessa såsom en styggelse, de skola icke ätas, de äro en styggelse: örnen, lammgamen, havsörnen,
gladan, falken med dess arter,
alla slags korpar efter deras arter,
strutsen, tahemasfågeln, fiskmåsen, höken med dess arter,
ugglan, dykfågeln, uven,
tinsemetfågeln, pelikanen,
asgamen, hägern, regnpiparen med dess arter, härfågeln och flädermusen.
Alla de flygande smådjur som gå på fyra fötter skola vara en styggelse för eder.
Av alla flygande smådjur, som gå på fyra fötter fån I allenast äta dem som ovanför sina fötter hava två ben att hoppa med på jorden.
Dessa fån I äta bland gräshopporna: arbe med dess arter, soleam med dess arter, hargol med dess arter och hagab med dess arter.
Men alla andra flygande smådjur som hava fyra fötter skola vara en styggelse för eder.
Genom följande djur ådragen I eder orenhet; var och en som kommer vid deras döda kroppar skall vara oren ända till aftonen,
och var och en som har burit bort någon sådan död kropp skall två sina kläder och vara oren ända till aftonen:
alla de fyrfotadjur som hava klövar, men icke helkluvna, och som icke idissla, de skola gälla för eder såsom orena.
Var och en som kommer vid dem bliver oren.
Och alla slags fyrfotade djur som gå på tassar skola gälla för eder såsom orena.
Var och en som kommer vid deras döda kroppar skall vara oren ända till aftonen.
Och den som har burit bort en sådan död kropp, han skall två sina kläder och vara oren ända till aftonen; de skola gälla för eder såsom orena.
Och bland de smådjur som röra sig på jorden skola dessa gälla för eder såsom orena: vesslan, jordråttan, ödlan med dess arter,
anakan, koadjuret, letaan, hometdjuret och kameleonten.
Dessa äro de som skola gälla för eder såsom orena bland alla smådjur.
Var och en som kommer vid dem, sedan de äro döda, skall vara oren ända till aftonen.
Och allt varpå något sådant djur faller, sedan det är dött, bliver orent, vare sig det är något slags träkärl, eller det är kläder, eller något av skinn, eller en säck, eller vilken annan sak det vara må, som användes till något behov.
Man skall lägga det i vatten, och det skall vara orent ända till aftonen; så bliver det rent.
Och om något sådant faller i något slags lerkärl, så bliver allt som är i detta orent, och kärlet skolen I slå sönder.
Allt slags mat däri, allt som man äter tillrett med vatten, det bliver orent; och allt slags dryck i något slags kärl, allt som man dricker, det bliver orent därav.
Och allt varpå någon sådan död kropp faller bliver orent.
Är det en ugn eller en härd, skall den förstöras, ty den bliver oren.
Och den skall gälla för eder såsom oren.
Men en källa eller en brunn, en plats dit vatten samlar sig, skall förbliva ren; men kommer någon vid själva den döda kroppen, bliver han oren.
Och om en sådan död kropp faller på något slags utsädeskorn, något man sår, då förbliver detta rent.
Men om vatten har kommit på säden och någon sådan död kropp sedan faller därpå, så skall den gälla för eder såsom oren.
Och om något fyrfotadjur som får ätas av eder dör, så skall den som kommer vid dess döda kropp vara oren ända till aftonen.
Och den som äter kött av en sådan död kropp, han skall två sina kläder och vara oren ända till aftonen.
Och den som har burit bort någon sådan död kropp, han skall två sina kläder och vara oren ända till aftonen.
Och alla slags smådjur som röra sig på jorden äro en styggelse; de skola icke ätas.
Varken av det som går på buken eller av det som går på fyra eller flera fötter, bland alla de smådjur som röra sig på jorden, skolen I äta något, ty de äro en styggelse.
Gören eder icke själva till en styggelse genom något sådant djur, och ådragen eder icke orenhet genom sådana, så att I bliven orenade genom dem.
Ty jag är HERREN, eder Gud; och I skolen hålla eder heliga och vara heliga, ty jag är helig.
Och I skolen icke ådraga eder orenhet genom något av de smådjur som röra sig på jorden.
Ty jag är HERREN, som har fört eder upp ur Egyptens land, för att jag skall vara eder Gud.
Så skolen I nu vara heliga, ty jag är helig.
Detta är lagen om fyrfotadjuren, och om fåglarna, och om alla slags levande varelser som röra sig i vattnet, och om alla slags smådjur på jorden,
för att man skall kunna skilja mellan orent och rent, mellan de djur som få ätas och de djur som icke få ätas.
Och HERREN talade till Mose och sade:
Tala till Israels barn och säg: När en kvinna föder barn och det är ett gossebarn som hon har fött, så skall hon vara oren i sju dagar; lika många dagar som vid sin månadsrening skall hon vara oren.
Och på åttonde dagen skall barnets förhud omskäras.
Och sedan skall hon stanna hemma trettiotre dagar, under sitt reningsflöde.
Hon skall icke komma vid något heligt och får icke heller komma till helgedomen, förrän hennes reningsdagar äro ute.
Men om det är ett flickebarn som hon har fött, så skall hon vara oren i två veckor, på samma sätt som vid sin månadsrening; och sedan skall hon stanna hemma i sextiosex dagar, under sitt reningsflöde.
Och när hennes reningsdagar äro ute, vare sig efter son eller efter dotter, skall hon föra fram ett årsgammalt lamm såsom brännoffer, och en ung duva eller en turturduva såsom syndoffer, till uppenbarelsetältets ingång, till prästen.
Och han skall offra detta inför HERRENS ansikte och bringa försoning för henne, så bliver hon ren från sitt blodflöde.
Detta är lagen om en barnaföderska, när hon har fött ett gossebarn, och när hon har fött ett flickebarn.
Och om hon icke förmår bekosta ett får, så skall hon taga två turturduvor eller två unga duvor, en till brännoffer och en till syndoffer.
Och prästen skall bringa försoning för henne, så bliver hon ren.
Och HERREN talade till Mose och Aron och sade:
När någon på sin kropps hud får en upphöjning eller ett utslag eller en ljus fläck, och därav uppstår ett spetälskeartat ont på hans kropps hud, så skall han föras till prästen Aron eller till en av hans söner, prästerna.
Om då prästen, när han beser det angripna stället på hans kropps hud, finner att håret på det angripna stället har vitnat, och att det angripna stället visar sig djupare än den övriga huden på kroppen, så är han angripen av spetälska; och sedan prästen har besett honom skall han förklara honom oren.
Och om det är en vit fläck som synes på hans kropps hud, men den icke visar sig djupare än den övriga huden, och håret därpå icke har vitnat, så skall prästen hålla den angripne innestängd i sju dagar.
Om då prästen, när han på sjunde dagen beser honom, finner att det angripna stället visar sig oförändrat, och att det onda icke har utbrett sig på huden, så skall prästen för andra gången hålla honom innestängd i sju dagar.
Om då prästen, när han på sjunde dagen beser honom för andra gången, finner att det angripna stället har bleknat, och att det onda icke har utbrett sig på huden, så skall prästen förklara honom ren, ty då är det ett vanligt utslag, och sedan han har tvått sina kläder, är han ren.
Men om utslaget utbreder sig på huden, sedan han har låtit bese sig av prästen för att förklaras ren, och han nu för andra gången låter bese sig av prästen
och prästen då, när han beser honom, finner att utslaget har utbrett sig på huden, så skall prästen förklara honom oren, ty då är det spetälska.
När någon bliver angripen av spetälska, skall han föras till prästen.
Om då prästen, när han beser honom, finner en vit upphöjning på huden, och ser att håret där har vitnat, och att svallkött bildar sig i upphöjningen,
så är det gammal spetälska på hans kropps hud, och prästen skall förklara honom oren; han skall då icke stänga honom inne, ty han är oren.
Men om spetälskan så har brutit ut på huden, att på den angripne hela huden, från huvud till fötter, överallt där prästen ser, är betäckt av spetälska
och prästen alltså, när han beser honom, finner att spetälska betäcker hela hans kropp, så skall han förklara den angripne ren.
Hela hans kropp har blivit vit; han är ren.
Men så snart svallkött visar sig på honom, är han oren.
När prästen ser svallköttet, skall han förklara honom oren; svallköttet är orent, det är spetälska.
Men om svallköttet förändrar sig och stället bliver vitt, så skall han komma till prästen.
Om då prästen, när han beser honom, finner att det angripna stället har blivit vitt, så skall prästen förklara den angripne ren, han är då ren.
När någon på sin kropps hud har haft en bulnad som har blivit läkt,
men sedan, på det ställe där bulnaden var, en vit upphöjning eller en rödvit fläck visar sig, så skall han låta bese sig av prästen.
Om då prästen, när han beser honom, finner att stället visar sig lägre än den övriga huden, och att håret därpå har vitnat, så skall prästen förklara honom oren; ty då är han angripen av spetälska, som har brutit ut där bulnaden var.
Men om prästen, när han beser stället, finner att vitt hår saknas där, och att stället icke är lägre än den övriga huden, och att det är blekt, så skall prästen hålla honom innestängd i sju dagar.
Om då det onda utbreder sig på huden, så skall prästen förklara honom oren, ty då är han angripen.
Men om den ljusa fläcken bliver oförändrad där den är och icke utbreder sig, då är det ett märke efter bulnaden, och prästen skall förklara honom ren.
Men om någon på sin kropps hud får ett brännsår, och om av ärrbildningen i brännsåret sedan bliver en rödvit eller vit fläck
och prästen, när han beser stället, finner att håret på fläcken har vitnat, och att den visar sig djupare än den övriga huden, så är mannen angripen av spetälska, som har brutit ut där brännsåret var; och prästen skall förklara honom oren, ty då är han angripen av spetälska.
Men om prästen, när han beser stället, finner att vitt hår saknas på den ljusa fläcken, och att stället icke är lägre än den övriga huden, och att det är blekt, så skall prästen hålla honom innestängd i sju dagar.
Om då prästen, när han på sjunde dagen beser honom, finner att det onda har utbrett sig på huden, så skall prästen förklara honom oren ty då är han angripen av spetälska.
Men om den ljusa fläcken bliver oförändrad där den är och icke utbreder sig på huden och förbliver blek, då är det en upphöjning efter brännsåret, och prästen skall förklara honom ren, ty det är ett märke efter brännsåret.
När på en man eller en kvinna något ställe på huvudet eller på hakan bliver angripet
och prästen, då han beser det angripna stället, finner att det visar sig djupare än den övriga huden och att gulaktigt tunt hår finnes där, så skall prästen förklara den angripne oren, ty då är det spetälskeskorv, huvud- eller hakspetälska.
Men om prästen, när han beser det angripna stället med skorven, finner, att om det än icke visar sig djupare än den övriga huden, svart hår likväl saknas där, så skall prästen hålla den av skorven angripne innestängd i sju dagar.
Om då prästen, när han på sjunde dagen beser det angripna stället, finner att skorven icke har utbrett sig, och att där icke finnes något gulaktigt hår, och att skorven icke visar sig djupare än den övriga huden,
så skall den sjuke raka sig, utan att dock raka det skorviga stället, och prästen skall för andra gången hålla den skorvsjuke innestängd i sju dagar.
Om då prästen, när han på sjunde dagen beser den skorvsjuke, finner att skorven icke har utbrett sig på huden, och att den icke visar sig djupare än den övriga huden, så skall prästen förklara honom ren, och sedan han har tvått sina kläder, är han ren.
Men om skorven utbreder sig på huden, sedan han har blivit förklarad ren,
och prästen, när han beser honom, finner att skorven har utbrett sig på huden, så behöver prästen icke efterforska om där finnes något gulaktigt hår, ty han är oren.
Men om skorven visar sig oförändrad, och svart hår har vuxit upp på stället, då är skorven läkt, och han är ren, och prästen skall förklara honom ren.
När någon, man eller kvinna, på sin kropps hud får fläckar, vita fläckar,
och prästen, när han beser den angripne, finner att fläckarna på hans kropps hud äro blekvita, då är det ett ofarligt utslag som har kommit fram på huden; han är ren.
När på en mans huvud håret utan vidare faller av, är det vanlig bakskallighet; han är ren.
Och om håret utan vidare faller av på främre delen av huvudet, så är det vanlig framskallighet; han är ren.
Men när på det skalliga stället, baktill eller framtill, en rödvit fläck uppstår, då är det spetälska som har brutit ut på det skalliga stället baktill eller framtill.
Om alltså prästen, när han beser honom, finner att den upphöjda fläcken på det skalliga stället, baktill eller framtill, är rödvit, och att den visar sig lik spetälska på den övriga kroppens hud,
så är mannen spetälsk, han är oren; prästen skall strax förklara honom oren, ty han är angripen på sitt huvud.
Den som är angripen av spetälska skall gå med sönderrivna kläder, han skall hava sitt hår oordnat och skyla sitt skägg, och han skall ropa: »Oren!
Oren!»
Så länge han är angripen av spetälska, skall han vara oren; oren är han.
Han skall bo avskild; utanför lägret skall han hava sin bostad.
När en klädnad bliver angripen av spetälska, vare sig klädnaden är av ylle eller av linne,
eller när så sker med något vävt eller virkat tyg, vare sig av linne eller av ylle, eller med skinn eller med något, vad det vara må, som är förfärdigat av skinn,
och det angripna stället visar sig grönaktigt eller rödaktigt, på klädnaden eller skinnet, eller på det vävda eller virkade tyget, eller på skinnsaken, vad det vara må, då är stället angripet av spetälska och skall visas för prästen.
Och när prästen har besett det angripna stället, skall han hava den angripna saken inlåst i sju dagar.
Om han då, när han på sjunde dagen beser det angripna stället, finner att skadan har utbrett sig på klädnaden, eller på det vävda eller virkade tyget, eller på skinnet, vadhelst det vara må, som är förfärdigat av skinnet, så är stället angripet av elakartad spetälska; sådant är orent.
Och man skall bränna upp klädnaden, eller det vävda eller virkade tyget, vare sig det år av ylle eller av linne, eller skinnsaken som är angripen, vad det vara må; ty det är en elakartad spetälska; allt sådant skall brännas upp i eld.
Men om prästen, när han beser stället, finner att fläcken icke har utbrett sig på klädnaden, eller på det vävda eller virkade tyget, eller på skinnsaken, vad det vara må,
så skall prästen bjuda att man tvår den sak på vilken det angripna stället finnes, och han skall för andra gången hava den inlåst i sju dagar.
Om då prästen, när han efter tvagningen beser det angripna stället, finner att det angripna stället icke har förändrat sitt utseende, så är en sådan sak oren, om ock fläcken icke vidare har utbrett sig; du skall bränna upp den i eld; det är en frätfläck, vare sig den sitter på avigsidan eller på rätsidan.
Men om prästen, när han beser det angripna stället, finner att det efter tvagningen har bleknat, så skall han riva bort det från klädnaden eller skinnet, eller från det vävda eller virkade tyget.
Om likväl sedan en fläck åter visar sig på klädnaden, eller på det vävda eller virkade tyget, eller på skinnsaken, vad det vara må, så är det spetälska som har brutit ut; den sak på vilken det angripna stället finnes skall du bränna upp i eld.
Men om genom tvagningen fläcken har gått bort på klädnaden, eller på det vävda eller virkade tyget, eller på skinnsaken, vad det vara må, så skall det för andra gången tvås, och så bliver det rent.
Detta är lagen om det som bliver angripet av spetälska, antingen det är en klädnad av ylle eller linne, eller det är vävt eller virkat tyg, eller någon skinnsak, vad det vara må -- den lag efter vilken det skall förklaras rent eller orent.
Och HERREN talade till Mose och sade:
Detta vare lagen om huru man skall förfara, när den som har haft spetälska skall renas: Han skall föras till prästen;
och prästen skall gå ut utanför lägret.
Om då prästen, när han beser den spetälske, finner att han är botad från den spetälska varav han var angripen,
så skall prästen bjuda att man för dens räkning, som skall renas, tager två levande rena fåglar, cederträ, rosenrött garn och isop.
Och prästen skall bjuda att man slaktar den ena fågeln över ett lerkärl med friskt vatten i.
Sedan skall han taga den levande fågeln, så ock cederträet, det rosenröda garnet och isopen, och detta alltsammans, jämväl den levande fågeln, skall han doppa i den fågelns blod, som har blivit slaktad över det friska vattnet.
Och han skall stänka sju gånger på den som skall renas från spetälskan; och sedan han så har renat honom, skall han slappa den levande fågeln fri ute på marken.
Och den som skall renas skall två sina kläder och raka av allt sitt hår och bada sig i vatten, så bliver han ren och får sedan gå in i lägret.
Dock skall han stanna utanför sitt tält i sju dagar.
Och på sjunde dagen skall han raka av allt sitt hår, både huvudhåret och skägget och ögonbrynen: allt sitt hår skall han raka av.
Och han skall två sina kläder och bada sin kropp i vatten, så bliver han ren.
Och på åttonde dagen skall han taga två felfria lamm av hankön och ett årsgammalt felfritt lamm av honkön, så ock tre tiondedels efa fint mjöl, begjutet med olja, till spisoffer, och därtill en log olja.
Och prästen som förrättar reningen skall ställa den som skall renas och allt det andra fram inför HERRENS ansikte, vid ingången till uppenbarelsetältet.
Och prästen skall taga det ena lammet och offra det till ett skuldoffer, jämte tillhörande log olja, och vifta detta såsom ett viftoffer inför HERRENS ansikte.
Och man skall slakta lammet på samma plats där man slaktar synd- och brännoffersdjuren, på en helig plats; ty skuldoffret tillhör prästen, likasom syndoffret; det är högheligt.
Och prästen skall taga något av skuldoffrets blod, och därmed skall prästen bestryka högra örsnibben på den som skall renas, så ock tummen på hans högra hand och stortån på hans högra fot.
Sedan skall prästen taga av tillhörande log olja och gjuta i sin vänstra hand,
och prästen skall doppa sitt högra pekfinger i oljan som han har i sin vänstra hand och stänka något av oljan med sitt finger sju gånger inför HERRENS ansikte.
Och med det som bliver över av oljan i hans hand skall prästen bestryka högra örsnibben på den som skall renas, så ock tummen på hans högra hand och stortån på hans högra fot, ovanpå skuldoffersblodet.
Och det som sedan är över av oljan i prästens hand skall han gjuta på dens huvud, som skall renas; så skall prästen bringa försoning för honom inför HERRENS ansikte.
Därefter skall prästen offra syndoffret och bringa försoning för den som skall renas, så att han bliver fri ifrån sin orenhet; sedan skall han slakta brännoffersdjuret.
Och prästen skall offra brännoffret på altaret och tillika spisoffret.
När så prästen bringar försoning för honom, då bliver han ren.
Men om han är fattig och icke kan anskaffa så mycket, så skall han taga allenast ett lamm till skuldoffer, och vifta det för att bringa försoning för sig, och allenast en tiondedels efa fint mjöl, begjutet med olja, till spisoffer, och därtill en log olja,
så ock två turturduvor eller två unga duvor, efter som han kan anskaffa; den ena skall vara till syndoffer, den andra till brännoffer.
Och han skall, för att förklaras ren, bära allt detta till prästen på åttonde dagen, till uppenbarelsetältets ingång, inför HERRENS ansikte.
Och prästen skall taga skuldofferslammet och tillhörande log olja, och detta skall prästen vifta såsom ett viftoffer inför HERRENS ansikte.
Och man skall slakta skuldofferslammet, och prästen skall taga av skuldoffrets blod och bestryka högra örsnibben på den som skall renas, så ock tummen på hans högra hand och stortån på hans högra fot.
Sedan skall prästen gjuta något av oljan i sin vänstra hand,
och prästen skall stänka med sitt högra pekfinger något av oljan som han har i sin vänstra hand sju gånger inför HERRENS ansikte.
Och prästen skall med oljan som han har i sin hand bestryka högra örsnibben på den som skall renas, så ock tummen på hans högra hand och stortån på hans högra fot, ovanpå skuldoffersblodet.
Och det som är över av oljan i prästens hand skall han gjuta på dens huvud, som skall renas, till att bringa försoning för honom inför HERRENS ansikte.
Därefter skall han offra den ena av turturduvorna eller av de unga duvorna, vad han nu har kunnat anskaffa;
efter som han har kunnat anskaffa: skall han offra den ena till syndoffer och den andra till brännoffer, tillika med spisoffret.
Så skall prästen bringa försoning inför HERRENS ansikte för den som skall renas.
Detta är lagen om den som har varit angripen av spetälska, men icke kan anskaffa vad som rätteligen hör till hans rening.
Och HERREN talade till Mose och Aron och sade:
När I kommen in i Kanaans land, som jag vill giva eder till besittning, och jag låter något hus i det land I fån till besittning bliva angripet av spetälska,
så skall husets ägare gå och anmäla det för prästen och säga: »Det synes som om mitt hus vore angripet av spetälska.»
Då skall prästen bjuda att man, innan prästen går in för att bese det angripna stället, utrymmer huset, för att icke allt som är i huset skall bliva orent.
Och därefter skall prästen gå in för att bese huset.
Om han då, när han beser det angripna stället, finner att det angripna stället på husets vägg bildar grönaktiga eller rödaktiga fördjupningar, som visa sig lägre än den övriga väggen,
så skall prästen gå ut ur huset, till dörren på huset, och stänga huset för sju dagar.
Om då prästen, när han på sjunde dagen kommer igen och beser det, finner att fläcken har utbrett sig på husets vägg,
så skall prästen bjuda att man bryter ut de stenar som äro angripna, och kastar dem utanför staden på någon oren plats.
Men huset skall man skrapa överallt innantill och kasta det avskrapade murbruket utanför staden på någon oren plats.
Och man skall taga andra stenar och sätta in dem i de förras ställe och taga annat murbruk och rappa huset därmed.
Om likväl en fläck åter kommer fram på huset, sedan man har brutit ut stenarna, och sedan man har skrapat huset, och sedan det har blivit rappat,
så skall prästen gå in och bese det, och om han då finner att fläcken har utbrett sig på huset, så är detta en elakartad spetälska på huset, det är orent.
Och man skall riva ned huset, med dess stenar och trävirke och allt murbruk på huset, och föra bort alltsammans utanför staden till någon oren plats.
Och om någon har gått in i huset under den tid det skulle vara stängt, så skall han vara oren ända till aftonen.
Och om någon har legat i huset, skall han två sina kläder, och om någon har ätit i huset, skall också han två sina kläder.
Men om prästen, när han går in och beser huset, finner att fläcken icke har utbrett sig på huset, sedan det har blivit rappat, så skall han förklara huset rent, ty då är det onda hävt.
Och han skall till husets rening taga två fåglar, cederträ, rosenrött garn och isop.
Och han skall slakta den ena fågeln över ett lerkärl med friskt vatten i.
Sedan skall han taga cederträet, isopen, det rosenröda garnet och den levande fågeln, och doppa alltsammans i den slaktade fågelns blod och det friska vattnet, och stänka på huset sju gånger.
Så skall han rena huset med fågelns blod och det friska vattnet och med den levande fågeln, cederträet, isopen och det rosenröda garnet.
Och han skall släppa den levande fågeln fri ute på marken utanför staden.
När han så bringar försoning för huset, då bliver det rent.
Detta är lagen om allt slags spetälskesjukdom och spetälskeskorv,
om spetälska på kläder och på hus,
om upphöjningar på huden, utslag och ljusa fläckar,
till undervisning om när något är orent eller rent.
Detta är lagen om spetälska.
Och HERREN talade till Mose och Aron och sade:
Talen till Israels barn och sägen till dem:
Om någon får flytning ur sitt kött, så är sådan flytning oren.
Och angående hans orenhet, medan flytningen varar, gäller följande: Evad hans kött avsöndrar flytningen, eller det tillsluter sig för flytningen, så är han oren.
Allt varpå den sjuke ligger bliver orent, och allt varpå han sitter bliver orent.
Och den som kommer vid det varpå han har legat skall två sina kläder och bada sig i vatten och vara oren ända till aftonen.
Och den som sätter sig på något varpå den sjuke har suttit skall två sina kläder och bada sig i vatten och vara oren ända till aftonen.
Och den som kommer vid den sjukes kropp skall två sina kläder och bada sig i vatten och vara oren ända till aftonen.
Och om den sjuke spottar på någon som är ren, skall denne två sina kläder och bada sig i vatten och vara oren ända till aftonen.
Och allt varpå den sjuke sitter när han färdas någonstädes, bliver orent.
Och var och en som kommer vid något, vad det vara må, som har legat under honom skall vara oren ända till aftonen; och den som bär bort något sådant skall två sina kläder och bada sig i vatten och vara oren ända till aftonen.
Och var och en som den sjuke kommer vid, utan att hava sköljt sina händer i vatten, skall två sina kläder och bada sig i vatten och vara oren ända till aftonen.
Och ett lerkärl som den sjuke kommer vid skall sönderslås; men är det ett träkärl, skall det sköljas med vatten.
När den som har flytning bliver ren från sin flytning, skall han, för att förklaras ren, räkna sju dagar och därefter två sina kläder, och sedan skall han bada sin kropp i rinnande vatten, så bliver han ren.
Och på åttonde dagen skall han taga sig två turturduvor eller två unga duvor och komma inför HERRENS ansikte, till uppenbarelsetältets ingång, och giva dem åt prästen.
Och prästen skall offra dem, den ena till syndoffer och den andra till brännoffer; så skall prästen bringa försoning för honom inför HERRENS ansikte, till rening från hans flytning.
Och om en man har haft sädesutgjutning, så skall han bada hela sin kropp i vatten och vara oren ända till aftonen.
Och allt slags klädnad och allt av skinn, varpå sådan sädesutgjutning har skett, skall tvås i vatten och vara orent ända till aftonen.
Och när en man har legat hos en kvinna och sädesutgjutning har skett, så skola de båda bada sig i vatten och vara orena ända till aftonen.
Och när en kvinna har sin flytning, i det att blod avgår ur hennes kött, skall hon vara oren i sju dagar, och var och en som kommer vid henne skall vara oren ända till aftonen.
Och allt varpå hon ligger under sin månadsrening bliver orent, och allt varpå hon sitter bliver orent.
Och var och en som kommer vid det varpå hon har legat skall två sina kläder och bada sig i vatten och vara oren ända till aftonen.
Och var och en som kommer vid något varpå hon har suttit skall två sina kläder och bada sig i vatten och vara oren ända till aftonen.
Och om någon sak lägges på det varpå hon har legat eller suttit, och någon då kommer vid denna sak, så skall han vara oren ända till aftonen.
Och om en man ligger hos henne, och något av hennes månadsflöde kommer på honom, skall han vara oren i sju dagar, och allt varpå han ligger bliver orent.
Och om en kvinna har blodflöde under en längre tid, utan att det är hennes månadsrening, eller om hon har flöde utöver tiden för sin månadsrening, så skall om henne, så länge hennes orena flöde varar, gälla detsamma som under hennes månadsreningstid; hon är oren.
Om allt varpå hon ligger, så länge hennes flöde varar, skall gälla detsamma som om det varpå hon ligger under sin månadsrening; och allt varpå hon sitter bliver orent, likasom under hennes månadsrening.
Och var och en som kommer vid något av detta bliver oren; han skall två sina kläder och bada sig i vatten och vara oren ända till aftonen.
Men om hon bliver ren från sitt flöde, skall hon räkna sju dagar och sedan vara ren.
Och på åttonde dagen skall hon taga sig två turturduvor eller två unga duvor och bära dem till prästen, till uppenbarelsetältets ingång.
Och prästen skall offra den ena till syndoffer och den andra till brännoffer; så skall prästen bringa försoning för henne inför HERRENS ansikte, till rening från hennes orena flöde.
Så skolen I bevara Israels barn från orenhet, på det att de icke må dö i sin orenhet, om de orena mitt tabernakel, som står mitt ibland dem.
Detta är lagen om den som har flytning och om den som har sädesutgjutning, så att han därigenom bliver oren,
och om den kvinna som har sin månadsrening, och om den som har någon flytning, evad det är man eller kvinna, så ock om en man som ligger hos en oren kvinna.
Och HERREN talade till Mose, sedan Arons två söner voro döda, de båda som träffats av döden, när de trädde fram inför HERRENS ansikte.
Och HERREN sade till Mose: Säg till din broder Aron att han icke på vilken tid som helst får gå in i helgedomen innanför förlåten, framför nådastolen som är ovanpå arken, på det att han icke må dö; ty i molnskyn vill jag uppenbara mig över nådastolen.
Så skall förfaras, när Aron skall gå in i helgedomen: Han skall taga en ungtjur till syndoffer och en vädur till brännoffer;
han skall ikläda sig en helig livklädnad av linne och hava benkläder av linne över sitt kött, och han skall omgjorda sig med ett bälte av linne och vira en huvudbindel av linne om sitt huvud; detta är de heliga kläderna, och innan han ikläder sig dem, skall han bada sin kropp i vatten.
Och av Israels barns menighet skall han mottaga två bockar till syndoffer och en vädur till brännoffer.
Och Aron skall föra fram sin egen syndofferstjur och bringa försoning för sig och sitt hus.
Sedan skall han taga de två bockarna och ställa dem inför HERRENS ansikte, vid ingången till uppenbarelsetältet.
Och Aron skall draga lott om de två bockarna: en lott för HERREN och en lott för Asasel.
Och den bock som lotten bestämmer åt HERREN skall Aron föra fram och offra till syndoffer.
Men den bock som lotten bestämmer åt Asasel skall ställas levande inför HERRENS ansikte, för att försoning må bringas för honom, på det att han må släppas fri ut till Asasel i öknen.
Aron skall alltså föra fram sin syndofferstjur och bringa försoning för sig och sitt hus, han skall slakta sin syndofferstjur.
Sedan skall han taga ett fyrfat fullt med glöd från altaret som står inför HERRENS ansikte, och fylla sina händer med stött välluktande rökelse; och han skall bära in detta innanför förlåten.
Och rökelsen skall han lägga på elden inför HERRENS ansikte, så att ett moln av rökelse skyler nådastolen, ovanpå vittnesbördet, på det att han icke må dö.
Och han skall taga av tjurens blod och stänka med sitt finger framtill på nådastolen; och framför nådastolen skall han stänka blodet sju gånger med sitt finger.
Sedan skall han slakta folkets syndoffersbock och bära in hans blod innanför förlåten; och han skall göra med hans blod såsom han gjorde med tjurens blod: han skall tänka därmed på nådastolen och framför nådastolen.
Så skall han bringa försoning för helgedomen och rena den från Israels barns orenheter och överträdelser, vad de än må hava syndat.
Och på samma sätt skall han göra ned uppenbarelsetältet, som har sin plats hos dem mitt ibland deras orenheter.
Och ingen människa får vara i uppenbarelsetältet, från den stund på han går in för att bringa försoning i helgedomen, ända till dess han har gått ut.
Så skall han bringa försoning för sig och sitt hus och för Israels hela församling.
Sedan skall han gå ut till altaret som står inför HERRENS ansikte och bringa försoning för det; han skall taga av tjurens blod och av bockens blod och stryka på altarets horn runt omkring,
och han skall stänka blodet därpå med sitt finger sju gånger, och rena och helga det från Israels barns orenheter.
När han så har fullbordat försoningen för helgedomen, uppenbarelsetältet och altaret, skall han föra fram den levande bocken.
Och Aron skall lägga båda sina händer på den levande bockens huvud, och bekänna över honom Israels barns alla missgärningar och alla deras överträdelser, vad de än må hava syndat; han skall lägga dem på bockens huvud och genom en man som hålles redo därtill släppa honom ut i öknen.
Så skall bocken bära alla deras missgärningar på sig ut i vildmarken; man skall släppa bocken ute i öknen.
Därefter skall Aron gå in i uppenbarelsetältet och taga av sig linnekläderna, som han hade iklätt sig när han gick in i helgedomen; och han skall lämna dem där.
Och han skall bada sin kropp i vatten på en helig plats och ikläda sig sina vanliga kläder; sedan skall han gå ut och offra sitt eget brännoffer och folkets brännoffer och bringa försoning för sig och för folket.
Och fettet av syndoffersdjuret skall han förbränna på altaret.
Men den som släppte bocken ut till Asasel skall två sina kläder och bada sin kropp i vatten; därefter får han gå in i lägret.
Och syndofferstjuren och syndoffersbocken, vilkas blod blev inburet för att bringa försoning i helgedomen, skola föras bort utanför lägret, och man skall bränna upp dem i eld med deras hud och kött och orenlighet.
Och den som bränner upp detta skall två sina kläder och bada sin kropp i vatten; därefter får han gå in i lägret.
Och detta skall vara för eder en evärdlig stadga: I sjunde månaden, på tionde dagen i månaden, skolen I späka eder och icke göra något arbete, varken infödingen eller främlingen som bor ibland eder.
Ty på den dagen skall försoning bringas för eder, till att rena eder; från alla edra synder skolen I renas inför HERRENS ansikte.
En vilosabbat skall den vara för eder, och I skolen då späka eder.
Detta skall vara en evärdlig stadga.
Och den präst, som har blivit smord och mottagit handfyllning till att vara präst i sin faders ställe skall bringa denna försoning; han skall ikläda sig linnekläderna, de heliga kläderna,
och han skall bringa försoning för det allraheligaste och försoning för uppenbarelsetältet och altaret, och han skall bringa försoning för prästerna och allt folket i församlingen.
Detta skall vara för eder en evärdlig stadga, att försoning skall bringas för Israels barn, till rening från alla deras synder, en gång om året.
Och han gjorde såsom HERREN hade bjudit Mose.
Och HERREN talade till Mose och sade:
Tala till Aron och hans söner och alla Israels barn och säg till dem Detta är vad HERREN har bjudit och sagt:
Om någon av Israels hus, i lägret eller utanför lägret, slaktar ett fäkreatur eller ett lamm eller en get,
utan att föra fram djuret till uppenbarelsetältets ingång för att frambära det såsom en offergåva åt HERREN framför HERRENS tabernakel, så skall detta tillräknas den mannen såsom blodskuld, ty blod har han utgjutit, och den mannen skall utrotas ur sitt folk.
Därför skola Israels barn föra sina slaktdjur, som de pläga slakta ute på marken, fram till HERREN, till uppenbarelsetältets ingång, till prästen, och där slakta dem såsom tackoffer åt HERREN.
Och prästen skall stänka blodet på HERRENS altare, vid ingången till uppenbarelsetältet, och förbränna fettet till en välbehaglig lukt för HERREN.
Och de skola icke mer offra sina slaktoffer åt de onda andar som de i trolös avfällighet löpa efter.
Detta skall vara en evärdlig stadga för dem från släkte till släkte.
Och du skall säga till dem: Om någon av Israels hus, eller av främlingarna som bo ibland dem, offrar ett brännoffer eller ett slaktoffer
och icke för det fram till uppenbarelsetältets ingång för att offra det åt HERREN, så skall den mannen utrotas ur sin släkt.
Och om någon av Israels hus, eller av främlingarna som bo ibland dem, förtär något blod, så skall jag vända mitt ansikte mot honom som förtär blodet och utrota honom ur hans folk.
Ty allt kötts själ är i blodet, och jag har givit eder det till altaret, till att bringa försoning för edra själar; ty blodet är det som bringar försoning, genom själen som är däri.
Därför säger jag till Israels barn: Ingen av eder skall förtära blod; och främlingen som bor ibland eder skall icke heller förtära blod.
Och om någon av Israels barn, eller av främlingarna som bo ibland dem, fäller ett villebråd av fyrfotadjur eller en fågel, sådant som får ätas, så skall han låta blodet rinna ut och övertäcka det med jord.
Ty så är det med allt kötts själ, att blodet är det som innehåller själen; därför säger jag till Israels barn: I skolen icke förtära något kötts blod.
Ty blodet är allt kötts själ; var och en som förtär det skall utrotas.
Och var och en som äter ett självdött eller ihjälrivet djur, evad han är inföding eller främling, skall två sina kläder och bada sig i vatten och vara oren ända till aftonen; då bliver han ren.
Men om han icke tvår sina kläder och icke badar sin kropp kommer han att bära på missgärning.
Och HERREN talade till Mose och sade:
Tala till Israels barn och säg till dem: Jag är HERREN, eder Gud.
I skolen icke göra såsom man gör i Egyptens land, där I haven bott.
Ej heller skolen I göra såsom man gör i Kanaans land, dit jag vill föra eder; I skolen icke vandra efter deras stadgar.
Efter mina rätter skolen I göra och mina stadgar skolen I hålla, och skolen vandra efter dem.
Jag är HERREN, eder Gud.
Ja, I skolen hålla mina stadgar och rätter, ty den människa som gör efter dem skall leva genom dem.
Jag är HERREN.
Ingen bland eder skall komma vid någon kvinna som år hans nära blodsförvant och blotta hennes blygd.
Jag är HERREN.
Du skall icke blotta din faders blygd genom att blotta din moders blygd; hon är din moder, du skall icke blotta hennes blygd.
Du skall icke blotta någon annan kvinnas blygd, som är din faders hustru, ty det är din faders blygd.
Du skall icke blotta din systers blygd, evad hon är din faders dotter eller din moders dotter, evad hon är född hemma eller född ute.
Du skall icke blotta din sondotters eller din dotterdotters blygd, ty det är din egen blygd.
Du skall icke blotta din faders hustrus dotters blygd, ty hon är av din faders släkt, hon är din syster.
Du skall icke blotta din faders systers blygd; hon är din faders nära blodsförvant.
Du skall icke blotta din moders systers blygd, ty hon är din moders nära blodsförvant.
Du skall icke blotta din faders broders blygd: vid hans hustru skall du icke komma; hon är din faders syster.
Du skall icke blotta din svärdotters blygd; hon är din sons hustru, hennes blygd skall du icke blotta.
Du skall icke blotta din broders hustrus blygd, ty det är din broders blygd.
Du skall icke blotta en kvinnas blygd och tillika hennes dotters; du skall icke heller taga till hustru hennes sondotter eller dotterdotter och blotta dennas blygd, de äro ju nära blodsförvanter; sådant vore en skändlighet.
Och du skall icke till hustru taga en kvinna jämte hennes syster, så att du uppväcker fiendskap mellan dem, i det att du blottar den enas blygd och tillika den andras, medan den förra lever.
Du skall icke komma vid en kvinna och blotta hennes blygd, när hon är oren under sin månadsrening.
Med din nästas hustru skall du icke beblanda dig, så att du genom henne bliver oren.
Du skall icke giva någon av dina avkomlingar till offer åt Molok; du skall icke ohelga din Guds namn.
Jag är HERREN.
Du skall icke ligga hos en man såsom man ligger hos en kvinna; det är en styggelse.
Du skall icke beblanda där med något djur, så att du genom detta bliver oren.
Och ingen kvinna skall hava att skaffa med något djur, så att hon beblandar sig därmed; det är en vederstygglighet.
I skolen icke orena eder med något av allt detta, ty med allt sådant hava de hedningar orenat sig, som jag fördriver för eder.
Därigenom har landet blivit orenat, och jag har på det hemsökt dess missgärning, så att landet har utspytt sina inbyggare.
Så hållen då I mina stadgar och rätter, och ingen av eder, evad han är inföding eller en främling som bor ibland eder, må göra någon av alla dessa styggelser.
Ty alla dessa styggelser hava landets inbyggare, som hava varit där före eder, bedrivit, så att landet har blivit orenat.
Gören intet sådant, på det att landet icke må utspy eder, om I så orenen det, likasom det utspyr det folk som har bott där före eder.
Ty var och en som gör någon av alla dessa styggelser skall utrotas ur sitt folk, ja, var och en som gör sådant.
Iakttagen därför vad jag har bjudit eder iakttaga, så att I icke gören efter någon av de styggeliga stadgar som man har följt före eder, och så orenen eder genom dem.
Jag är HERREN, eder Gud.
Och HERREN talade till Mose och sade:
Tala till Israels barns hela menighet och säg till dem: I skolen vara heliga, ty jag, HERREN, eder Gud, är helig.
Var och en av eder frukte sin moder och sin fader.
Mina sabbater skolen I hålla.
Jag är HERREN, eder Gud.
I skolen icke vända eder till avgudar och icke göra eder gjutna gudar.
Jag är HERREN, eder Gud.
När I viljen offra tackoffer åt HERREN, skolen I offra det på sådant sätt att I bliven välbehagliga.
Samma dag I offren det skall det ätas, eller ock den följande dagen; men det som bliver över till tredje dagen skall brännas upp i eld.
Om det ätes på tredje dagen, så är det en vederstygglighet; det bliver då icke välbehagligt.
Den som äter därav kommer att bära på missgärning, ty han har ohelgat det som var helgat åt HERREN, och han skall utrotas ur sin släkt.
När I inbärgen skörden av edert land, skall du icke skörda intill yttersta kanten av din åker, icke heller skall du göra någon axplockning efter din skörd.
Och i din vingård skall du icke göra någon efterskörd, och de avfallna druvorna i din vingård skall du icke plocka upp; du skall lämna detta kvar åt den fattige och åt främlingen.
Jag är HERREN, eder Gud.
I skolen icke stjäla eller ljuga eller begå något svek mot varandra.
I skolen icke svärja falskt vid mitt namn; då ohelgar du din Guds namn.
Jag är HERREN.
Du skall icke med orätt avhända din nästa något, eller taga något ifrån honom med våld.
Du skall icke förhålla dagakarlen hans lön över natten till morgonen.
Du skall icke uttala förbannelser över en döv, och för en blind skall du icke lägga något varpå han kan falla; du skall frukta din Gud.
Jag är HERREN.
I skolen icke göra orätt i domen; du skall icke hava anseende till den ringes person, ej heller vara partisk för den mäktige; du skall döma din nästa rätt.
Du skall icke gå med förtal bland dina fränder; du skall icke stå efter din nästas blod.
Jag är HERREN.
Du skall icke hava hat till din broder i ditt hjärta, men väl må du tillrättavisa din nästa, så att du icke för hans skull kommer att bära på synd.
Du skall icke hämnas och icke hysa agg mot någon av ditt folk, utan du skall älska din nästa såsom dig själv.
Jag är HERREN.
Mina stadgar skolen I hålla: Du skall icke låta två slags djur av din boskap para sig med varandra; din åker skall du icke beså med två slags säd; en klädnad av två olika slags garn får icke komma på dig.
Om en man har legat hos en kvinna och beblandat sig med henne, och hon är trälinna i en annan mans våld, och hon icke har blivit friköpt eller frigiven, så skola de straffas, men icke dödas, eftersom hon icke var fri.
Och han skall föra fram sitt skuldoffer inför HERREN, till uppenbarelsetältets ingång, en skuldoffersvädur.
När så prästen medelst skuldoffersväduren bringar försoning för honom inför HERRENS ansikte för den synd han har begått, då bliver den synd han har begått honom förlåten.
När I kommen in i landet och planteren träd av olika slag med ätbar frukt, skolen I anse deras frukt såsom deras förhud.
I tre år skolen I hålla dem för oomskurna och icke äta av dem;
men under det fjärde året skall all deras frukt vara helgad till HERRENS lov,
och först under det femte skolen I äta deras frukt.
Så skolen I göra, för att de må giva så mycket större avkastning åt eder.
Jag är HERREN, eder Gud.
I skolen icke äta något med blod i.
I skolen icke befatta eder med spådom eller teckentyderi.
I skolen icke rundklippa kanten av edert huvudhår, ej heller skall du avstympa kanten av ditt skägg.
I skolen icke göra något märke på eder kropp för någon död, ej heller bränna in skrifttecken på eder.
Jag är HERREN.
Du skall icke ohelga din dotter med att låta henne bliva en sköka, på det att icke landet må förfalla i skökoväsende och bliva uppfyllt av skändlighet.
Mina sabbater skolen I hålla, och för min helgedom skolen I hava fruktan.
Jag är HERREN.
I skolen icke vända eder till andar som tala genom besvärjare eller spåmän.
Söken icke sådana, så att I bliven orena genom dem.
Jag är HERREN, eder Gud.
För ett grått huvud skall du stå upp, och den gamle skall du ära; du skall frukta din Gud.
Jag är HERREN.
När en främling bor hos eder i edert land, skolen I icke förtrycka honom.
Främlingen som bor hos eder skall räknas såsom en inföding bland eder, du skall älska honom såsom dig själv; I haven ju själva varit främlingar i Egyptens land.
Jag är HERREN, eder Gud.
I skolen icke göra orätt i domen, icke i fråga om mått, vikt eller mål.
Riktig våg, riktiga vikter, riktig efa, riktigt hin-mått skolen I hava.
Jag är HERREN, eder Gud, som har fört eder ut ur Egyptens land.
Så skolen I nu hålla alla mina stadgar och alla mina rätter och göra efter dem.
Jag är HERREN.
Och HERREN talade till Mose och sade:
Du skall ock säga till Israels barn: Om någon av Israels barn, eller av främlingarna som bo i Israel, giver någon av sina avkomlingar åt Molok, så skall han straffas med döden; folket i landet skall stena honom.
Och jag skall vända mitt ansikte mot den mannen och utrota honom ur hans folk, därför att han har givit en av sina avkomlingar åt Molok, och därmed orenat min helgedom och ohelgat mitt heliga namn.
Om folket i landet ser genom fingrarna med den mannen, när han giver en av sina avkomlingar åt Molok, så att de icke döda honom,
då skall jag själv vända mitt ansikte mot den mannen och mot hans släkt; och honom och alla dem som hava följt honom och i trolös avfällighet lupit efter Molok skall jag utrota ur deras folk.
Och om någon vänder sig till andar som tala genom besvärjare eller spåmän, för att i trolös avfällighet löpa efter dem, så skall jag vända mitt ansikte mot honom och utrota honom ur hans folk.
Så skolen I nu hålla eder heliga, och vara heliga; ty jag är HERREN, eder Gud.
Och I skolen hålla mina stadgar och göra efter dem.
Jag är HERREN, som helgar eder.
Om någon uttalar förbannelser över sin fader eller sin moder, skall han straffas med döden; över sin fader och sin moder har han uttalat förbannelser, blodskuld låder vid honom.
Om någon begår äktenskapsbrott med en annan mans hustru, om han begår äktenskapsbrott med sin nästas hustru, så skola de straffas med döden, både mannen och kvinnan som hava begått äktenskapsbrottet.
Om någon ligger hos en kvinna som är hans faders hustru, så blottar han sin faders blygd; de skola båda straffas med döden, blodskuld låder vid dem.
Om någon ligger hos sin svärdotter, så skola de båda straffas med döden; de hava bedrivit en vederstygglighet, blodskuld låder vid dem.
Om en man ligger hos en annan man såsom man ligger hos en kvinna, så göra de båda en styggelse; de skola straffas med döden, blodskuld låder vid dem.
Om någon till hustru tager en kvinna och tillika hennes moder, så är det en skändlighet; man skall bränna upp både honom och dem i eld, för att icke någon skändlighet må finnas bland eder.
Om en man beblandar sig med något djur, så skall han straffas med döden, och djuret skolen I dräpa.
Och om en kvinna kommer vid något djur och beblandar sig därmed, så skall du dräpa både kvinnan och djuret; de skola straffas med döden, blodskuld låder vid dem.
Om någon tager till hustru sin syster, sin faders dotter eller sin moders dotter, och ser hennes blygd och hon ser hans blygd, så är det en skamlig gärning, och de skola utrotas inför sitt folks ögon; han har blottat sin systers blygd, han bär på missgärning.
Om någon ligger hos en kvinna som har sin månadsrening och blottar hennes blygd, i det att han avtäcker hennes brunn och hon blottar sitt blods brunn, så skola de båda utrotas ur sitt folk.
Du skall icke blotta din moders systers eller din faders systers blygd.
Ty den så gör avtäcker sin nära blodsförvants blygd; de komma att bära på missgärning.
Om någon ligger hos sin farbroders hustru, så blottar han sin farbroders blygd; de komma att bära på synd, barnlösa skola de dö.
Om någon tager sin broders hustru, så är det en oren gärning; han blottar då sin broders blygd, barnlösa skola de bliva.
Så skolen I nu hålla alla mina stadgar och alla mina rätter och stadgar och göra efter dem, för att landet icke må utspy eder, det land dit jag vill föra eder, så att I fån bo där.
Och I skolen icke vandra efter det folks stadgar, som jag vill fördriva för eder; ty just därför att de hava bedrivit allt sådant, har jag blivit led vid dem.
Och därför har jag sagt till eder I skolen besitta deras land, ty jag skall giva eder det till besittning, ett land som flyter av mjölk och honung.
Jag är HERREN, eder Gud, som har avskilt eder från andra folk.
Gören alltså skillnad mellan rena fyrfotadjur och orena, och mellan rena fåglar och orena, så att I icke gören eder själva till styggelse för de fyrfotadjurs eller fåglars skull eller för de kräldjurs, skull på marken, som jag har avskilt, för att I skolen hålla dem för orena.
I skolen vara mig heliga, ty jag, HERREN, är helig, och jag har avskilt eder från andra folk, för att I skolen höra mig till.
När någon, man eller kvinna, befattar sig med andebesvärjelse eller spådom, skall denne straffas med döden; man skall stena honom, blodskuld låder vid honom.
Och HERREN sade till Mose: Säg till prästerna, Arons söner, säg till dem så: En präst får icke ådraga sig orenhet genom någon död bland sina fränder,
utom genom sina närmaste blodsförvanter: sin moder, sin fader, sin dotter, sin broder; son, sin dotter, sin broder;
så ock genom sin syster, om hon var jungfru och stod honom närmare och icke tillhörde någon man, i sådant fall må han ådraga sig orenhet genom henne.
Eftersom han är en herre bland sina fränder, får han icke ådraga sig orenhet och göra sig ohelig.
Prästerna skola icke raka någon del av sitt huvud skallig eller avraka kanten av sitt skägg eller rista något märke på sin kropp.
De skola vara helgade åt sin Guds och må icke ohelga sin Guds namn, ty de bära fram HERRENS eldsoffer sin Guds spis; därför skola de heliga.
Ingen av dem skall taga till hustru en sköka eller en vanärad kvinna, ej heller skall någon taga till hustru en kvinna som har blivit förskjuten av sin man, ty prästen är helgad åt sin Gud.
Därför skall du akta honom helig, ty han bär fram din Guds spis; han skall vara dig helig, ty jag, HERREN, som helgar eder, är helig.
Om en prästs dotter ohelgar sig genom skökolevnad, så ohelgar hon sin fader; hon skall brännas upp i eld.
Den som är överstepräst bland sina bröder, den på vilkens huvud smörjelseoljan har blivit utgjuten, och som har mottagit handfyllning till att ikläda sig prästkläderna, han skall icke hava sitt hår oordnat, ej heller riva sönder sina kläder;
och han skall icke gå in till någon död; icke ens genom sin fader eller genom sin moder får han ådraga sig orenhet.
Och ur helgedomen skall han icke gå ut, på det att han icke må ohelga sin Guds helgedom, ty hans Guds smörjelseolja, varmed han har blivit invigd, är på honom.
Jag är HERREN.
Till hustru skall han taga en kvinna som är jungfru.
En änka eller en förskjuten hustru eller en vanärad kvinna, en sköka -- en sådan får han icke taga, utan en jungfru bland sina fränder skall han taga till hustru,
för att han icke må ohelga sin livsfrukt bland sina fränder; ty jag är HERREN, som helgar honom.
Och HERREN talade till Mose och sade:
Tala till Aron och säg: Av dina avkomlingar i kommande släkten skall ingen som har något lyte träda fram för att frambära sin Guds spis.
Ingen skall träda fram, som har något lyte, varken en blind eller en halt, eller en som har lyte i ansiktet, eller som har någon lem för stor,
ingen som har brutit arm eller ben,
ingen som är puckelryggig eller förkrympt, eller som har fel på ögat, eller som har skabb eller annat utslag, eller som är snöpt.
Av prästen Arons avkomlingar skall ingen som har något lyte gå fram för att frambära HERRENS eldsoffer; han har ett lyte, han skall icke gå fram för att frambära sin Guds spis.
Sin Guds spis må han äta, både det som är högheligt och det som är heligt,
men eftersom han har ett lyte, skall han icke gå in till förlåten, ej heller skall han gå fram till altaret, på det att han icke må ohelga mina heliga ting; ty jag är HERREN, som helgar dem.
Och Mose talade detta till Aron och hans söner och alla Israels barn.
Och HERREN talade till Mose och sade:
Tala till Aron och hans söner och säg att de skola hålla sig ifrån de heliga gåvor som Israels barn bära fram åt mig, på det att de icke må ohelga mitt heliga namn.
Jag är HERREN.
Säg till dem: Om i kommande släkten någon av edra avkomlingar, medan orenhet låder vid honom, kommer vid de heliga gåvor som Israels barn bära fram åt HERREN, så skall han utrotas ur min åsyn Jag är HERREN.
Om någon av Arons avkomlingar är spetälsk eller har flytning, skall han icke äta av de heliga gåvorna, förrän han har blivit ren; ej heller den som kommer vid någon som har blivit oren genom en död, eller den som har haft sädesutgjutning;
ej heller den som kommer vid något slags smådjur genom vilket man bliver oren, eller vid en människa genom vilken man bliver oren, på vad sätt denna än må hava blivit oren.
Den som kommer vid något sådant, han skall vara oren ända till aftonen, och skall icke äta av de heliga gåvorna, förrän han har badat sin kropp i vatten.
Men när solen har gått ned, är han ren, och sedan må han äta av de heliga gåvorna, ty det är hans spis.
Ett självdött eller ihjälrivet djur skall han icke äta, så att han därigenom bliver oren.
Jag är HERREN.
De skola iakttaga vad jag har bjudit dem iakttaga, på det att de icke för det heligas skull må komma att bära på synd och träffas av döden därför att de ohelga det.
Jag är HERREN, som helgar dem.
Ingen främmande får äta av det heliga; en inhysesman hos prästen eller en hans legodräng skall icke äta av det heliga.
Men när en präst har köpt en träl för sina penningar, må denne äta därav, så ock den träl som är född i hans hus; dessa må äta av hans spis.
När en prästs dotter har blivit en främmande mans hustru, skall hon icke äta av det heliga som gives till offergärd.
Men om en prästs dotter har blivit änka eller blivit förskjuten, och hon är utan livsfrukt, och hon så kommer åter till sin faders hus och är där såsom i sin ungdom, då må hon äta av sin faders spis; men ingen främmande får äta därav.
Och om någon ouppsåtligen äter av det heliga, skall han lägga femtedelen därtill och giva prästen ersättning för det heliga.
Prästerna skola icke ohelga de heliga gåvorna, det som Israels barn göra såsom gärd åt HERREN,
och därigenom draga över dem missgärning och skuld, när de äta av deras heliga gåvor; ty jag är HERREN, som helgar dem.
Och HERREN talade till Mose och sade:
Tala till Aron och hans söner och alla Israels barn och säg till dem: Om någon av Israels hus eller av främlingarna i Israel vill offra något offer, vare sig det är ett löftesoffer eller ett frivilligt offer som de vilja offra åt HERREN såsom brännoffer, så skolen I göra det på sådant sätt att I bliven välbehagliga;
offret skall vara ett felfritt handjur, av fäkreaturen eller av fåren eller av getterna;
I skolen icke därtill taga ett djur som har något lyte, ty genom ett sådant bliven I icke välbehagliga.
Och när någon vill offra ett tackoffer åt HERREN av fäkreaturen eller av småboskapen, vare sig det gäller att fullgöra ett löfte, eller det gäller ett frivilligt offer, då skall det vara felfritt far att bliva välbehagligt; intet lyte får finnas därpå.
Det som är blint eller brutet eller stympat eller sårigt, eller det som har skabb eller annat utslag sådant skolen I icke offra åt HERREN; eldsoffer av sådant skolen I icke lägga på altaret åt HERREN.
Ett djur av fäkreaturen eller av småboskapen, som har någon lem för stor eller för liten, må du väl offra såsom frivilligt offer, men såsom löftesoffer bliver det icke välbehagligt.
Och I skolen icke offra åt HERREN något som har blivit snöpt genom klämning eller krossning eller avslitning eller utskärning; sådant skolen I icke göra i edert land.
Icke heller av en utlännings hand skolen I mottaga och offra sådana djur till eder Guds spis, ty de äro skadade, de hava ett lyte; genom sådana bliven I icke välbehagliga.
Och HERREN talade till Mose och sade:
När en kalv eller ett får eller en get har blivit född, skall djuret dia sin moder i sju dagar.
Men allt ifrån den åttonde dagen är det välbehagligt såsom eldsoffersgåva åt HERREN.
I skolen icke slakta något djur, vare sig av fäkreaturen eller av småboskapen, på samma dag som dess avföda.
När I viljen offra ett lovoffer åt HERREN, skolen I offra det på sådant sätt att I bliven välbehagliga.
Det skall ätas samma dag; I skolen icke lämna något därav kvar till följande morgon.
Jag är HERREN.
I skolen hålla mina bud och göra efter dem.
Jag är HERREN.
I skolen icke ohelga mitt heliga namn, ty jag vill bliva helgad bland Israels barn.
Jag är HERREN, som helgar eder,
han som har fört eder ut ur Egyptens land, för att jag skall vara eder Gud.
Jag är HERREN.
Och HERREN talade till Mose och sade:
Tala till Israels barn och säg till dem: Dessa äro HERRENS högtider, vilka I skolen utlysa såsom heliga sammankomster; mina högtider äro dessa:
Sex dagar skall arbete göras, men på sjunde dagen är vilosabbat, en dag för helig sammankomst; intet arbete skolen I då göra.
Det är HERRENS sabbat, var I än ären bosatta.
Dessa äro HERRENS högtider, de heliga sammankomster som I skolen utlysa på bestämda tider:
I första månaden, på fjortonde dagen i månaden, vid aftontiden, är HERRENS påsk.
Och på femtonde dagen i samma månad är HERRENS osyrade bröds högtid; då skolen I äta osyrat bröd, i sju dagar.
På den första dagen skolen I hålla en helig sammankomst; ingen arbetssyssla skolen I då göra.
Och I skolen offra eldsoffer åt HERREN i sju dagar.
På den sjunde dagen skall åter hållas en helig sammankomst; ingen arbetssyssla skolen I då göra.
Och HERREN talade till Mose och sade:
Tala till Israels barn och säg till dem: När I kommen in i det land som jag vill giva eder, och I inbärgen dess skörd, då skolen I bära till prästen den kärve som är förstlingen av eder skörd.
Och den kärven skall han vifta inför HERRENS ansikte, för att I mån bliva välbehagliga; dagen efter sabbaten skall prästen vifta den.
Och på den dag då I låten vifta kärven skolen I offra ett felfritt årsgammalt lamm till brännoffer åt HERREN,
och såsom spisoffer därtill två tiondedels efa fint mjöl, begjutet med olja, ett eldsoffer åt HERREN till en välbehaglig lukt, och såsom drickoffer därtill en fjärdedels hin vin.
Och intet av det nya, varken bröd eller rostade ax eller korn av grönskuren säd, skolen I äta förrän på denna samma dag, icke förrän I haven burit fram offergåvan åt eder Gud.
Detta skall vara en evärdlig stadga för eder från släkte till släkte, var I än ären bosatta.
Sedan skolen I räkna sju fulla veckor från dagen efter sabbaten, från den dag då I buren fram viftofferskärven;
femtio dagar skolen I räkna intill dagen efter den sjunde sabbaten; då skolen I bära fram ett offer av den nya grödan åt HERREN.
Från de orter där I bon skolen I bära fram viftoffersbröd, två kakor av två tiondedels efa fint mjöl, bakade med surdeg: en förstlingsgåva åt HERREN.
Och jämte brödet skolen I föra fram sju felfria årsgamla lamm, en ungtjur och två vädurar, till att offras såsom brännoffer åt HERREN, med tillhörande spisoffer och drickoffer: ett eldsoffer till en välbehaglig lukt för HERREN.
Därtill skolen I offra en bock till syndoffer och två årsgamla lamm till tackoffer.
Och prästen skall vifta dem såsom ett viftoffer inför HERRENS ansikte, jämte förstlingsbröden som bäras fram tillika med de båda lammen de skola vara helgade åt HERREN och tillhöra prästen.
Och till denna samma dag skolen I utlysa en helig sammankomst att hållas av eder; ingen arbetssyssla skolen I då göra.
Detta skall vara en evärdlig stadga för eder från släkte till släkte, var I än ären bosatta.
Och när I inbärgen skörden av edert land, skall du icke skörda intill yttersta kanten av din åker, icke heller skall du göra någon axplockning efter din skörd, du skall lämna detta kvar åt den fattige och åt främlingen.
Jag är HERREN, eder Gud.
Och HERREN talade till Mose och sade:
Tala till Israels barn och säg: I sjunde månaden, på första dagen i månaden, skolen I hålla sabbatsvila, en högtid med basunklang, till att bringa eder i åminnelse inför HERREN, en helig sammankomst.
Ingen arbetssyssla skolen I då göra, och I skolen offra eldsoffer åt HERREN.
Och HERREN talade till Mose och sade:
Men på tionde dagen i samma sjunde månad är försoningsdagen; då skolen I hålla en helig sammankomst, och I skolen då späka eder; och I skolen offra eldsoffer åt HERREN.
Och I skolen intet arbete göra på denna samma dag, ty det är en försoningsdag, då försoning bringas för eder inför HERRENS, eder Guds, ansikte.
Och var och en som icke späker sig på denna samma dag skall utrotas ur sin släkt.
Och var och en som gör något arbete på denna samma dag, honom skall jag förgöra ur hans folk.
Intet arbete skolen I då göra Detta skall vara en evärdlig stadga för eder från släkte till släkte, var I än ären bosatta.
En vilosabbat skall den vara för eder, och I skolen då späka eder.
På nionde dagen i månaden, om aftonen, skolen I hålla denna eder sabbatsvila, från afton till afton.
Och HERREN talade till Mose och sade:
Tala till Israels barn och säg: På femtonde dagen i samma sjunde månad är HERRENS lövhyddohögtid, i sju dagar.
På den första dagen skall man hålla en helig sammankomst; ingen arbetssyssla skolen I då göra.
I sju dagar skolen I offra eldsoffer åt HERREN.
På den åttonde dagen skolen I hålla en helig sammankomst och skolen offra eldsoffer åt HERREN.
Då är högtidsförsamling; ingen arbetssyssla skolen I då göra.
Dessa äro HERRENS högtider, vilka I skolen utlysa såsom heliga sammankomster, och på vilka I skolen offra eldsoffer åt HERREN, brännoffer och spisoffer, slaktoffer och drickoffer, var dag de för den dagen bestämda offren --
detta förutom HERRENS sabbater, och förutom edra övriga gåvor, och förutom alla edra löftesoffer, och förutom alla frivilliga offer som I given åt HERREN.
Men på femtonde dagen i sjunde månaden, när I inbärgen avkastningen av landet, skolen I fira HERRENS högtid, i sju dagar.
På den första dagen är sabbatsvila, på den åttonde dagen är ock sabbatsvila.
Och I skolen på den första dagen taga frukt av edra skönaste träd, kvistar av palmer och grenar av lummiga träd och av pilträd, och skolen så vara glada i sju dagar inför HERRENS, eder Guds, ansikte.
I skolen fira denna högtid såsom en HERRENS högtid sju dagar om året.
Detta skall vara en evärdlig stadga för eder från släkte till släkte; i sjunde månaden skolen I fira den.
Då skolen I bo i lövhyddor i sju dagar; alla de som äro infödingar i Israel skola bo i lövhyddor,
för att edra efterkommande må veta huru jag lät Israels barn bo i lövhyddor, när jag förde dem ut ur Egyptens land Jag är HERREN, eder Gud.
Och Mose talade till Israels barn om dessa HERRENS högtider.
Och HERREN talade till Mose och sade:
Bjud Israels barn att bära till dig ren olja, av stötta oliver, till ljusstaken, så att lamporna dagligen kunna sättas upp.
Utanför den förlåt som hänger framför vittnesbördet, i uppenbarelsetältet, skall Aron beständigt sköta den, från aftonen till morgonen, inför HERRENS ansikte.
Detta skall vara en evärdlig stadga för eder från släkte till släkte.
Lamporna på den gyllene ljusstaken skall han beständigt sköta inför HERRENS ansikte.
Och du skall taga fint mjöl och därav baka tolv kakor; var kaka skall innehålla två tiondedels efa.
Och du skall lägga upp dem i två rader, sex i var rad, på det gyllene bordet inför HERRENS ansikte.
Och på vardera raden skall du lägga ren rökelse, för att denna må utgöra själva altaroffret av bröden, ett eldsoffer åt HERREN.
Sabbatsdag efter sabbatsdag skall man beständigt lägga upp dem inför HERRENS ansikte: en gärd av Israels barn, till ett evigt förbund.
De skola tillhöra Aron och hans söner och skola ätas av dem på en helig plats, ty de äro högheliga och äro hans evärdliga rätt av HERRENS eldsoffer.
Och en man som var son till en israelitisk kvinna, men till fader hade en egyptisk man, gick ut bland Israels barn; och den israelitiska kvinnans son och en israelitisk man kommo i träta med varandra i lägret.
Och den israelitiska kvinnans son smädade Namnet och hädade.
Då förde de honom fram till Mose.
Och hans moder hette Selomit, dotter till Dibri, av Dans stam.
Och de satte honom i förvar, för att de skulle få hans dom bestämd efter HERRENS befallning.
Och HERREN talade till Mose och sade:
För ut hädaren utanför lägret; sedan må alla som hörde det lägga sina händer på hans huvud, och må så hela menigheten stena honom.
Och till Israels barn skall du tala och säga: Om någon hädar sin Gud, kommer han att bära på synd.
Och den som smädar HERRENS namn skall straffas med döden; hela menigheten skall stena honom.
Evad det är en främling eller en inföding som smädar Namnet, skall han dödas.
Om någon slår ihjäl någon människa, skall han straffas med döden;
och den som slår ihjäl ett boskapsdjur skall ersätta det: liv för liv.
Och om någon vållar att hans nästa får ett lyte, så skall man göra mot honom såsom han själv har gjort:
bruten lem för bruten lem, öga för öga, tand för tand; samma lyte han har vållat att en annan fick skall han själv få.
Den som slår ihjäl ett boskapsdjur skall ersätta det, och den som slår ihjäl en människa skall dödas.
En och samma lag skall gälla för eder, den skall gälla lika väl för främlingen som för infödingen; ty jag är HERREN, eder Gud.
Och Mose talade detta till Israels barn; och de förde ut hädaren utanför lägret och stenade honom.
Alltså gjorde Israels barn såsom HERREN hade bjudit Mose.
Och HERREN talade till Mose på Sinai berg och sade:
Tala till Israels barn och säg till dem: När I kommen in i det land som jag vill giva eder, skall landet hålla sabbat åt HERREN.
I sex år skall du beså din åker, och i sex år skära din vingård och inbärga avkastningen av landet,
men under det sjunde året skall landet hava vilosabbat, en HERRENS sabbat; då skall du icke beså din åker och icke skära din vingård.
Vad som växer upp av spillsäden efter din skörd skall du icke skörda, och de druvor som växa på dina oskurna vinträd skall du icke avbärga.
Det skall vara ett sabbatsvilans år för landet.
Och vad landets sabbat ändå giver skolen I hava till föda: du själv, din tjänare och din tjänarinna, din daglönare och din inhysesman, de som bo hos dig.
Din boskap och de vilda djuren i ditt land skola ock hava sin föda av all dess avkastning.
Och du skall räkna sju årsveckor, det är sju gånger sju år, så att tiden för de sju årsveckorna bliver fyrtionio år.
Då skall du i sjunde månaden, på tionde dagen i månaden, låta blåsa i larmbasun; på försoningsdagen skolen I blåsa i basun över hela edert land.
Och I skolen helga det femtionde året och utropa frihet i landet för alla dess inbyggare.
Det skall vara ett jubelår för eder; var och en av eder skall då återfå sin arvsbesittning, var och en av eder skall återfå sin släktegendom.
Ett jubelår skall detta femtionde år vara för eder; då skolen I icke så något, och vad som då växer upp av spillsäden skolen I icke skörda, och I skolen då icke avbärga edra oskurna vinträd.
Ty det är ett jubelår; heligt skall det vara för eder.
Från själva marken skolen I hämta eder föda, av dess avkastning.
Under ett sådant jubelår skall var och en av eder återfå sin arvsbesittning.
Om I alltså säljer något åt eder nästa eller köpen något av eder nästa, skolen I icke göra varandra orätt:
efter antalet år från jubelåret skall du betala din nästa, efter antalet årsgrödor skall han få betalning av dig.
Alltefter som åren äro flera skall du betala högre pris, och alltefter som åren äro färre skall du betala lägre pris; ty ett visst antal grödor är det han säljer till dig.
I skolen icke göra varandra orätt du skall frukta din Gud; ty jag är HERREN, eder Gud.
Och I skolen göra efter mina stadgar, och mina rätter skolen I hålla och skolen göra efter dem; då skolen I bo trygga i landet.
Och landet skall giva sin frukt, så att I haven nog att äta, och I skolen bo trygga däri.
Och om I frågen: »Vad skola vi äta under det sjunde året, om vi icke få så och icke få inbärga vår gröda?»,
så mån I veta att jag skall bjuda min välsignelse komma över eder under det sjätte året, så att det giver gröda för de tre åren.
Och ännu när I under det åttonde året sån, skolen I hava av den gamla grödan att äta; ända till dess att grödan på det nionde året har kommit in, skolen I hava gammalt att äta.
När I säljen jord, skolen I icke sälja den för evärdlig tid, ty landet är mitt; I ären ju främlingar och gäster hos mig.
I hela det land I fån till besittning skolen I medgiva rätt att återbörda jordegendom.
Om din broder råkar i armod och säljer något av sin arvsbesittning, så må hans närmaste bördeman komma till honom och återbörda det brodern har sålt.
Och om någon icke har någon bördeman, men han själv kommer i tillfälle att anskaffa vad som behöves för att återbörda,
så skall han räkna efter, huru många år som hava förflutit ifrån försäljningen, och betala lösen för de återstående åren åt den man till vilken han sålde, och han skall så återfå sin besittning.
Men om han icke förmår anskaffa vad som behöves till att betala honom, så skall det han har sålt förbliva i köparens hand intill jubelåret.
Men på jubelåret skall det frånträdas, och han skall då återfå sin besittning.
Om någon säljer ett boningshus i en stad som är omgiven med murar, så skall han hava rätt att återbörda det innan ett år har förflutit, sedan han sålde det; hans rätt att återbörda det är då inskränkt till viss tid.
Men om det icke har blivit återbördat, förrän hela året är ute, så skall huset, om det ligger i en stad som är omgiven med murar, förbliva köparens och hans efterkommandes egendom för evärdlig tid; det skall då icke frånträdas på jubelåret.
Men hus i sådana byar som icke hava murar omkring sig skola räknas till landets åkermark; de skola kunna återbördas, och på jubelåret skola de frånträdas.
Dock skola leviterna inom de städer som äro deras arvsbesittning hava evärdlig rätt att återbörda husen i städerna
Också om någon annan av leviterna inlöser det sålda huset i den stad där han har sin besittning, skall det dock frånträdas på jubelåret; ty husen i levitstäderna äro leviternas arvsbesittning bland Israels barn.
Och ett fält som är utmark omkring någon av deras städer får icke säljas, ty det är deras evärdliga besittning.
Om din broder råkar i armod och kommer på obestånd hos dig, så skall du taga dig an honom; såsom en främling eller en inhysesman skall han få leva hos dig.
Du skall icke ockra på honom eller taga ränta, ty du skall frukta din Gud, och du skall låta din broder leva hos dig.
Du skall icke lämna honom dina penningar på ocker eller lämna honom av dina livsmedel mot ränta.
Jag är HERREN, eder Gud, som har fört eder ut ur Egyptens land, för att giva eder Kanaans land och vara eder Gud.
Om din broder råkar i armod hos dig och säljer sig åt dig, skall du icke låta honom göra trälarbete;
såsom en daglönare och en inhysesman skall han vara hos dig; intill jubelåret skall han tjäna hos dig.
Då skall du giva honom fri, honom själv och hans barn med honom; och han skall återfå sin släktegendom, sin fädernebesittning skall han återfå.
Ty de äro mina tjänare, som jag har fört ut ur Egyptens land; de skola icke säljas såsom man säljer trälar.
Du skall icke med hårdhet bruka din makt över dem; du skall frukta din Gud.
Men om du vill skaffa dig en verklig träl eller trälinna, så skall du köpa en sådan träl eller trälinna från hedningarna som bo runt omkring eder.
I mån ock köpa sådana ibland barnen till inhysesmännen som bo hos eder och bland personer av deras släkt, som I haven hos eder, och som äro födda i edert land; sådana skola förbliva eder egendom.
Och dem mån I hava att lämna såsom arv åt edra barn efter eder, till egendom och besittning; dem kunnen I hava till trälar evärdligen.
Men ibland edra bröder, Israels barn, skall ingen med hårdhet bruka sin makt över den andre.
Om en främling eller en inhysesman hos dig kommer till välstånd, och en din broder råkar i armod hos honom och säljer sig åt främlingen som bor inhyses hos dig, eller eljest åt någon som tillhör en främlingssläkt,
så skall han sedan, efter det att han har sålt sig, kunna lösas ut; någon av hans bröder må lösa honom;
eller ock må hans farbroder eller hans farbroders son lösa honom, eller må någon annan nära blodsförvant av hans släkt lösa honom; eller om han kommer i tillfälle därtill, må han själv lösa sig.
Därvid skall han, jämte den som har köpt honom, räkna efter, huru lång tid som har förflutit ifrån det år då han sålde sig åt honom till jubelåret; och det pris för vilket han såldes skall uppskattas efter årens antal; hans arbetstid hos honom skall beräknas till samma värde som en daglönares.
Om ännu många år äro kvar, skall han såsom lösen för sig betala en motsvarande del av det penningbelopp som han köptes för.
Om däremot allenast få år återstå till jubelåret, så skall han räkna efter detta, sig till godo, och betala lösen för sig efter antalet av sina år.
Såsom en daglönare som är lejd för år skall man behandla honom ingen må inför dina ögon med hårdhet bruka sin makt över honom.
Men om han icke bliver löst på något av de nämnda sätten, så skall han på jubelåret givas fri, han själv och hans barn med honom.
Ty Israels barn äro mina tjänare; de äro mina tjänare, som jag har fört ut ur Egyptens land.
Jag är HERREN, eder Gud.
I skolen icke göra eder några av gudar, ej heller uppresa åt eder något beläte eller någon stod, eller uppsätta i edert land stenar med inhuggna bilder, för att tillbedja vid dem; ty jag är HERREN, eder Gud.
Mina sabbater skolen I hålla, och för min helgedom skolen I hava fruktan.
Jag är HERREN.
Om I vandren efter mina stadgar och hållen mina bud och gören efter dem,
så skall jag giva eder regn i rätt tid, så att jorden giver sin gröda och träden på marken bära sin frukt.
Och trösktiden skall hos eder räcka intill vinbärgningen, och vinbärgningen skall räcka intill såningstiden, och I skolen hava bröd nog att äta och skolen bo trygga i edert land.
Och jag skall skaffa frid i landet, och I skolen få ro, och ingen skall förskräcka eder.
Jag skall göra slut på vilddjuren i landet, och intet svärd skall gå fram genom edert land.
I skolen jaga edra fiender framför eder, och de skola falla för edra svärd.
Fem av eder skola jaga hundra framför sig, och hundra av eder skola jaga tiotusen, och edra fiender skola falla för edra svärd.
Och jag skall vända mig till eder och göra eder fruktsamma och för öka eder, och jag skall upprätthålla mitt förbund med eder.
Och gammal gröda, som länge har legat inne, skolen I hava att äta; I skolen nödgas skaffa den gamla undan för den nya.
Och jag skall uppresa min boning mitt ibland eder, och min själ skall icke försmå eder.
Jag skall vandra mitt ibland eder och vara eder Gud, och I skolen vara mitt folk.
Jag är HERREN, eder Gud, som förde eder ut ur Egyptens land, för att I icke skullen vara trälar där; och jag har brutit sönder edert ok och låtit eder gå med upprätt huvud.
Men om I icke hören mig och icke gören efter alla dessa bud,
om I förkasten mina stadgar, och om edra själar försmå mina rätter, så att I icke gören efter alla mina bud, utan bryten mitt förbund,
då skall ock jag handla på samma sätt mot eder: jag skall hemsöka eder med förskräckliga olyckor, med tärande sjukdom och feber, så att edra ögon försmäkta och eder själ förtvinar; och I skolen förgäves så eder säd, ty edra fiender skola äta den.
Jag skall vända mitt ansikte mot eder, och I skolen bliva slagna av edra fiender; och de som hata eder skola råda över eder, och I skolen fly, om ock ingen förföljer eder.
Om I, detta oaktat, icke hören mig, så skall jag tukta eder sjufalt värre för edra synders skull.
Jag skall krossa eder stolta makt.
Jag skall låta eder himmel bliva såsom järn och eder jord såsom koppar.
Och eder möda skall vara förspilld, ty eder jord skall icke giva sin gröda, och träden i landet skola icke bära sin frukt.
Om I ändå vandren mig emot och icke viljen höra mig, så skall jag slå eder sjufalt värre, såsom edra synder förtjäna.
Jag skall sända över eder vilddjur, som skola döda edra barn och fördärva eder boskap och minska edert eget antal, så att edra vägar bliva öde.
Om I, detta oaktat, icke låten varna eder av mig, utan vandren mig emot,
så skall också jag vandra eder emot och slå eder sjufalt för edra synders skull.
Jag skall låta eder drabbas av ett hämndesvärd, som skall hämnas mitt förbund, och I skolen nödgas församla eder i städerna; men där skall jag sända pest bland eder, och I skolen bliva givna i fiendehand.
Jag skall så fördärva edert livsuppehälle, att edert bröd skall kunna bakas i en enda ugn av tio kvinnor, och edert bröd skall lämnas ut efter vikt, och när I äten, skolen I icke bliva mätta.
Om I, detta oaktat, icke hören mig, utan vandren mig emot,
så skall också jag i vrede vandra eder emot och tukta eder sjufalt för edra synders skull.
I skolen nödgas äta edra söners kött och äta edra döttrars kött.
Jag skall ödelägga edra offerhöjder och utrota edra solstoder; jag skall kasta edra döda kroppar på edra eländiga avgudars döda kroppar, ty min själ skall försmå eder.
Och jag skall göra edra städer till ruiner och föröda edra helgedomar, och jag skall icke mer med välbehag känna lukten av edra offer.
Jag skall själv ödelägga landet, så att edra fiender, som bo däri, skola häpna däröver.
Men eder skall jag förströ bland hedningarna, och jag skall förfölja eder med draget svärd; så skall edert land bliva en ödemark, och edra städer skola bliva ruiner.
Då skall landet få gottgörelse för sina sabbater, då, under hela den tid det ligger öde och I ären i edra fienders land.
Ja, då skall landet hålla sabbat och giva gottgörelse för sina sabbater.
Hela den tid det ligger öde skall det hålla sabbat och få den vila det icke fick på edra sabbater, då I bodden däri.
Och åt dem som bliva kvar av eder skall jag giva försagda hjärtan i deras fienders länder, så att de jagas på flykten av ett prasslande löv som röres av vinden, och fly, såsom flydde de för svärd, och falla, om ock ingen förföljer dem.
Och de skola stupa på varandra, likasom för svärd, om ock ingen förföljer dem.
Ja, I skolen icke kunna hålla stånd mot edra fiender.
I skolen förgås bland hedningarna, och edra fienders land skall förtära eder.
Och de som bliva kvar av eder skola försmäkta i edra fienders land, genom sin egen missgärning, och försmäkta tillika genom sina fäders missgärning, likasom dessa hava gjort.
Och de skola nödgas bekänna den missgärning de själva hava begått, och den deras fäder hava begått, genom att handla trolöst mot mig, och huru de hava vandrat mig emot
-- varför också jag måste vandra dem emot och föra dem bort i deras fienders land -- ja, då skola deras oomskurna hjärtan nödgas ödmjuka sig, då skola de få umgälla sin missgärning.
Och då skall jag tänka på mitt förbund med Jakob, då skall jag ock tänka på mitt förbund med Isak och på mitt förbund med Abraham, och på landet skall jag tänka.
Ty landet måste bliva övergivet av dem och så få gottgörelse för sina sabbater genom att bliva öde när folket är borta, och själva skola de få umgälla sin missgärning, därför, ja, därför att de förkastade mina rätter, och därför att deras själar försmådde mina stadgar.
Men detta oaktat skall jag, medan de äro i sina fienders land, icke så förkasta eller försmå dem, att jag förgör dem och bryter mitt förbund med dem; ty jag är HERREN, deras Gud.
Nej, till fromma för dem skall jag tänka på förbundet med förfäderna, som jag förde ut ur Egyptens land, inför hedningarnas ögon, på det att jag skulle vara deras Gud.
Jag är HERREN.
Dessa äro de stadgar och rätter och lagar som HERREN fastställde mellan sig och Israels barn, på Sinai berg genom Mose.
Och HERREN talade till Mose och sade:
Tala till Israels barn och säg till dem: Om någon skall fullgöra ett löfte, ett sådant varvid du har att bestämma värdet på personer som lovas åt HERREN, så gäller följande:
Om värdet skall bestämmas för en man som är mellan tjugu och sextio år gammal, så skall du bestämma detta till femtio siklar silver, efter helgedomssikelns vikt.
Om frågan gäller en kvinna, så skall du bestämma värdet till trettio siklar.
Om frågan gäller någon som är mellan fem år och tjugu år gammal, så skall det värde du bestämmer vara för mankön tjugu siklar och för kvinnkön tio siklar.
Om frågan gäller någon som är mellan en månad och fem år gammal, så skall det värde du bestämmer vara för mankön fem siklar silver och för kvinnkön tre siklar silver.
Om frågan gäller någon som är sextio år gammal eller därutöver, så skall det värde du bestämmer vara, om det är en man, femton siklar, men för en kvinna skall det vara tio siklar.
Är någon i sådant armod att han icke kan betala det värde du bestämmer, så skall han ställas fram inför prästen, och prästen skall då bestämma ett värde för honom; efter vad den som har gjort löftet kan anskaffa skall prästen bestämma värdet för honom.
Om frågan gäller boskap, av de lag man får bära fram såsom offer åt HERREN, så skall allt sådant, när man har givit det åt HERREN, vara heligt;
man skall icke utväxla eller utbyta det, vare sig ett bättre mot ett sämre eller ett sämre mot ett bättre.
Om någon likväl utbyter ett djur mot ett annat, så skall både det förra och det som har blivit lämnat i utbyte vara heligt.
Men om frågan gäller något slags orent djur, ett sådant som man icke får bära fram såsom offer åt HERREN, så skall djuret ställas fram inför prästen;
och prästen skall bestämma dess värde, alltefter som det är bättre eller sämre.
Såsom du -- prästen -- bestämmer det, så skall det vara.
Och om ägaren vill lösa djuret, så skall han till det värde du har bestämt lägga femtedelen av värdet.
Om någon helgar sitt hus, för att det skall vara helgat åt HERREN, så skall prästen bestämma dess värde, alltefter som det är bättre eller sämre.
Såsom prästen bestämmer dess värde, så skall det förbliva.
Och om den som har helgat sitt hus vill lösa det, så skall han till det värde i penningar du har bestämt lägga femtedelen därav; då bliver det hans.
Om någon helgar åt HERREN ett stycke åker av sin arvsbesittning så skall du bestämma dess värde efter utsädet därpå: mot var homer utsädeskorn skola svara femtio siklar silver.
Om han helgar sin åker ända från jubelåret, så skall det förbliva vid det värde du bestämmer.
Men om han helgar sin åker efter jubelåret, då skall prästen åt honom beräkna penningvärdet efter antalet av de år som återstå till nästa jubelår; och ett motsvarande avdrag skall göras på det värde du förut har bestämt.
Och om den som har helgat åkern vill lösa den, så skall han till det värde i penningar du har bestämt lägga femtedelen därav; då förbliver den hans.
Om han icke löser åkern, men säljer den åt någon annan, så får åkern sedan icke lösas,
utan när åkern frånträdes på jubelåret, skall den vara helgad åt HERREN, likasom en tillspillogiven åker; hans arvsbesittning tillfaller då prästen.
Om någon helgar åt HERREN en åker som han har köpt, en som icke hör till hans arvsbesittning,
så skall prästen åt honom räkna ut beloppet av det bestämda värdet intill jubelåret; och han skall samma dag erlägga detta värde, som du har bestämt; det skall vara helgat åt HERREN.
Men på jubelåret skall åkern återgå till den av vilken den har blivit köpt, och vilkens arvejord den är.
Och när du bestämmer något värde, skall det alltid bestämmas i helgedomssiklar, sikeln räknad till tjugu gera.
Men det som är förstfött ibland boskap, och som tillhör HERREN redan såsom förstfött, det skall ingen helga; vare sig det är ett djur av fäkreaturen eller ett djur av småboskapen, tillhör det redan HERREN
Men om frågan gäller något orent djur, så skall man lösa det efter det värde du bestämmer och lägga femtedelen av värdet därtill.
Om det icke löses, så skall det säljas efter det värde du bestämmer.
Och om frågan gäller något tillspillogivet, vad någon har givit till spillo åt HERREN av sin egendom, det må vara en människa eller ett boskapsdjur eller den åker som är hans arvsbesittning, så får sådant varken säljas eller lösas; allt tillspillogivet är högheligt och tillhör HERREN.
En människa som har blivit tillspillogiven får aldrig lösas; en sådan måste dödas.
Och all tionde av jorden, vare sig av säden på jorden eller av trädens frukt, tillhör HERREN; den är helgad åt HERREN.
Om någon vill lösa något av sin tionde, så skall han lägga femtedelen av värdet därtill.
Och vad beträffar tionde av fäkreatur eller av småboskap, allt som går under herdestaven, så skall av allt detta vart tionde djur vara helgat åt HERREN;
man skall icke efterforska om det är bättre eller sämre, och man får icke utbyta det.
Om någon likväl utbyter djuret, så skall både detta och det som har blivit lämnat i utbyte vara heligt; det får icke lösas.
Dessa äro de bud som HERREN på Sinai berg gav Israels barn genom Mose.
Och HERREN talade till Mose i Sinais öken, i uppenbarelsetältet, på första dagen i andra månaden av det andra året efter deras uttåg ur Egyptens land; han sade:
»Räknen antalet av Israels barn, deras hela menighet, efter deras släkter och efter deras familjer, vart namn räknat särskilt, allt mankön, var person för sig;
alla stridbara män i Israel, de män som äro tjugu år gamla eller därutöver, dem skolen I inmönstra efter deras häravdelningar, du och Aron.
I skolen därvid taga till eder en man av var stam, den som är huvudman för sin stams familjer.
Och dessa äro namnen på de män som skola biträda eder: av Ruben: Elisur, Sedeurs son;
av Simeon: Selumiel, Surisaddais son;
av Juda: Naheson, Amminadabs son;
av Isaskar: Netanel, Suars son;
av Sebulon: Eliab, Helons son;
av Josefs barn: av Efraim: Elisama, Ammihuds son; av Manasse: Gamliel, Pedasurs son;
av Benjamin: Abidan, Gideonis son;
av Dan: Ahieser, Ammisaddais son;
av Aser: Pagiel, Okrans son;
av Gad: Eljasaf, Deguels son;
av Naftali: Ahira, Enans son.»
Dessa voro ombud för menigheten, hövdingar för sina fädernestammar, huvudmän för Israels ätter.
Och Mose och Aron togo till sig dessa namngivna män;
och sedan de hade församlat hela menigheten på första dagen i andra månaden, blev folket infört i förteckningen efter sina släkter och efter sina familjer, vart namn räknat särskilt, de som voro tjugu år gamla eller därutöver, var person för sig,
allt såsom HERREN hade bjudit Mose; och han mönstrade dem i Sinais öken.
Och avkomlingarna av Rubens, Israels förstföddes, söner, upptecknade efter sina släkter och efter sina familjer, vart namn räknat särskilt, var person för sig, alla av mankön som voro tjugu år gamla eller därutöver, alla stridbara män,
så många av Rubens stam som inmönstrades, utgjorde fyrtiosex tusen fem hundra.
Avkomlingarna av Simeons söner, upptecknade efter sina släkter och efter sina familjer, så många som inmönstrades, vart namn räknat särskilt, var person för sig, alla av mankön som voro tjugu år gamla eller därutöver, alla stridbara män,
så många av Simeons stam som inmönstrades, utgjorde femtionio tusen tre hundra.
Avkomlingarna av Gads söner, upptecknade efter sina släkter och efter sina familjer, vart namn räknat särskilt, de som voro tjugu år gamla eller därutöver, alla stridbara män,
så många av Gads stam som inmönstrades, utgjorde fyrtiofem tusen sex hundra femtio.
Avkomlingarna av Judas söner, upptecknade efter sina släkter och efter sina familjer, vart namn räknat särskilt, de som voro tjugu år gamla eller därutöver, alla stridbara män,
så många av Juda stam som inmönstrades, utgjorde sjuttiofyra tusen sex hundra.
Avkomlingarna av Isaskars söner, upptecknade efter sina släkter och efter sina familjer, vart namn räknat särskilt, de som voro tjugu år gamla eller därutöver, alla stridbara män,
så många av Isaskars stam son inmönstrades, utgjorde femtiofyra tusen fyra hundra.
Avkomlingarna av Sebulons söner upptecknade efter sina släkter och efter sina familjer, vart namn räknat särskilt, de som voro tjugu år gamla eller därutöver, alla stridbara män,
så många av Sebulons stam som inmönstrades, utgjorde femtiosju tusen fyra hundra.
Avkomlingarna av Josefs söner: Avkomlingarna av Efraims söner, upptecknade efter sina släkter och efter sina familjer, vart namn räknat särskilt, de som voro tjugu år gamla eller därutöver, alla stridbara män,
så många av Efraims stam som inmönstrades; utgjorde fyrtio tusen fem hundra.
Avkomlingarna av Manasses söner, upptecknade efter sina släkter och efter sina familjer, vart namn räknat särskilt, de som voro tjugu år gamla eller därutöver, alla stridbara män,
så många av Manasse stam som inmönstrades, utgjorde trettiotvå tusen två hundra.
Avkomlingarna av Benjamins söner, upptecknade efter sina släkter och efter sina familjer, vart namn räknat särskilt, de som voro tjugu år gamla eller därutöver, alla stridbara män,
så många av Benjamins stam som inmönstrades, utgjorde trettiofem tusen fyra hundra.
Avkomlingarna av Dans söner, upptecknade efter sina släkter och efter sina familjer, vart namn räknat särskilt, de som voro tjugu år gamla eller därutöver, alla stridbara män,
så många av Dans stam som inmönstrades, utgjorde sextiotvå tusen sju hundra.
Avkomlingarna av Asers söner, upptecknade efter sina släkter och efter sina familjer, vart namn räknat särskilt, de som voro tjugu år gamla eller därutöver, alla stridbara män,
så många av Asers stam som inmönstrades, utgjorde fyrtioett tusen fem hundra.
Avkomlingarna av Naftalis söner, upptecknade efter sina släkter och efter sina familjer, vart namn räknat särskilt, de som voro tjugu år gamla eller därutöver, alla stridbara män,
så många av Naftali stam som inmönstrades, utgjorde femtiotre tusen fyra hundra.
Dessa voro de inmönstrade, de som blevo inmönstrade av Mose och Aron och Israels hövdingar, tolv män, som företrädde var och en sin stamfamilj.
Och alla de av Israels barn som inmönstrades, efter deras familjer, de som voro tjugu år gamla eller därutöver, alla stridbara män i Israel,
alla dessa inmönstrade utgjorde sex hundra tre tusen fem hundra femtio.
Men leviterna i sin fädernestam blevo icke inmönstrade med de övriga.
Ty HERREN talade till Mose och sade:
Levi stam allenast skall du icke inmönstra, och du skall icke räkna antalet av dem med de övriga israeliterna;
utan du skall förordna leviterna att förestå vittnesbördets tabernakel med alla dess redskap och alla dess tillbehör.
De skola bära tabernaklet och alla dess redskap och göra tjänst därvid; och runt omkring tabernaklet skola de hava sitt läger.
När tabernaklet skall bryta upp, skola leviterna nedtaga det, och när tabernaklet skall slås upp, skola leviterna uppsätta det; men om någon främmande kommer därvid, skall han dödas.
De övriga israeliterna skola lägra sig var och en i sitt läger, och var och en under sitt baner, efter sina häravdelningar;
men leviterna skola lägra sig runt omkring vittnesbördets tabernakel, för att icke förtörnelse må komma över Israels barns menighet; och leviterna skola iakttaga vad som är att iakttaga vid vittnesbördets tabernakel.
Och Israels barn gjorde så; de gjorde i alla stycken såsom HERREN hade bjudit Mose.
Och HERREN talade till Mose och Aron och sade:
Israels barn skola lägra sig var och en under sitt baner, vid de fälttecken som höra till deras särskilda familjer; runt omkring uppenbarelsetältet skola de lägra sig så, att de hava det framför sig.
På framsidan, österut, skall Juda lägra sig under sitt baner, efter sina häravdelningar: Juda barns hövding Naheson, Amminadabs son
med de inmönstrade som utgöra hans här, sjuttiofyra tusen sex hundra man.
Bredvid honom skall Isaskars stam lägra sig: Isaskars barns hövding Netanel, Suars son,
med de inmönstrade som utgöra hans här, femtiofyra tusen fyra hundra man.
Därnäst Sebulons stam: Sebulons barns hövding Eliab, Helons son,
med de inmönstrade som utgöra hans här, femtiosju tusen fyra hundra man.
De inmönstrade som tillhöra Juda läger utgöra alltså tillsammans ett hundra åttiosex tusen fyra hundra man, delade i sina häravdelningar.
De skola vid uppbrott tåga främst.
Ruben skall lägra sig under sitt baner söderut, efter sina häravdelningar: Rubens barns hövding Elisur, Sedeurs son,
med de inmönstrade som utgöra hans här, fyrtiosex tusen fem hundra man.
Bredvid honom skall Simeons stam lägra sig: Simeons barns hövding Selumiel, Surisaddais son,
med de inmönstrade som utgöra hans här, femtionio tusen tre hundra man.
Därnäst Gads stam: Gads barns hövding Eljasaf, Reguels son
med de inmönstrade som utgöra hans här, fyrtiofem tusen sex hundra femtio man.
De inmönstrade som tillhöra Rubens läger utgöra alltså tillsammans ett hundra femtioett tusen fyra hundra femtio man, delade i sina häravdelningar.
Och de skola vid uppbrott tåga i andra rummet.
Sedan skall uppenbarelsetältet med leviternas läger hava sin plats i tåget, mitt emellan de övriga lägren.
I den ordning de lägra sig skola de ock tåga, var och en på sin plats, under sina baner.
Efraim skall lägra sig under sitt baner västerut, efter sina häravdelningar: Efraims barns hövding Elisama, Ammihuds son,
med de inmönstrade som utgöra hans här, fyrtio tusen fem hundra man.
Bredvid honom skall Manasse stam lägra sig: Manasse barns hövding Gamliel, Pedasurs son,
med de inmönstrade som utgöra hans här, trettiotvå tusen två hundra man.
Därnäst Benjamins stam: Benjamins barns hövding Abidan, Gideonis son,
med de inmönstrade som utgöra hans här, trettiofem tusen fyra hundra man.
De inmönstrade som tillhöra Efraims läger utgöra alltså tillsammans ett hundra åtta tusen ett hundra man, delade i sina häravdelningar.
Och de skola vid uppbrott tåga i tredje rummet.
Dan skall lägra sig under sitt baner norrut, efter sina häravdelningar: Dans barns hövding Ahieser, Ammisaddais son,
med de inmönstrade som utgöra hans här, sextiotvå tusen sju hundra man.
Bredvid honom skall Asers stam lägra sig: Asers barns hövding Pagiel, Okrans son,
med de inmönstrade som utgöra hans har, fyrtioett tusen fem hundra man.
Därnäst Naftali stam: Naftali barns hövding Ahira, Enans son,
med de inmönstrade som utgöra hans här, femtiotre tusen fyra hundra man.
De inmönstrade som tillhöra Dans läger utgöra alltså tillsammans ett hundra femtiosju tusen sex hundra man.
De skola vid uppbrott tåga sist, under sina baner.
Dessa voro, efter sina familjer, de av Israels barn som inmönstrades.
De som inmönstrades i lägren, efter sina häravdelningar, utgjorde tillsammans sex hundra tre tusen fem hundra femtio man.
Men leviterna blevo icke inmönstrade med de övriga israeliterna, ty så hade HERREN: bjudit Mose.
Och Israels barn gjorde så; alldeles så, som HERREN hade bjudit Mose, lägrade de sig under sina baner, och så tågade de ock, var och en i sin släkt, efter sin familj.
Detta är berättelsen om Arons och Moses släkt, vid den tid då HERREN talade med Mose på Sinai berg.
Dessa äro namnen på Arons söner: Nadab, den förstfödde, och Abihu, Eleasar och Itamar.
Dessa voro namnen på Arons söner, de smorda prästerna, som hade mottagit handfyllning till att vara präster.
Men Nadab och Abihu föllo döda ned inför HERRENS ansikte, när de framburo främmande eld inför HERRENS ansikte i Sinais öken; och de hade inga söner.
Sedan voro Eleasar och Itamar präster under sin fader Aron.
Och HERREN talade till Mose och sade:
Levi stam skall du låta få tillträde hit; du skall låta dem stå inför prästen Aron för att betjäna honom.
De skola iakttaga vad han har att iakttaga, och vad hela menigheten har att iakttaga, inför uppenbarelsetältet, i det att de förrätta tjänsten vid tabernaklet.
Och de skola hava vården om alla uppenbarelsetältets tillbehör, och iakttaga vad Israels barn hava att iakttaga, i det att de förrätta tjänsten vid tabernaklet.
Alltså skall du giva leviterna åt Aron och hans söner; de skola vara honom givna såsom gåva av Israels barn.
Men Aron och hans söner skall du anbefalla att iakttaga vad som hör till deras prästämbete.
Om någon främmande kommer därvid, skall han dödas.
Och HERREN talade till Mose och sade:
Se, jag har själv bland Israels barn uttagit leviterna i stället för allt förstfött bland Israels barn, allt som öppnar moderlivet, så att leviterna skola tillhöra mig.
Ty mig tillhör allt förstfött; på den dag då jag slog allt förstfött i Egyptens land helgade jag åt mig allt förstfött i Israel, såväl människor som boskap.
Mig skola de tillhöra.
Jag är HERREN.
Och HERREN talade till Mose i Sinais öken och sade:
Mönstra Levi barn, efter deras familjer och efter deras släkter; alla av mankön som äro en månad gamla eller därutöver skall du inmönstra.
och Mose inmönstrade dem efter HERRENS befallning, såsom honom hade blivit bjudet.
Och dessa voro Levis söner, efter deras namn: Gerson, Kehat och Merari.
Och dessa voro namnen på Gersons söner, efter deras släkter: Libni och Simei.
Och Kehats söner efter sina släkter voro Amram och Jishar, Hebron och Ussiel.
Och Meraris söner efter sina släkter voro Maheli och Musi.
Dessa voro leviternas släkter, efter deras familjer.
Från Gerson härstammade libniternas släkt och simeiternas släkt; dessa voro gersoniternas släkter.
De av dem som inmönstrades, i det att man räknade alla dem av mankön som voro en månad gamla eller därutöver dessa inmönstrade utgjorde sju tusen fem hundra.
Gersoniternas släkter hade sitt läger bakom tabernaklet, västerut.
Och hövding för gersoniternas stamfamilj var Eljasaf, Laels son.
Och Gersons barn skulle vid uppenbarelsetältet hava vården om själva tabernaklet och dess täckelse, om dess överdrag och om förhänget för ingången till uppenbarelsetältet,
vidare om förgårdens omhängen och om förhänget för ingången till förgården, som omgav tabernaklet och altaret, så ock om dess streck -- vad arbete nu kunde förekomma därvid.
Från Kehat härstammade amramiternas släkt, jishariternas släkt hebroniternas släkt och ussieliternas släkt; dessa voro kehatiternas släkter.
När man räknade alla dem av mankön som voro en månad gamla eller därutöver, utgjorde de åtta tusen sex hundra; dessa voro de som skulle hava vården om de heliga föremålen.
Kehats barns släkter hade sitt läger vid sidan av tabernaklet, söderut.
Och hövding för de kehatitiska släkternas stamfamilj; var Elisafan, Ussiels son.
De skulle hava vården om arken, bordet, ljusstaken, altarna och de tillbehör till de heliga föremålen, som begagnades vid gudstjänsten, så ock om förhänget och om allt arbete därvid.
Men överhövding över alla leviterna var Eleasar, prästen Arons son; han var förman för dem som skulle hava vården om de heliga föremålen.
Från Merari härstammade maheliternas släkt och musiternas släkt; dessa voro merariternas släkter.
Och de av dem som inmönstrades, i det att man räknade alla dem av mankön som voro en månad gamla eller därutöver, utgjorde sex tusen två hundra.
Och hövding för de meraritiska släkternas stamfamilj var Suriel, Abihails son.
De hade sitt läger vid sidan av tabernaklet, norrut.
Och Meraris barn fingo till åliggande att hava vården om bräderna till tabernaklet, om dess tvärstänger, stolpar och fotstycken och om alla dess tillbehör och om allt arbete därvid,
så ock om stolparna till förgården runt omkring med deras fotstycken, deras pluggar och streck.
Men mitt för tabernaklet, på framsidan, mitt för uppenbarelsetältet, österut, hade Mose och Aron och hans söner sitt läger; dessa skulle iakttaga vad som var att iakttaga vid helgedomen, vad Israels barn hade att iakttaga; men om någon främmande kom därvid, skulle han dödas.
De inmönstrade av leviterna som Mose och Aron inmönstrade efter deras släkter, enligt HERRENS befallning, alla av mankön som voro en månad gamla eller därutöver, utgjorde tillsammans tjugutvå tusen.
Och HERREN sade till Mose: Mönstra allt förstfött av mankön bland Israels barn, alla som äro en månad gamla eller därutöver, och räkna antalet av deras namn.
Och tag ut åt mig -- ty jag är HERREN -- leviterna i stället för allt förstfött bland Israels barn, så ock leviternas boskap i stället för allt förstfött bland Israels barns boskap.
Och Mose mönstrade allt förstfött bland Israels barn, såsom HERREN hade bjudit honom.
Och de förstfödde av mankön, vart namn räknat särskilt, de som voro en månad gamla eller därutöver, utgjorde, så många som inmönstrades, tillsammans tjugutvå tusen två hundra sjuttiotre.
Och HERREN talade till Mose och sade:
Du skall uttaga leviterna i stället för allt förstfött bland Israels barn, så ock leviternas boskap i stället för dessas boskap; så att leviterna skola tillhöra mig.
Jag är HERREN.
Men till lösen för de två hundra sjuttiotre personer med vilka antalet av Israels barns förstfödde överstiger leviternas antal,
skall du taga fem siklar för var person; du skall taga upp dessa efter helgedomssikelns vikt, sikeln räknad till tjugu gera.
Och du skall giva penningarna åt Aron och hans söner såsom lösen för de övertaliga bland folket.
Och Mose tog lösesumman av dem som voro övertaliga, när man räknade dem som voro lösta genom leviterna.
Av Israels barns förstfödde tog han penningarna, ett tusen tre hundra sextiofem siklar, efter helgedomssikelns vikt.
Och Mose gav lösesumman åt Aron och hans söner, efter HERRENS befallning, såsom HERREN hade bjudit Mose.
Och HERREN talade till Mose och Aron och sade:
Räknen bland Levi barn antalet av Kehats barn, efter deras släkter och efter deras familjer,
dem som äro trettio år gamla eller därutöver, ända till femtio år, alla tjänstbara män som kunna förrätta sysslor vid uppenbarelsetältet.
Och detta skall vara Kehats barns tjänstgöring vid uppenbarelsetältet: de skola hava hand om de högheliga föremålen.
När lägret skall bryta upp, skola Aron och hans söner gå in och taga ned den förlåt som hänger framför arken och med den övertäcka vittnesbördets ark;
däröver skola de lägga ett överdrag av tahasskinn och över detta ytterligare breda ett kläde, helt och hållet mörkblått; sedan skola de sätta in stängerna.
Och över skådebrödsbordet skola de breda ett mörkblått kläde och ställa därpå faten, skålarna och bägarna, ävensom kannorna till drickoffren; »det beständiga brödet» skall ock läggas därpå.
Häröver skola de breda ett rosenrött kläde och betäcka detta med ett överdrag av tahasskinn; sedan skola de sätta in stängerna.
Och de skola taga ett mörkblått kläde och därmed övertäcka ljusstaken och dess lampor, lamptänger och brickor, så ock alla tillhörande oljekärl som begagnas under tjänstgöringen därvid;
och de skola lägga den med alla dess tillbehör i ett överdrag av tahasskinn och sedan lägga alltsammans på en bår.
Över det gyllene altaret skola de likaledes breda ett mörkblått kläde och betäcka detta med ett överdrag av tahasskinn, sedan skola de sätta in stängerna.
Och de skola taga alla gudstjänstredskap, som begagnas vid tjänstgöringen i helgedomen, och lägga dem i ett mörkblått kläde och betäcka dem med ett överdrag av tahasskinn, och sedan lägga dem på en bår.
Och de skola taga bort askan från altaret och breda över det ett purpurrött kläde
och lägga därpå alla tillbehör som begagnas under tjänstgöringen därvid, fyrfaten, gafflarna, skovlarna och skålarna, korteligen, altarets alla tillbehör; och däröver skola de breda ett överdrag av tahasskinn och så sätta in stängerna.
Sedan nu Aron och hans söner, när lägret skall bryta upp, så hava övertäckt de heliga föremålen och alla tillbehör till dessa heliga föremål, skola därefter Kehats barn komma för att bära; men de må icke röra vid de heliga föremålen, ty då skola de dö.
Detta är vad Kehats barn hava att bära av det som hör till uppenbarelsetältet.
Och Eleasars, prästen Arons sons åliggande skall vara att hava vården om oljan till ljusstaken, om den välluktande rökelsen, om det dagliga spisoffret och om smörjelseoljan; hans åliggande skall vara att hava vården om hela tabernaklet och om allt vad däri är, de heliga föremålen och deras tillbehör.
Och HERREN talade till Mose och Aron och sade:
Låten icke kehatiternas släktgren utrotas ur leviternas stam.
Utan gören på följande sätt med dem, för att de må leva och icke dö, när de nalkas de högheliga föremålen: Aron och hans söner skola gå in och anvisa var och en av dem vad han har att göra eller bära
men själva må de icke gå in och se de heliga föremålen, icke ens ett ögonblick, ty då skola de dö.
Och HERREN talade till Mose och sade:
Räkna ock antalet av Gersons barn, efter deras familjer och efter deras släkter.
Dem som äro trettio år gamla eller därutöver, ända till femtio år, skall du inmönstra, alla tjänstbara män som kunna förrätta arbete vid uppenbarelsetältet.
Detta skall vara gersoniternas släkters tjänstgöring, vad de hava att göra och vad de hava att bära:
de skola bära de tygvåder av vilka tabernaklet bildas, uppenbarelsetältets täckelse, dess överdrag och det överdrag av tahasskinn som ligger ovanpå detta, förhänget för ingången till uppenbarelsetältet,
vidare omhängena till förgården, förhänget för porten till förgården, som omgiver tabernaklet och altaret, så ock tillhörande streck och alla redskap till arbetet därvid; och allt som härvid är att göra skola de förrätta.
På det sätt Aron och hans söner bestämma skall Gersons barns hela tjänstgöring försiggå, i fråga om allt vad de hava att bära och göra; och I skolen överlämna i deras vård allt vad de hava att bära.
Detta är den tjänstgöring som Gersons barns släkter skola hava vid uppenbarelsetältet; och vad de hava att iakttaga skola de utföra under ledning av Itamar, prästen Arons son
Meraris barn skall du inmönstra, efter deras släkter och efter deras familjer.
Dem som äro trettio år gamla eller därutöver, ända till femtio år, skall du inmönstra, alla tjänstbara män som kunna förrätta arbete vid uppenbarelsetältet.
Och detta är vad som skall åligga dem att bära, allt vad som hör till deras tjänstgöring vid uppenbarelsetältet: bräderna till tabernaklet, dess tvärstänger, stolpar och fotstycken,
så ock stolparna till förgården runt omkring med deras fotstycken, pluggar och streck, korteligen, alla deras tillbehör och allt som hör till arbetet därvid; och I skolen lämna dem uppgift på de särskilda föremål som det åligger dem att bära.
Detta skall vara de meraritiska släkternas tjänstgöring, allt vad som hör till deras tjänstgöring vid uppenbarelsetältet; och det skall utföras under ledning av Itamar, prästen Arons son.
Och Mose och Aron och menighetens hövdingar inmönstrade Kehats barn, efter deras släkter och efter deras familjer,
dem som voro trettio år gamla eller därutöver, ända till femtio år alla tjänstbara män som kunde göra arbete vid uppenbarelsetältet.
Och de av dem som inmönstrades, efter deras släkter, utgjorde två tusen sju hundra femtio.
Så många voro de av kehatiternas släkter som inmönstrades, summan av dem som skulle göra tjänst vid uppenbarelsetältet, de som Mose och Aron inmönstrade, efter HERRENS befallning genom Mose.
Och de av Gersons barn som inmönstrades, efter deras släkter och efter deras familjer,
de som voro trettio år gamla eller därutöver, ända till femtio år, alla tjänstbara män som kunde göra arbete vid uppenbarelsetältet,
dessa som inmönstrades efter sina släkter och efter sina familjer utgjorde två tusen sex hundra trettio.
Så många voro de av Gersons barns släkter som inmönstrades, summan av dem som skulle göra tjänst vid uppenbarelsetältet, de som Mose och Aron inmönstrade, efter HERRENS befallning.
Och de av Meraris barns släkter som inmönstrades, efter deras släkter och efter deras familjer,
de som voro trettio år gamla eller därutöver, ända till femtio år, alla tjänstbara män som kunde göra arbete vid uppenbarelsetältet,
dessa som inmönstrades efter sina släkter utgjorde tre tusen två hundra.
Så många voro de av Meraris barns släkter som inmönstrades, de som Mose och Aron inmönstrade efter HERRENS befallning genom Mose.
De av leviterna som Mose och Aron och Israels hövdingar inmönstrade, efter deras släkter och efter deras familjer,
de som voro trettio år gamla eller därutöver, ända till femtio år, alla som kunde förrätta något tjänstgöringsarbete eller något bärarearbete vid uppenbarelsetältet,
dessa som inmönstrades utgjorde tillsammans åtta tusen fem hundra åttio.
Efter HERRENS befallning blevo de inmönstrade genom Mose, var och en till det som han hade att göra eller bära, och var och en fick det åliggande som HERREN hade bjudit Mose.
Och HERREN talade till Mose och sade:
Bjud Israels barn att de skaffa bort ur lägret var och en som är spetälsk eller har flytning och var och en som har blivit oren genom någon död.
En sådan, vare sig man eller kvinna, skolen I skaffa bort; till något ställe utanför lägret skolen I skicka honom, för att han icke må orena deras läger; jag har ju min boning mitt ibland dem.
Och Israels barn gjorde så; de skickade dem till ett ställe utanför lägret; såsom HERREN hade tillsagt Mose, så gjorde Israels barn.
Och HERREN talade till Mose och sade:
Tala till Israels barn: Om någon, vare sig man eller kvinna, begår någon synd -- vad det nu må vara, vari en människa kan försynda sig -- i det han gör sig skyldig till en orättrådighet mot HERREN, och denna person alltså ådrager sig skuld,
så skall han bekänna den synd han har begått, och ersätta det han har förbrutit sig på till dess fulla belopp och lägga femtedelen av värdet därtill; och detta skall han giva åt den som han har förbrutit sig emot.
Men om denne icke har efterlämnat någon bördeman, åt vilken ersättning kan givas för det han har förbrutit sig på, då skall ersättningen för detta givas åt HERREN och tillhöra prästen, utom försoningsväduren, med vilken försoning bringas för den skyldige.
Och alla heliga gåvor som Israels barn giva såsom en gärd, vilken de bära fram till prästen, skola tillhöra denne;
honom skola allas heliga gåvor tillhöra; vad någon giver åt prästen skall tillhöra denne.
Och HERREN talade till Mose och sade:
Tala till Israels barn och säg till dem: Om en hustru har svikit sin man och varit honom otrogen,
i det att någon annan har legat hos henne och beblandat sig med henne, utan att hennes man har fått veta därav, och utan att hon har blivit röjd, fastän hon verkligen har låtit skända sig; om alltså intet vittne finnes mot henne och hon icke har blivit gripen på bar gärning,
men misstankens ande likväl kommer över honom, så att han får misstanke mot sin hustru, och det verkligen är så, att hon har låtit skända sig; eller om misstankens ande kommer över honom, så att han får misstanke mot sin hustru, och detta fastän hon icke har låtit skända sig:
så skall mannen föra sin hustru till prästen och såsom offer för henne bära fram en tiondedels efa kornmjöl, men ingen olja skall han gjuta därpå och ingen rökelse lägga därpå, ty det är ett misstankeoffer, ett åminnelseoffer, som bringar en missgärning i åminnelse.
Och prästen skall föra henne fram och ställa henne inför HERRENS ansikte.
Och prästen skall taga heligt vatten i ett lerkärl, och sedan skall prästen taga något av stoftet på tabernaklets golv och lägga i vattnet.
Och prästen skall ställa kvinnan fram inför HERRENS ansikte och lösa upp kvinnans hår och lägga på hennes händer åminnelseoffret, det är misstankeoffret; men prästen själv skall hålla i sin hand det förbannelsebringande olycksvattnet.
Därefter skall prästen besvärja kvinnan och säga till henne: »Om ingen har lägrat dig och du icke har svikit din man genom att låta skända dig, så må detta förbannelsebringande olycksvatten icke skada dig.
Men om du har svikit din man och låtit skända dig, i det att någon annan än din man har beblandat sig med dig»
(prästen besvärjer nu kvinnan med förbannelsens ed, i det han säger till kvinnan:) »Då må HERREN göra dig till ett exempel som man nämner, när man förbannar och svär bland ditt folk; HERREN må då låta din länd förvissna och din buk svälla upp;
ja, när du har fått detta förbannelsebringande vatten in i ditt liv, då må det komma din buk att svälla upp och din länd att förvissna.»
Och kvinnan skall säga: »Amen, amen.»
Sedan skall prästen skriva upp dessa förbannelser på ett blad och därefter avtvå dem i olycksvattnet
och giva kvinnan det förbannelsebringande olycksvattnet att dricka, för att detta förbannelsebringande vatten må bliva henne till olycka, när hon har fått det i sig.
Och prästen skall taga misstankeoffret ur kvinnans hand och vifta detta offer inför HERRENS ansikte och bära det fram till altaret.
Och prästen skall av offret taga en handfull, det som utgör själva altaroffret, och förbränna det på altaret; därefter skall han giva kvinnan vattnet att dricka.
Och när han så har givit henne vattnet att dricka, då skall detta ske: om hon har låtit skända sig och varit sin man otrogen, så skall det förbannelsebringande vattnet, när hon har fått det i sig, bliva henne till olycka, i det att hennes buk sväller upp och hennes länd förvissnar; och kvinnan skall bliva ett exempel som man nämner, när man förbannar bland hennes folk.
Men om kvinnan icke har låtit skända sig, utan är ren, då skall hon förbliva oskadd och kunna undfå livsfrukt.
Detta är misstankelagen, om huru förfaras skall, när en kvinna har svikit sin man och låtit skända sig,
eller när eljest misstankens ande kommer över en man, så att han misstänker sin hustru; han skall då ställa hustrun fram inför HERRENS ansikte, och prästen skall med henne göra allt vad denna lag stadgar.
Så skall mannen vara fri ifrån missgärning, men hustrun kommer att bära på missgärning.
Och HERREN talade till Mose och sade:
Tala till Israels barn och säg till dem: Om någon, vare sig man eller kvinna, har att fullgöra ett nasirlöfte, ett löfte att vara HERRENS nasir,
så skall han avhålla sig från vin och starka drycker; han skall icke dricka någon syrad dryck av vin eller någon annan syrad stark dryck; intet slags druvsaft skall han dricka, ej heller skall han äta druvor, vare sig friska eller torra.
Så länge hans nasirtid varar, skall han icke äta något som kommer av vinträdet, icke ens dess kartar eller späda skott.
Så länge hans nasirlöfte varar, skall ingen rakkniv komma på hans huvud; till dess att den tid är ute, under vilken han skall vara HERRENS nasir, skall han vara helig och låte håret växa långt på sitt huvud.
Så länge han är HERRENS nasir, skall han icke nalkas någon död.
Icke ens genom sin fader eller sin moder, sin broder eller sin syster får han ådraga sig orenhet, om de dö ty han bär på sitt huvud tecknet till att han är sin Guds nasir;
så länge hans nasirtid varar, är han helgad åt HERREN.
Men om någon oförtänkt och plötsligt dör i hans närhet, och därmed orenar hans huvud, på vilket han bär nasirtecknet, så skall han raka sitt huvud den dag han bliver ren; han skall raka det på sjunde dagen.
Och på åttonde dagen skall han bära fram till prästen två turturduvor eller två unga duvor, till uppenbarelsetältets ingång.
Och prästen skall offra en till syndoffer och en till brännoffer och bringa försoning för honom, till rening från den synd han har dragit över sig genom den döde; sedan skall han samma dag åter helga sitt huvud;
han skall inviga sig till nasir åt HERREN för lika lång tid som han förut hade lovat.
Och han skall föra fram ett årsgammalt lamm till skuldoffer.
Den förra löftestiden skall vara ogill, därför att hans nasirat blev orenat.
Och detta är lagen om en nasir: Den dag hans nasirtid är ute skall han föras fram till uppenbarelsetältets ingång;
och han skall såsom sitt offer åt HERREN frambära ett årsgammalt felfritt lamm av hankön till brännoffer och ett årsgammalt felfritt lamm av honkön till syndoffer och en felfri vädur till tackoffer,
därjämte en korg med osyrat bröd, kakor av fint mjöl, begjutna med olja, och osyrade tunnkakor, smorda med olja, så ock tillhörande spis offer och drickoffer.
Och prästen skall bära fram detta inför HERRENS ansikte och offra hans syndoffer och hans brännoffer.
Och väduren skall han offra till tackoffer åt HERREN, jämte korgen med de osyrade bröden; prästen skall ock offra tillhörande spisoffer och drickoffer.
Och nasiren skall vid ingången till uppenbarelsetältet raka sitt huvud, på vilket han bär nasirtecknet, och taga sitt huvudhår, sitt nasirtecken, och lägga det på elden som brinner under tackoffret.
Och prästen skall taga den kokta vädursbogen, och därjämte ur korgen en osyrad kaka och en osyrad tunnkaka, och lägga detta på nasirens händer, sedan denne har rakat av sig nasirtecknet.
Och prästen skall vifta detta såsom ett viftoffer inför HERRENS ansikte; det skall vara helgat åt prästen, jämte viftoffersbringan och offergärdslåret.
Sedan får nasiren åter dricka vin.
Detta är lagen om den som har avlagt ett nasirlöfte, och om vad han på grund av nasirlöftet skall offra åt HERREN, förutom vad han eljest kan anskaffa; efter innehållet i det löfte han har avlagt skall han göra, enligt lagen om hans nasirat.
Och HERREN talade till Mose och sade:
Tala till Aron och hans söner och säg: När I välsignen Israels barn, skolen I säga så till dem:
HERREN välsigne dig och bevare dig.
HERREN låte sitt ansikte lysa över dig och vare dig nådig.
HERREN vände sitt ansikte till dig och give dig frid.
Så skola de lägga mitt namn på Israels barn, och jag skall då välsigna dem.
Då nu Mose hade satt upp tabernaklet och smort och helgat det, med alla dess tillbehör, och hade satt upp altaret med alla dess tillbehör, och smort och helgat detta,
framburos offergåvor av Israels hövdingar, huvudmännen för stamfamiljerna, det är stamhövdingarna, som stodo i spetsen för de inmönstrade.
De förde fram såsom sin offergåva inför HERRENS ansikte sex övertäckta vagnar och tolv oxar: två hövdingar tillhopa en vagn och var hövding en oxe; dessa förde de fram inför tabernaklet.
Och HERREN sade till Mose:
»Tag emot detta av dem för att bruka det till uppenbarelsetältets tjänst; och lämna det åt leviterna, alltefter beskaffenheten av vars och ens tjänst.»
Och Mose tog emot vagnarna och oxarna och gav dem åt leviterna.
Två vagnar och fyra oxar gav han åt Gersons barn, efter beskaffenheten av deras tjänst;
fyra vagnar och åtta oxar gav han åt Meraris barn, efter beskaffenheten av den tjänst de förrättade under ledning av Itamar, prästen Arons son;
men åt Kehats barn gav han icke något, ty dem ålåg att hava hand om de heliga föremålen, och dessa skulle bäras på axlarna.
Och hövdingarna förde fram skänker till altarets invigning, när det smordes; hövdingarna förde fram dessa sina offergåvor inför altaret.
Och HERREN sade till Mose: »Låt hövdingarna, en i sänder, var och en på sin dag, föra fram sina offergåvor till altarets invigning.»
Och den som på första dagen förde fram sin offergåva var Naheson, Amminadabs son, av Juda stam
Hans offergåva var ett silverfat, ett hundra trettio siklar i vikt, och en silverskål om sjuttio siklar, efter helgedomssikelns vikt, båda fulla med fint mjöl, begjutet med olja, till spisoffer,
vidare en skål av guld om tio siklar, full med rökelse,
vidare en ungtjur, en vädur och ett årsgammalt lamm till brännoffer
och en bock till syndoffer,
samt till tackoffret två tjurar, fem vädurar, fem bockar och fem årsgamla lamm.
Detta var Nahesons, Amminadabs sons, offergåva.
På andra dagen förde Netanel, Suars son, hövdingen för Isaskar, fram sin gåva;
han framförde såsom sin offergåva ett silverfat, ett hundra trettio siklar i vikt, och en silverskål om sjuttio siklar, efter helgedomssikelns vikt, båda fulla med fint mjöl, begjutet med olja, till spisoffer,
vidare en skål av guld om tio siklar, full med rökelse,
vidare en ungtjur, en vädur och ett årsgammalt lamm till brännoffer
och en bock till syndoffer,
samt till tackoffret två tjurar, fem vädurar, fem bockar och fem årsgamla lamm.
Detta var Netanels, Suars sons, offergåva.
På tredje dagen kom hövdingen för Sebulons barn, Eliab, Helons son;
hans offergåva var ett silverfat, ett hundra trettio siklar i vikt, och en silverskål om sjuttio siklar, efter helgedomssikelns vikt, båda fulla med fint mjöl, begjutet med olja, till spisoffer
vidare en skål av guld om tio siklar, full med rökelse,
vidare en ungtjur, en vädur och ett årsgammalt lamm till brännoffer
och en bock till syndoffer,
samt till tackoffret två tjurar, fem vädurar, fem bockar och fem årsgamla lamm.
Detta var Eliabs, Helons sons, offergåva.
På fjärde dagen kom hövdingen för Rubens barn, Elisur, Sedeurs son;
hans offergåva var ett silverfat, ett hundra trettio siklar i vikt, och en silverskål om sjuttio siklar, efter helgedomssikelns vikt, båda fulla med fint mjöl, begjutet med olja, till spisoffer,
vidare en skål av guld om tio siklar, full med rökelse,
vidare en ungtjur, en vädur och ett årsgammalt lamm till brännoffer
och en bock till syndoffer,
samt till tackoffret två tjurar, fem vädurar, fem bockar och fem årsgamla lamm.
Detta var Elisurs, Sedeurs sons, offergåva.
På femte dagen kom hövdingen för Simeons barn, Selumiel, Surisaddais son;
hans offergåva var ett silverfat, ett hundra trettio siklar i vikt, och en silverskål om sjuttio siklar, efter helgedomssikelns vikt, båda fulla med fint mjöl, begjutet med olja, till spisoffer,
vidare en skål av guld om tio siklar, full med rökelse,
vidare en ungtjur, en vädur och ett årsgammalt lamm till brännoffer
och en bock till syndoffer,
samt till tackoffret två tjurar, fem vädurar, fem bockar och fem årsgamla lamm.
Detta var Selumiels, Surisaddais sons, offergåva.
På sjätte dagen kom hövdingen för Gads barn, Eljasaf, Deguels son;
hans offergåva var ett silverfat, ett hundra trettio siklar i vikt, och en silverskål om sjuttio siklar, efter helgedomssikelns vikt, båda fulla med fint mjöl, begjutet med olja, till spisoffer,
vidare en skål av guld om tio siklar, full med rökelse,
vidare en ungtjur, en vädur och ett årsgammalt lamm till brännoffer
och en bock till syndoffer,
samt till tackoffret två tjurar, fem vädurar, fem bockar och fem årsgamla lamm.
Detta var Eljasafs, Deguels sons, offergåva.
På sjunde dagen kom hövdingen för Efraims barn, Elisama, Ammihuds son;
hans offergåva var ett silverfat, ett hundra trettio siklar i vikt, och en silverskål om sjuttio siklar, efter helgedomssikelns vikt, båda fulla med fint mjöl, begjutet med olja, till spisoffer,
vidare en skål av guld om tio siklar, full med rökelse,
vidare en ungtjur, en vädur och ett årsgammalt lamm till brännoffer
och en bock till syndoffer,
samt till tackoffret två tjurar, fem vädurar, fem bockar och fem årsgamla lamm.
Detta var Elisamas, Ammihuds sons, offergåva.
På åttonde dagen kom hövdingen för Manasse barn, Gamliel, Pedasurs son;
hans offergåva var ett silverfat, ett hundra trettio siklar i vikt, och en silverskål om sjuttio siklar, efter helgedomssikelns vikt, båda fulla med fint mjöl, begjutet med olja, till spisoffer,
vidare en skål av guld om tio siklar, full med rökelse,
vidare en ungtjur en vädur och ett årsgammalt lamm till brännoffer
och en bock till syndoffer,
samt till tackoffret två tjurar, fem vädurar, fem bockar och fem årsgamla lamm.
Detta var Gamliels Pedasurs sons, offergåva.
På nionde dagen kom hövdingen för Benjamins barn, Abidan, Gideonis son;
hans offergåva var ett silverfat, ett hundra trettio siklar i vikt, och en silverskål om sjuttio siklar, efter helgedomssikelns vikt, båda fulla med fint mjöl, begjutet med olja, till spisoffer,
vidare en skål av guld om tio siklar, full med rökelse,
vidare en ungtjur, en vädur och ett årsgammalt lamm till brännoffer
och en bock till syndoffer,
samt till tackoffret två tjurar, fem vädurar, fem bockar och fem årsgamla lamm.
Detta var Abidans, Gideonis sons, offergåva.
På tionde dagen kom hövdingen för Dans barn, Ahieser, Ammisaddais son;
hans offergåva var ett silverfat, ett hundra trettio siklar i vikt, och en silverskål om sjuttio siklar, efter helgedomssikelns vikt, båda fulla med fint mjöl, begjutet med olja, till spisoffer,
vidare en skål av guld om tio siklar, full med rökelse,
vidare en ungtjur, en vädur och ett årsgammalt lamm till brännoffer
och en bock till syndoffer,
samt till tackoffret två tjurar, fem vädurar, fem bockar och fem årsgamla lamm.
Detta var Ahiesers, Ammisaddais sons, offergåva.
På elfte dagen kom hövdingen för Asers barn, Pagiel, Okrans son;
hans offergåva var ett silverfat, ett hundra trettio siklar i vikt, och en silverskål om sjuttio siklar, efter helgedomssikelns vikt, båda fulla med fint mjöl, begjutet med olja, till spisoffer,
vidare en skål av guld om tio siklar, full med rökelse,
vidare en ungtjur, en vädur och ett årsgammalt lamm till brännoffer
och en bock till syndoffer,
samt till tackoffret två tjurar, fem vädurar, fem bockar och fem årsgamla lamm.
Detta var Pagiels, Okrans sons, offergåva.
På tolfte dagen kom hövdingen för Naftali barn, Ahira, Enans son;
hans offergåva var ett silverfat, ett hundra trettio siklar i vikt, och en silverskål om sjuttio siklar, efter helgedomssikelns vikt, båda fulla med fint mjöl, begjutet med olja, till spisoffer,
vidare en skål av guld om tio siklar, full med rökelse,
vidare en ungtjur, en vädur och ett årsgammalt lamm till brännoffer
och en bock till syndoffer,
samt till tackoffret två tjurar, fem vädurar, fem bockar och fem årsgamla lamm.
Detta var Ahiras, Enans sons, offergåva.
Detta var vad Israels hövdingar skänkte till altarets invigning, när det smordes: tolv silverfat, tolv silverskålar och tolv guldskålar.
Vart fat kom på ett hundra trettio silversiklar och var skål på sjuttio siklar, så att silvret i dessa kärl sammanlagt utgjorde två tusen fyra hundra siklar, efter helgedomssikelns vikt.
Av de tolv guldskålarna, som voro fulla med rökelse, vägde var och en tio siklar, efter helgedomssikelns vikt, så att guldet i skålarna sammanlagt utgjorde ett hundra tjugu siklar.
Brännoffers-fäkreaturen utgjorde tillsammans tolv tjurar, vartill kommo tolv vädurar, tolv årsgamla lamm, med tillhörande spisoffer, och tolv bockar till syndoffer.
Och tackoffers-fäkreaturen utgjorde tillsammans tjugufyra tjurar, vartill kommo sextio vädurar, sextio bockar och sextio årsgamla lamm.
Detta var vad som skänktes till altarets invigning, sedan det hade blivit smort.
Och när Mose gick in i uppenbarelsetältet för att tala med honom, hörde han rösten tala till sig från nådastolen ovanpå vittnesbördets ark, från platsen mellan de två keruberna; där talade rösten till honom.
Och HERREN talade till Mose och sade:
»Tala till Aron och säg till honom: När du sätter upp lamporna, skall detta ske så, att de sju lamporna kasta sitt sken över platsen framför ljusstaken.»
Och Aron gjorde så; han satte upp lamporna så, att de kastade sitt sken över platsen framför ljusstaken, såsom HERREN hade bjudit Mose.
Och ljusstaken var gjord på följande sätt: den var av guld i drivet arbete; också dess fotställning och blommorna därpå voro i drivet arbete.
Efter det mönster som HERREN hade visat Mose hade denne låtit göra ljusstaken.
Och HERREN talade till Mose och sade:
Du skall bland Israels barn uttaga leviterna och rena dem.
Och på följande sätt skall du göra med dem för att rena dem: Du skall stänka reningsvatten på dem; och de skola låta raka hela sin kropp och två sina kläder och skola så rena sig.
Sedan skola de taga en ungtjur, med tillhörande spisoffer av fint mjöl, begjutet med olja; därjämte skall du taga en annan ungtjur till syndoffer.
Och du skall föra leviterna fram inför uppenbarelsetältet, och du skall församla Israels barns hela menighet
Och när du har fört leviterna fram inför HERRENS ansikte, skola Israels barn lägga sina händer på dem.
Och Aron skall vifta leviterna inför HERRENS ansikte såsom ett viftoffer från Israels barn, och de skola sedan hava till åliggande att förrätta HERRENS tjänst.
Och leviterna skola lägga sina händer på tjurarnas huvuden, och den ena skall du offra till syndoffer och den andra till brännoffer åt HERREN, för att bringa försoning för leviterna.
Så skall du ställa leviterna inför Aron och hans söner och vifta dem såsom ett viftoffer åt HERREN.
På detta sätt skall du bland Israels barn avskilja leviterna, så att leviterna skola tillhöra mig.
Därefter skola leviterna gå in och göra tjänst vid uppenbarelsetältet, sedan du har renat dem och viftat dem såsom ett viftoffer;
ty bland Israels barn äro de givna åt mig såsom gåva; i stället för allt som öppnar moderlivet, allt förstfött bland Israels barn, har jag uttagit dem åt mig.
Ty mig tillhör allt förstfött bland, Israels barn, både människor och boskap; på den dag då jag slog allt förstfött i Egyptens land helgade jag det åt mig.
Och jag har tagit leviterna i stället för allt förstfött bland Israels barn.
Och jag har bland Israels barn givit leviterna såsom gåva åt Aron och hans söner, till att förrätta Israels barns tjänst vid uppenbarelsetältet och bringa försoning för Israels barn, på det att ingen hemsökelse må drabba Israels barn, därigenom att Israels barn nalkas helgedomen.
Och Mose och Aron och Israels barns hela menighet gjorde så med leviterna; Israels barn gjorde med leviterna i alla stycken såsom HERREN hade bjudit Mose angående dem.
Och leviterna renade sig och tvådde sina kläder, och Aron viftade dem såsom ett viftoffer inför HERRENS ansikte, och Aron bragte försoning för dem och renade dem.
Därefter gingo leviterna in och förrättade sin tjänst vid uppenbarelsetältet under Aron och hans söner.
Såsom HERREN hade bjudit Mose angående leviterna, så gjorde de med dem.
och HERREN talade till Mose och sade:
Detta är vad som skall gälla angående leviterna: Den som är tjugufem år gammal eller därutöver skall infinna sig och göra tjänst med arbete vid uppenbarelsetältet.
Men när leviten bliver femtio år gammal, skall han vara fri ifrån att tjäna med arbete; han skall då icke längre arbeta.
Han må betjäna sina bröder vid uppenbarelsetältet med att iakttaga vad som där är att iakttaga; men något bestämt arbete skall han icke förrätta.
Så skall du förfara med leviterna i vad som angår deras åligganden.
Och HERREN talade till Mose Sinais öken, i första månaden av det andra året efter deras uttåg ur Egyptens land; han sade:
Israels barn skola ock hålla påsk högtid på den bestämda tiden.
På fjortonde dagen i denna månad, vid aftontiden, skolen I hålla den, på bestämd tid.
Enligt alla stadgar och föreskrifter därom skolen I hålla den.
Så sade då Mose till Israels barn att de skulle hålla påskhögtid.
Och de höllo påskhögtid i först månaden, på fjortonde dagen i månaden, vid aftontiden, i Sinais öken Israels barn gjorde i alla stycken såsom HERREN hade bjudit Mose
Men där voro några män som hade blivit orena genom en död människa, så att de icke kunde hålla påskhögtid på den dagen; dessa trädde på den dagen fram inför Mose och Aron.
Och männen sade till honom: »Vi hava blivit orena genom en död människa; skall det därför förmenas oss att bland Israels barn bära fram HERRENS offergåva på bestämd?»
Mose svarade dem: »Stannen så vill jag höra vad HERREN bjuder angående eder.»
Och HERREN talade till Mose och sade:
Tala till Israels barn och säg: Om någon bland eder eller edra efterkommande har blivit oren genom en död, eller är ute på resa långt borta, och han ändå vill hålla HERRENS påskhögtid
så skall han hålla den i andra månaden, på fjortonde dagen, vid aftontiden.
Med osyrat bröd och bittra örter skall han äta påskalammet.
Intet därav skall lämnas kvar till morgonen, och intet ben skall sönderslås därpå.
I alla stycken skall påskhögtiden hållas såsom stadgat är därom.
Men om någon som är ren, och som icke är ute på resa ändå underlåter att hålla påskhögtid, så skall han utrotas ur sin släkt, eftersom han icke har burit fram HERRENS offergåva på bestämd tid; den mannen bär på synd.
Och om någon främling bor hos eder och vill hålla HERRENS påskhögtid, så skall han hålla den enligt den stadga och föreskrift som gäller för påskhögtiden.
En och samma stadga skall gälla för eder, lika väl för främlingen som för infödingen i landet.
Och på den dag då tabernaklet sattes upp övertäckte molnskyn tabernaklet, vittnesbördets tält, och om aftonen, och sedan ända till morgonen, var det såsom såge man en eld över tabernaklet.
Så var det beständigt: molnskyn övertäckte det, och om natten var det såsom såge man en eld.
Och så ofta molnskyn höjde sig från tältet, bröto Israels barn strax upp, och på det ställe där molnskyn stannade, där slogo Israels barn läger.
Efter HERRENS befallning bröto Israels barn upp, och efter HERRENS befallning slogo de läger.
Så länge molnskyn vilade över tabernaklet, lågo de i läger.
Och om molnskyn en längre tid förblev över tabernaklet, så iakttogo Israels barn vad HERREN bjöd dem iakttaga och bröto icke upp.
Stundom kunde det hända att molnskyn allenast några få dagar stannade över tabernaklet; då lågo de efter HERRENS befallning i läger och bröto sedan upp efter HERRENS befallning.
Stundom kunde det ock hända att molnskyn stannade allenast från aftonen till morgonen; när då molnskyn om morgonen höjde sig, bröto de upp; eller om så var, att molnskyn stannade en dag och en natt och sedan höjde sig, så bröto de upp då.
Eller om den stannade två dagar, eller en månad, eller vilken tid som helst, så att molnskyn länge förblev vilande över tabernaklet, så lågo Israels barn stilla i läger och bröto icke upp; men när den sedan höjde sig, bröto de upp.
Efter HERRENS befallning slogo de läger, och efter HERRENS befallning bröto de upp.
Vad HERREN bjöd dem iakttaga, det iakttogo de, efter HERRENS befallning genom Mose.
Och HERREN talade till Mose och sade:
»Gör dig två trumpeter av silver; i drivet arbete skall du göra dem.
Dessa skall du bruka, när menigheten skall sammankallas, och när lägren skola bryta upp.
När man stöter i dem båda, skall hela menigheten församla sig till dig, vid ingången till uppenbarelsetältet.
Men när man stöter allenast i den ena, skola hövdingarna, huvudmännen för Israels ätter, församla sig till dig.
Och när I blåsen en larmsignal, skola de läger bryta upp, som ligga österut.
Men när I blåsen larmsignal för andra gången, skola de läger bryta upp, som ligga söderut.
När lägren skola bryta upp, skall man blåsa larmsignal,
men när församlingen skall sammankallas, skolen I icke blåsa larmsignal, utan stöta i trumpeterna.
Och Arons söner, prästerna, äro de som skola blåsa i trumpeterna.
Detta skall vara en evärdlig stadga för eder från släkte till släkte.
Och om I, i edert land, dragen ut till strid mot någon eder ovän som angriper eder, så skolen I blåsa larmsignal med trumpeterna; härigenom skolen I då bringas i åminnelse inför HERRENS, eder Guds, ansikte, och I skolen så bliva frälsta ifrån edra fiender.
Och när I haven en glädjedag och haven edra högtider och nymånader, skolen I stöta i trumpeterna, då I offren edra brännoffer och tackoffer; så skola de bringa eder i åminnelse inför eder Guds ansikte.
Jag är HERREN, eder Gud.»
I andra året, i andra månaden, på tjugonde dagen i månaden höjde sig molnskyn från vittnesbördets tabernakel.
Då bröto Israels barn upp från Sinais öken och tågade från lägerplats till lägerplats; och molnskyn stannade i öknen Paran.
Och när de nu första gången bröto upp, efter HERRENS befallning genom Mose,
var Juda barns läger under sitt baner det första som bröt upp, häravdelning efter häravdelning; och anförare för denna här var Naheson, Amminadabs son.
Och anförare för den här som utgjordes av Isaskars barns stam var Netanel, Suars son.
Och anförare för den här som utgjordes av Sebulons barns stam var Eliab, Helons son.
Därefter, sedan tabernaklet hade blivit nedtaget, bröto Gersons barn och Meraris barn upp och buro tabernaklet.
Därefter bröt Rubens läger upp under sitt baner, häravdelning efter häravdelning; och anförare för denna här var Elisur, Sedeurs son.
Och anförare för den här som utgjordes av Simeons barns stam var Selumiel, Surisaddais son.
Och anförare för den här som utgjordes av Gads barns stam var Eljasaf, Deguels son.
Därefter bröto kehatiterna upp och buro de heliga tingen, och de andra satte upp tabernaklet, innan dessa hunno fram.
Därefter bröt Efraims barns läger upp under sitt baner, häravdelning efter häravdelning; och anförare för denna här var Elisama, Ammihuds son.
Och anförare för den här som utgjordes av Manasse barns stam var Gamliel, Pedasurs son.
Och anförare for den här som utgjordes av Benjamins barns stam var Abidan, Gideonis son.
Därefter bröt Dans barns läger upp under sitt baner, såsom eftertrupp i hela lägertåget, häravdelning efter häravdelning; och anförare för denna här var Ahieser, Ammisaddais son.
Och anförare för den här som utgjordes av Asers barns stam var Pagiel, Okrans son.
Och anförare för den här som utgjordes av Naftali barns stam var Ahira, Enans son.
I denna ordning bröto Israels barn upp, häravdelning efter häravdelning.
Och de bröto nu upp.
Och Mose sade till Hobab, som var son till midjaniten Reguel, Moses svärfader: »Vi bryta nu upp och tåga till det land om vilket HERREN har sagt: 'Det vill jag giva eder.'
Följ du med oss, så vilja vi göra dig gott, ty HERREN har lovat Israel vad gott är.
Men han svarade honom: »Jag vill icke följa med, utan jag vill gå hem till mitt land och till min släkt.»
Då sade han: »Ack nej, övergiv oss icke.
Du vet ju bäst var vi kunna lägra oss i öknen; bliv du därför nu vårt öga.
Om du följer med oss, skola vi låta också dig få gott av det goda som HERREN gör mot oss.
Så bröto de upp och tågade från HERRENS berg tre dagsresor.
Och HERRENS förbundsark gick framför dem tre dagsresor, för att utse viloplats åt dem.
Och HERRENS molnsky svävade över dem om dagen, när de bröto upp från sitt lägerställe.
Och så ofta arken bröt upp, sade Mose: »Stå upp, HERRE; må dina fiender varda förskingrade, och må de som hata dig fly för ditt ansikte.»
Och när den sattes ned, sade han: »Kom tillbaka, HERRE, till Israels ätters mångtusenden.»
Men folket knorrade, och detta misshagade HERREN.
Ty när HERREN hörde det, upptändes hans vrede, och HERRENS eld begynte brinna ibland dem och förtärde de som voro ytterst i lägret.
Då ropade folket till Mose, och Mose bad till HERREN, och så stannade elden av.
Och detta ställe fick namnet Tabeera, därför att HERRENS eld hade brunnit ibland dem.
Och den blandade folkhop som åtföljde dem greps av lystnad; Israels barn själva begynte då ock åter att gråta och sade: »Ack om vi hade kött att äta!
Vi komma ihåg fisken som vi åt i Egypten för intet, så ock gurkorna, melonerna, purjolöken, rödlöken och vitlöken.
Men nu försmäkta våra själar, ty här finnes alls intet; vi få intet annat se än manna.
Men mannat liknade korianderfrö och hade samma utseende som bdelliumharts.
Folket gick omkring och samlade sådant, och malde det därefter på handkvarn eller stötte sönder det i mortel, och kokte det sedan i gryta och bakade kakor därav; och det smakade såsom fint bakverk med olja.
När daggen om natten föll över lägret, föll ock mannat där.
Och Mose hörde huru folket i sina särskilda släkter grät, var och en vid ingången till sitt tält; och HERRENS vrede upptändes storligen, och Mose själv blev misslynt.
Och Mose sade till HERREN: »Varför har du gjort så illa mot din tjänare, och varför har jag så litet funnit nåd för dina ögon, att du har lagt på mig bördan av hela detta folk?
Är då jag moder eller fader till hela detta folk, eftersom du säger till mig att jag skall bära det i min famn, såsom spenabarnet bäres av sin vårdare, in i det land som du med ed har lovat åt deras fäder?
Varifrån skall jag få kött att giva åt hela detta folk?
De gråta ju och vända sig mot mig och säga: 'Giv oss kött, så att vi få äta.'
Jag förmår icke ensam bära hela detta folk, ty det bliver mig för tungt.
Vill du så handla mot mig, så dräp mig hellre med ens, om jag har funnit nåd för dina ögon, och låt mig slippa detta elände.»
Då sade HERREN till Mose: »Samla ihop åt mig sjuttio män av de äldste i Israel, dem som du vet höra till de äldste i folket och till dess tillsyningsmän; och för dessa fram till uppenbarelsetältet och låt dem ställa sig där hos dig.
Där vill jag då stiga ned och tala med dig, och jag vill taga av den ande som är över dig och låta komma över dem; sedan skola de bistå dig med att bära på bördan av folket, så att du slipper bära den ensam.
Och till folket skall du säga: Helgen eder till i morgon, så skolen I få kött att äta, eftersom I haven gråtit inför HERREN och sagt: 'Ack om vi hade kött att äta!
I Egypten var oss gott att vara!'
Så skall nu HERREN giva eder kött att äta.
Icke allenast en dag eller två dagar skolen I få äta det, icke allenast fem dagar eller tio dagar eller tjugu dagar,
utan en hel månads tid, till dess att det går ut genom näsan på eder och bliver eder vämjeligt; detta därför att I haven förkastat HERREN, som är mitt ibland eder, och haven gråtit inför hans ansikte och sagt: 'Varför drogo vi då ut ur Egypten?'»
Mose sade: »Av sex hundra tusen man till fots utgöres det folk som jag har omkring mig, och dock säger du: 'Kött vill jag giva dem, så att de hava att äta en månads tid!'
Finnas då får och fäkreatur att slakta åt dem i sådan mängd att det räcker till för dem?
Eller skall man samla ihop alla havets fiskar åt dem, så att det räcker till för dem?»
HERREN svarade Mose: »Är då HERRENS arm för kort?
Du skall nu få se om det som jag har sagt skall vederfaras dig eller icke.»
Och Mose gick ut och förkunnade för folket vad HERREN hade sagt.
Sedan samlade han ihop sjuttio män av de äldste i folket och lät dem ställa sig runt omkring tältet.
Då steg HERREN ned i molnskyn och talade till honom, och tog av den ande som var över honom och lät komma över de sjuttio äldste.
Då nu anden föll på dem, begynte de profetera, vilket de sedan icke mer gjorde.
Och två män hade stannat kvar i lägret; den ene hette Eldad och den andre Medad.
Också på dem föll anden, ty de voro bland de uppskrivna, men hade likväl icke gått ut till tältet; och de profeterade i lägret.
Då skyndade en ung man bort och berättade detta för Mose och sade: »Eldad och Medad profetera i lägret.»